BZh91AY&SYóG^�8_�`pc����ߠ����b@����           ���mU�-6�mi��1m��B�UUcЖ�ڬ�5�Z�SVkm�J��S[m!(6�[cmmM�ih��ҩ��R�J�* ��v[��cf�͵��e�M���-�fm4�jEIE[���I�KV�ml2���hS6V��٤��[�F�I�   �o�[*L�M��gs%�m1I���Ѐ%J�bvf�W�]L��em�;���5l����a��V3p;����̪�E4��&¯��5Rj0�^��AA@�����i_v�Xu���ۭۻv����mkn����b�׷�l�[k5k)˺�m�v�5&����;�ղ��e�i���wskk,ٵ�&�k����UJ�P���튐]l��T��  'U�3�U�Ӹ�UR����J�����=A�4��x�Wl�*���*���ǽ���F�uWU�Xe�3i�M��|�R�����éT"{|�=��@})UU3�����4����}WF��s_g��5�*�ܾ���� hV|�=��$��k���Ê�m���`��|�����@�*��`����v���b��UU"&�>��������
U�|��`����*��{�J(�����I R�q�uR�Ƃ��}pzf�TG�w�à4�F�qB���P�Zԩ��jʦ�-�2Ą�m��'ءD��j}_@z�EwGu.�u�a��Zm�T�û�Jj�k���u�բ�s��Z���`�UEY�giK� 'v͸5KZ��݅� �����͌�٩6D�ڍ5,�A��UUU����o��{U
V�V^��A�R+]Ng3CA��t�P�����2�����
(Qz�@#w�;#�h,��-��z�ʡ&��0��M����G���@���� =��= 
�Us� ��� ={��h��m� m]5à�M�`� n��Z�Xm�`��Z��i�����(��nӠ �� #w��hwC��� mp��wV� Н6� �\���ЩEle�٥��6xq���UTo.�t �S  9�s�@:��;�c��(�7��3��x�� )���F����w6�6a&ƛk,)�fֱo�!UJQ�} ;�q��h����w@��]�@Pq���C�]�{�G�S�� ���i�: 7π  T    � j`�*���      ��1))J�bh10L�����d�J�j       ��@���d�1L�#@�) ��4S���j6G�='�P*$C)SJ���  ��@ =�G�|��������#A̃I��|������IR:�T@�;i?�=��yEw��i��@xAS�T U��H*�����?��w��o��Og���?����"�+'�eUU��@ U���t
 ������^�_��h_�Y����"�Y��8S��,�c���L,8Rp�axY+��(�f�|S����������A=�'a"n'��M�D�dGK�$�I8XOK!�Ě*)$�RN �d|Y#��¤8T����Ap�I�Ȝ,�p�IK"p�8T��A*I�[�I��G$O$8T���E,�p�'
���zT��I8Y$�Dp�l�p�I�Bp�<,���'
�p�&�p�' �I,I��'�A �RNAe'8RN,
C��8Pp�8R(8T���,��A���D�Pp��*'
#��>*p��Ȝ)!¤�*'$8Q)�D�a0�C��p���!�`p�'
�p�,���N$�Pp�#��8RN��!��'
F�!p�' �HzT,I��8Y#E���8Y��)$�R�$�`p�§$�,I�a,�p�'Őp�8Y�I8Y,�¤8T��I8X"p�8Pp�8XN$�Q�a8Y!�A��'
��H�*C��8T�����p�&$�Dp�I�Ĝ,'
��d*I,�K�dG
D�A���bN���8X8Y"�$�*'
���p�'
I�a*I°�G
���p��bNI8Q$�I8T�)8TG
�¤�)��'ő8T���NF�(8Y
#��¢zY$�`p�I¤�(M�2	�I8PxT,I¤�*��'�D�Q4T��
I¢8Q*'
N8RR�p�8X)$�RN�I8RNJTp�'"8X*'
�¤�,I��8Yp�'
��H�I8P�(�� p�������l��Pp�p�8XG����p�Hp�I¤xY��8RG$�,I¤�,C��N
<,N%,���M�A¤8R,��bFʐ�RH�H����ҒXC�D�dNA��6S��'�Q8Y#�Ȝ)'!E�N�#�C�$zTG
A���d���8Y�N���g8S��)��p��p�S��,�Np�
p��p���Np�
p���p���\/
p�����¸a�,�N¸Y�ϊ�\,�c����a��¸W�p��p���
�d�g�8T��G'#�'
��*8W
���
p�
��8Y,�+��p�'8S��8S�|Y©xS�p�
p��p��8Y���xX�g8Y½,�Npѓ�8Y¸S���p�^p���,�\,��
p���.��g8S��'
p�K¸W
�~+�a\+��+�p��p�
�Nc��+�p�¾,�\+��)��W
p�
�g
�N���^�1´S��,�N8Y���c�����g8^p��8S��N���\+��p�
�\)����
�*8Y,�p��p���i\,�c�8Tp��I£����E�p�,�g
p���-,�Np��8Y,�g
��c��+��,p�p�)xY��p�
p�p�
p�^�Np���)�g)xX��4v?�MS�?�v��>~/���78&��B�T�Y��n+��v��Je�ò]F�`�zdQ
�V �MR���ݭJ��p���Xi֩�f9Z�9�:9";ꒉHS�ݩX�,Y%t���M&��r�X���*M��eL�	{��P���ePSF!I�g6�Rx�q����Ko�[���*�׃7��M���f!ra���p .n��7.�8m:y�Ӻ�q�A�S �M�̌a"���[�&e�5bEx�-�^�Bk��:�|NPyF[h�]��KZ�J�Ar��!�T�ݫ�)'"!�v��cV�nJ��#�kN��6Uٷ�f�X�Ì:�O��-�7
y���i[>���rS��"��˰����y�	����1�R�H�uW���=Nm�6�Ȅ��E����t^l	��X���҅a�n��ޖ�VU\u�JnЋQ�,B�v�OT�����3�p�ɧ0�ix�,%,虊7rXxJ�d��1�b"ꤒ�eK�aY���pM��eX�vk�a�Y��'��kWw�o-u��Mh��{$-�in9EU��t��\��l�WNR���ͬ��Kx���v�MJKQz.�e�e<L�.@�MOj����P��	a^##2�fYn-!��@������T�iX:�ul�^e�
�YS*�k�"�L��TVfK��6���-�#.L�s����+=z���]��;�F`37,!G��֩ust;bkoZ�$��n�Ǣ�%�n�]��6���&�DA�i�i��#�Ztݵ���ܥ���H��o4;�6�B&�M�Ū��eeEu2���n�l��U悶\jUٿ�Qʹ2�o5�9>�l�Uf���X���l�'L-v)��ͤ�k �ry��X/�TCG|��۬V+/j�,��"�m��Ŗ�؂ަ�/s/�KEJ��+Z.fQÄH�:�1)&(�͌�o)ث�Ѱ��2�[YQ�p�a(^z��*zU:0���Wò�H^2�h��#��n�ʪ�Ҫ�[6��k�T��Y����
�1$��嗸�l� �{M�[J�m�t�43�����Y�ֽ	�f���ը�ܻc�ؤ�$�)�+��Zp�����[��,�yIX�Wx�ְ�ʨ��/+ٙ�҂VQtRy!��l�q�t�2��b8ɷAK�ȅ��0;u����L���֚�Z+i�v�ʢ�^іQ)����d��Y^�<��rxܤ��rމZ�]ޚ�ܒ�Z����%���1s*�4�Z*#V����b�����;xu��ը2�t����صPe�%�e�Տ�q&Έ��<zv����dnCJ���'e�
S�j�T7m��M)uX�.C�j����֒-�heY��5M�a�i��Fe��zZ�����j՗wM��1Unek�ILb�)ndhVE.��ݱG*��1���r�Ȇ�)r�MR
�ƁM��欽't,��Rr�K7-A��)�S�lQ�q"M�v�����5�jO�]^n�c3m}J=gT���u�huo�D�bڎҺW�W[x�����eAX ��m�.dɱ���͖��nc�R��QoB8�
�I��m♗e�˱f�Ȯ)ۆ�VKQ;�˺Bҭ����Ԓ��B�Uy���b�<�Ռb�Y736T^�ͫI�y肃6��A�L�Qt�ZF1p�v�k�̥o������*Ua>�y���Af�*�q�ݤ����ǅ��wk[�����=�J�C4�PҤ-K�1[m�%n�f�Il射#^bA�!���"��Yq^����	�o�[�PTtQ����QG�B�I	ƅӷ6��)˷�����6��#����fЍ�úq�֬yam�v�s
%�"TPXЦ��2A��D��N����kwVr�v^Q�Y�eA��1�����UU�wIe�����p�6�5��Cx�����*ν�-ս��i;0Ip!n(3k�պuLSCM�טjº��4�'1�?e'�FY�x�s�I���¬E@��&p� ;*'(D�-�'���r?BEm�#U��K�f����:%VL���"K��YEi����h�l�-%���U�$9-�W�&�3X����Փ!�r��Z�V���0���Bŧ,�@븰mQt��v%�K^nB����YD�K�BM3�:m���<Af�&m^k�ŗ)���R�%IL�dkD�M�Y�7u�
����1O!֚;�!�a�}�4N�z�4i�f̽y{���,;�j�j΄�B��na�$�35��t�S7~^̭�4����m�m�T��qj�Up�Ӎ��c&P�,��a#{j�r^)ח�%.�����n�e?k5������⶜wƝk��fVvt�[�/�U4h��[P�cPV�t&ܳ��s��+��A�n�
>�n�<�2�WK�P���^�r��@��)����r��ۺ����.U�n�&.L��Mn�g)<����mURR��;���m;�W��Xz���OU-a�6*���d�jE�FM�EA^�4�?����J8�J�n�h+6��)���S�eSv`�4��T�-Y�P޽N�e����� cʰ�jܦucZ�F
rue䱆����(����MͭLܼ�.�+؞��T���	@�0���NC�Ot�X��l����"2���FSרf��e:���.Pgn	��^*��i�v�F�kI�y��[��V^�$��BST��/DZ�1�7�h��C]�ou�B^h���uZE&��%H���q�y��.�!UA8�ə �u�Ɨ1=ѧ�$Z��33Z�7��1d�o[ӗj�U�]���Y�jA�^��fߪ�Ds)Y�%ۨ�����X�
Lŕ	U!�����:��ZQ��X��9�SOq�fJ8�W&ZBa�45�")�1�(��a��mkj��,Ӹ�&i���a���F�Wm�9e3e�k��)KY)�OAw�Kq
*� �xn[�H���%Q�܁��Mm�V8���;�:b���)����ae�?�Vƪ;@P�D"B�V�L���XeVɗCa�M�I��.�J�y���J�N�� ����q&H^\!䨝�ebE	K]y6m:��CLU��4� �k
�u�!f�b���S��car�F�E�m��M��v�+{N�ԣ!�m��M������E��D�j�N�ФֳSY�wV	��5�d�TСSVC��Rf���E�����{x��L9N!�a�+Ud��v�AT(G�J�x2��T�v(edyW�k	Qb���(f� ��r�ZD��n���R�wpq	6���q Z݉m�s2B�#���:��O"���R�
!�)�q�Z*Z2�R�����ʨ�B��DZuq7d��q�2�.Fz1�C�M�.a9Ud�WJ��u�3+Ŷ��7�����K	kv�M]`6�n\y �v,�r��*�F�:^UI�R��,�4"�I/,�ܦ���3�t�b�X�Tz�1bUԛ��Ќ+s�3�:)Z� #(U����Ր(���^Eq�{y�^�ma�w>)k+!	��ׄ�����1���8��ϞP�0P$H�Z)3b�n�4��ե��I ��Mf9C-�Ǎ�P��e��%m��\5[�����"Ʈ/�M�ō�VM�I�Lj�5���ӆ�Q���K�u4�P)y���S�jL\��Ɋڭ��&��E�gI��*���lD�n�݅S�Fa�j�iY��qxD��;����ݶ��G`��Q�J��YV��YKj�5$T�ȸ����Xh�i+-�Ϡ���o�Y�z�^	R�jVU&B*�8ɢ$���Eۡ��e0����_�ncO<�G��B����'*�r�V��+Q��X+�v�
]�^$�^��_���풥V�m��!�do	:�a�5�/^�a,(^cR���\�fA�jCU<��C�I᠁v�ʤ]m�@ǚQ��d���,�a,�<)�`JV븶*ڰJ�-cB�x�I�h���Cn����������{K���++Z��1��yu��kr�"�[�Q������j�闵�ñBKZ�n�����)m�*�ܹi�ݧb��Ţ���C6ӥ��uVh�ou�X�آ���b���vbW)&��^!,T+/C)j3�V��J�/̙�6�OS$�.�ũqřyrb�hvۺHj$�2�e`E��k�[�#�ee�I����s(-�dXU3*���F�D�����l��@��y�$�,x�����Kop�ڤ�s.��l�jڬ�_f�l����u7r���ݳ�i�i�gj�J2څ�SJۥ��-���Zv:��zeEX�i�RJ�<��B6�6���Tk�V�k�H��fgT�v��1F[��,&H����F��E۩�$Yv;Dȓ������	�\��ss��ǲ PT�G�Vw�8��R��v�u�*�ń��#�βve7T�l{j�NF�:�4:�q=��X���i�&��f�ju3Sb�E¦��ر��`�̊�"i��n�k5d!˿]`�p�W6���#�Y������^�E�`r�n�-�JALK��rkx���X/6ݬ��z���7�2C5��%%�%U�V�K�{�MZ�����w�O�r��H���#���C\FVa�4[G�E$�Y�VU0�ZVU��<;lX��'�[N�SA�`�)�&-!jm��Ł�edcm�.�䩍�:�{���AH��"���MV��ұ[pٺ�*��l��5��U2M�0IKi��3%�2)u*��MJ�!YVX�5��1�;�=Y�T��EJ�sѷY{�[�ˇ0�ѫjl�Z�C�e���;��3��}N�����mǦ\�a�Q�Y2K����n�j���(��E����P�&]e��e��P2�4���+E%�U�{x(:֫e`W:+%P�J�y�țK�Xe�0=ͤ\���Q�2�Ƣŷ�j����e��1;[cCmJЪ�k[�:� ���L��Z�wQnfd׮�S���.�+Z,�ø%��Kdf�A�3�7��fQ^�Z�0�LV
�	G�LwJ��;�`q�t������ƕd���T�D�MZ�����U�8�Jf�-��k4'�ƈ\z�+�6��[�ڬ�)��z%6W�w-I���-�����-X��dr��7N�򜉕�`��H�U�R����*���I3N�V%3�Հ�L6���%e�����$]V�v�X�{Z^*�Su����i�JjT�L��u���À��!�� �&`y�MUeki��ŅܵU%���b
i؊SB�P����eh�u]k�3*S��YV�m�WwQ�M�Y��5P���'YKŁX*�9h]�W3X{v�t�"-���p���CX��g}�ajͷ*v��-fhj'r�&�ȥ�j�:�a��zň�V��bm^��,����'oEGNagX�D�bU�X�P��`���;uj�G2U��TjS ��c�`���j����u@�f(ƣi`8���#����R	�L;xH0��"A�*̚���\�l���Z�U��[T4nf�Ieʑ���%��#s�N�%f���R��T�0���n�5��хb��d�i	qQ�6+��֧�z�r6��Or5u/KT+qۤ�m�im`��Q���i�7����ݓ��k�S�t�M�qb���7�D&"HN����s�����N8��*fi����zjڰ�*��ܗ�RӀ�M$孱��`��$�"h̍�
�9�F�Z]���*r]e�*���<a�E�
���oq]�jê6�Y�XE��ʢ�C�@�{CD^@��~���ЯE�{�݂}��*��`��}� �G8"�����	X���i k�bn�%
����b��b_hC���7�������M���_B~�4XK�ք�L���k�_V*؋>l]����a*���`���8p���)���>CM�,!��A(�,W���l�+���R�g�O����I���/���AH*��+�m��|����U���g�����11����:A��
�8��O��[	�Z�y�E�di!�g��haB���t8��b��7 �O�`�Cp*`�3�C�0�a�����hz�U}B��3�IayG��$=PUh�E?�PR0n�wC6�#_�S}���h��
�r�$!�KD�H,a�T3�>�!������yd� �>HZ����U!3�kД�3�^أ��<$#2�V�_
|>phaU�ފįZ�b`��zDx-P�8-Cg/�DJ���ׂJ��7��pe�Y�f�vaτ��'��0e��`��:���n��	�����ˆu|_��l�)0�s�11���8	�U�&��のա"���|����A���P��M�;�w�Q�5C�	��ѥ�����}㠎���ƅZ�-?�z*�r�c�#�X���ऄ�)X샕
|.�H��[��DI�W^8w�=�Ff�y�7ӟ�D"���H�V$�R�1P��DMaa�p�x:bQHJ�����RA�	A�,�j9!i�j�J�Z�I|xZ���\ aTX��R��T�-��t%A���	`H�D5�`��,
�*��
Hj���DM_Y��$�H$Dx7`#G@��b8;hX�����غЯ�@�ǐ��X��Xբ,�k�f���/�CDic���&��d�Hg0������H��L����u�JC���s�<3��J[񰰈��`g�P�b�}�ᴅ�;,:>~���^��HV�{�1P�c�܁�4�
�/<�L<�����աU��3(V�K��#T
���>7�T`�Pja&91Ȉ�IP+"L�(�\-p�_=��b+�����uh|GJ��D]����n!�BV��|pW@�	���.���l5޺0K�>r�e
�*li@���t�g{xf�6��x���قh���m!��,5T"���H�;��po��������{~_{����C{�G����?��j��>m��(g%l�Uض�����ս��N[A���B�:�Y�]s]��)Ü��t�S͎���T�q�w��.Ά�^�ftќ���rױ-��'Cs.?�&ֺ�g$���yfDKztʋQy�2o�ʤ-���.�IS歍�7��&39P6暯dJ��m�1��N��D��R�fr$[u.oqz��b��)n��J��ą�%h���V�v*7��^�؊f�\��&Ɉ²KIw$(m+�,彟ǯ~Ys���Ե�j�8��c�d�f�2��Ǚr��3Jֶ�i�7��no�"����(9�]�d߶���J�X�\pGԏ,�:$*�;ۧ;'zlOM3�)�x��:a1��ܻ#Ǐp]�s%y�-y��J�m�p�-�٢����{�"O�`��+���Km]�NЭZ~�s
ɶ�Rc'bӘÇiڠo]���1���V<��5��w�)*a!��]n.m7���]W��R�k�ҕkp�b�k����y�e��ͼ�8��+^���-��-���q�\J�;o4��;�ڬU3ut�ԑǱ���6�O����R��O��^��Ý��z�e����%�Vv��X����V�u���r7k��j\8��U����W�.������B��܏���a�v���I\��Z�,�qa������N��v�5v�CS�����y����˩YR7���:�����eں�hu:&q�l�bŷr�]�M�i�Z�Hk���ש*��tZw��tU�,_c��4i�B�jR�כ�2�k.���ͥ�0m\�v��u���72fR�"�IM>B���B0Ty��4.<�Imu[�v�E�n�C�v��,T�w������;{ؒa[M׷����F7q����(��s�޳O���tt�ٮ_\��u����tw[R'����:�û��
�b��m��%�ӓ�k�۵���T
��I�wU� w�}ReV�Km�R�6r��0g.��U��+քLacԬ���ҭ���v���"�D)]����´�c+��"n��ѵ٫K�m��;��7�&�ۋ-���U�ܫp����;&n���ޛX��5��!�L|7U[f��\����8d�Fq1�B��l>]�
ׇ�mW:�;\���L�;�K-b��z`Ò�ٔB�1�A�֋���YC����>�m�
��Y��˵o���ab�(�U��Ug[聽it�Z�ʈ���P��q�/�E*&����N�۹�U��Y�L�:�Z��ѷ���u�z`����s���6̺��O)n�S��vS��Sm�x�����	��mQ��T0�.��ԍ^��s���X�F���:�-�w�ɯ
N��xs���Ǹ����Ô�6kd&j2G#�mm]��8�3S�R���TmXÎ+�],�4wg)r�h:��6���,}�U
������Jִ�����l�)�v��7��T�m2�kǯ�t{��7����3���6��Ⱥ�ޗS���;Y�a:���Y��<Z�WYN���_��6e{����b�b�Jv�ԏ>f��[~��Ƽ�at��qh�f�U�d���B�^S�pi�Y��s.̣8��۩8�fIL���-v�j�r�������2Nt��r��CG
��il{%�ľ�f4�&�K���ʼi�>���V:G��u}�Mj��н��pT�4p�Uq��0QiQC���ܟ�s���$���c!�m�o(��w#��u���c���7�]p�)}��n��ѽr9�鬥YQw#��T{��Ҿ|R:�˙�J�����k��\Sz's�e�U�R6�c8�:���\AgE��Y m�y����z��v�ҋ�9z�7�v�rŸ��R)��yuKk��f��Y���ׅ�D�'D�j"+[}��;�Ѳ7�UM齅��1eN�*[����s���YcqҖ�ώI��M�쾋e\�0�-�|q�v�c�:��W��V�A��}ҥ���(QDf��:Nom�v�]l���|����&���}Zs�p������zfe3Dw���!N�ӷ
�I=��_&.o������'2��8�R{}��Cv���e��s�wu���q-ܳJЩ�x7��c[��6Ҷ���[#sLF�����D��ŷ7��b��%�房b��^����I-�
�)��(�5�L;�����uAьp:$�ռ��W�"ܪ�Or�ӏ$���G��W5�(E�+�yqm���F�&[A�9n���H��d���<��=�j�3�7�g-Z��Y����:m���X�	�7�3����Z���<&�;�{8������a��e�t�nV��k��w*)p��O�P�����W�1�'+Xf1U8JklW��N�����\�DcV.��)j7��Rw�;�gp}ΤU����q	�HvB��O>9��e]=�Tl���^;"��5����NUa
''|�9]+R�Te���e���e��C��-[��ֻX��1Ej�9a4TN��կ@�T�`W.��/����ݫ�s�=U}�:��)`.=[�{��5Ϙ�]e<I��>��4Cq�Rҩf�P6��cٵ��3�GGV�L�tMp۸�fx��j�S¦L�svܣ,�w�or�yY�
eK!�N���qN�ġ��a�|9^���z�Z�Q��܍�1wona**�r)�w�|��M�A��ι�nc���Ύ�JH���;^��a��cשB���*�"�KX��A�A���c{�η�F�.:v��=��`|W(�]����n��!�-I0o[����]v"�]��g)�8.�.�GCK��O����fͶhk��	��YC��'V-5F�,�h�"�,f��I<j�Y�֦�������4�=ƥ-���ٷײ���z
5ii>X-�!����`j�$��A:Lr�_'`�u�Ui5w��}�M=�K��<1Y��r<����ޫ՝����P{S*�\���z���#������-9��t�>�[�r�c����٣�N���x��h*�u��5y�e��֯��诪�pٵ��$��_y�l���\�}xe��(N�q�2�J�I��N�Sp"q�rT�T9b�%��ƺI�z�#�Di�_*Agm���NY�.�Y� �Zs �B�4�<�HJ��DޙԋH�ͬ��}��\�v��L�9��7C��L#a�ݑ3V�++�'���zԕ�1�t���7w�+�$�騇��1�d�����e5.�ִ�@���*������nY�N��Fo4��2�������1�K?#�f�d=KK�
R�%%:�c�)u�x���v�֫���]���Ҿ��(��o�IqWNu|�h�N�[���V8>�b<W`hИ�V�e2`L���UR�Kd��B�{��%e����.��\�Cvs�6����\��v:����֢Yvw��¥c��r=1E٥�]��ҵ������h�}h�a/��jA9�7
!�����6{�p0�b%Tz���1N�f����2��v�H���v���^;�46ɼ�{�Q��(;BaP�S�E��AraW��{�.�g-��U�3݀���T.�2�v��a;����ۣ:��K^#ibZ�+-����粎:�u���DM�˻]6��M���2vsS�V���.���y��W%C�oW7]���:��a�&�����k��YQ�26�8H6S��b��b���O3��Y��am����B�_NC�*�1*c�ot~xc�Qefmq=ӴXQ
�s���y̮�{���h5��f`]�M̛���*t�AZcW�(G=��s�9*�lI]�f�g�WYUǥ��y�//y�$��JU3*c����8��t^s��$˝'�wҶ`UR����tUV[]�c�Ԉ�H�d*��nִ���ccu3�:��a`��l��}��c�M�JJBE,��J���k'Q౰s�ӛ��GVj�uY��X�$e��=V��fkE�!�%Z�q*�B�H8�������
�Nb��Z�M>W�QaV�̱?hY��G,Nt�%62�.;��TThcb�w���{�}��jQ�b����8�_Z��n�Zj^f��ST���� ��^�U��WL�8�l�[ִ11Iks(�o7Faj�/��"��ep'a#j�'i�r�,�l�g�1�6���35�7��=�z5V]�n�nZ#(KNͻ��I��n�W�v�R���VrW-�Vv�#]e�MG�ۋ&r�r�%���9ƉB'�ɻ�K��h����<Ň��ԗfs�b�@�,�c~��1ΜA�C�H� ��x�S�9)�\�̩/���8��h�VE��rk�G7L���s�_s0�R�c�ز��h=G���ֺ2���N�g��ϲ����I3�*Y�Gl�(��_[pJ90f�%W�[G��TT��o\�C�#.�ج�=���J�_e�r�(��jt�q�]�6����Pm��f�憷u&:���r����B���Aӕ�G�Zo�j�rN�e���D*s��)y�E0��Q����ү��N�s�K��sI�0�s���Ƴ��\kj����S�'�s-6p=�Ќs����Z��-p�QGH�P��������]Ԡ�5�-����p�q$YK�kB��kp=Hq��y����;9:�}���c��h���
�d[o;{�m¹�2>$�ﶈ���<\�9,��y���������i��]�C2��d����rG2���e�ms�|}c-_<]W'L�:��lm�(�F�W>搙�4l�p�	gB��+R,�.�o4���4���0]�YF{E���2)��ǗA��(y�
B2^lZɖ�R�B%�53R}:@p��o;�J8):Vz���� ��]�R
���)�����x�����5�vQ0�]G�\�UEG����\ʩ���'�����QlY&zU]m���mlMM�r��T)�ɸ6����Y��Lb�z/���de��}�9щ��uɭUM��e�˩��PZ�U�Mg����kwOڹcy���
ą�PMb���뇷�5�@p8�aFΘ��Xv4���w)۷W8wWkT�!�҆œ�[�h"��7�x)H�V)��QmFl���+vv;���s���mU"�p�Y�%��-�ۓ��4�eP��kȹ����c��=2VY�sF�ƕ�MU��!iVe�˹]�u^=�}mSI��ȋܰRɇv��772�7k}�']�$P}������Z�A��4�����9Ԝ�sk��Hrr�Xm�N.L�*Q�-�������)U�Y������-����!�CZ�wX��mw���/hSeƋWv�OeEX�n�T�'��aM���l�^�HJ��[�(����qf�lV-�Q���	��w�|녗�3*�� k,�Ӭ�dsd�s��N��i�B�+�;��w����]=�����ʫ��2��������j�O+�"} ��\�ҤP�s]Ϟ��oc�w\�|���
̎�ʫλӭ�����cu�_��Y����>r:��]ݺy�[X�������hv�qIs���fI��#߸fvџ37��YK�%P�����ˊ2�ỤW��NT�K=G�)��d�b�o*�\�������-v�q���n)�kv�w���"1��	:��OX9Ժ��Yr�o��_�n�o����Y��'���:q]��;yu�p\��/;�w1��Gwp���]�{]}��ܟN]ܰ��˻�}��l���ΧZ�W�w���+�'+�s]Z1躁�b��_h�����p�|��g����]:wu���;����������������������\(�W�6�S�m�Ǌ�M��i�mXګM��xǍ�x�獪�x�bx��jڶm��Zi������xƕ^iZz�>WU����V�i���xx����c�4�m��l�li�1^��lVʦ+�LW�Ux�զSjc0���ڥi�6�cI�F1�G�ǃ�cJx�ƚzұUX�M��0�X�V��l��EVi�h�SƘ��*��ٍ6��+ei�*Uclm�*�+cM�ƕU�TҶm[R�M��V��[O������U����ׯU��M0�ѥz�M1UX�Li�T��i�x�cMc��OSǇ�Lq�)��LW�6z���c��`���+׆=<xڶ�3I��0�ǆ�6c��J�q�>x�lm^+Ǎ*m����i�Ӭ4i�L1�q����ͽlڼRb��m*�x�z�U�UOUZu�4�*Um����5����SF2!�8���!�B���K(����95�P!̱w�Le���śIR}�G˩V (W��ƣM�@3Jvϋ�7p)�0�
-�������!����Ȇ�(�V��PJ
B�@��#�2�a�4b �M�� �i����Q1�B����eR�~1|$j�A?�a(Q��m-*R����"�(�M�"��H Ѩ�B����y@D(#,8\$� e@�h9���}ˆ6Ԉ"Ax�Ѩ�&|�!���$� ����Tm�g��Kxw���m�A�|�D@A:�����w�U?> q *
�� �����G�_����Hv����3�{���~�x}�$�>�ʝ�YR�%3]y-Sm:�ay�p��/���H��ˁq��ݓ�1��꧅S�Ŋc����gV�Iُm��m;�����It<�e����VU^H�s֞v�ie�m��JZR��9����V�׼�!o��w��e��i�E�u�ڗr͊���T�m38�,W&Λ�e��+�LU���wnO�0��NҪ��!�s��˖5Һ�G �Sy��T��eGq�1-��̑�˃1�N��2��Ͷ�n�m��p��MS�;������F��7C8yL#�nf���ug(�i�]�YV/�P��&�uy�I�sH)�^��J�Y��]h�j�G�Dp���Ƃ��on�d̮�����'��(/�����Y�^^M�r�+�&M5:Qp�������.ʭLc��op/pC�;رI]�[-I\0MWV�⥱WZu�BŴ�ڽч����T��I��Y�7��r�=]���!�q��0a$ʳݘLn�����괦ŕ/��IէtQ�;e888�HK�(�0V1$0V�Ǹ6�0�I�=����-b�gJ��HB�1l����æ�8t�ӧǧN�0�ӧN�:|t�N�:t�ӧN:zt��GN�:aӧN�6t�ӧO�:aӧN�:t��Ӧ��8C4䕓������C���4�O�7D鼪O���P흖^��q%�I m-7���ݿ�H��<��;���L����k�Ze�L�|)�u�b����m�r��0b�w>�SM'�B<(q���xQ�ŵ���Qn�i'�q5NWȢ�:�x=�h�Mʮ]�b��U^i(ړ^k��j}nuwXˬ)En�d�:ÂS���y.�-�%����[�V��}�k˳,r��9*���ꋺKDs�C����Y�ܬJhNn�`��g��N�R�71��Z�ki���ķS��vZ�BޘGm�a�6E�bm�7����W�ԥ�7��
؁�5Q���D4�X-ff@��^ĺ��%��˳��	��G7k��Œ}�褠{�jT��1Iܯ/F�Q���˦�D<	ŕ]�d*�F5ۭh������Y4�w��1�tl�sE(�e,�5㒘}���h���<KeE�U�)P�d�^J9J�Tfɨ؋#Y��z�R�#�)�G&g��\Z�Ԟ�S�Cه�Q��v��R�X2���xuTƃK-"%�&�+f�'�4���{��3���w�H�0q;9���k����k\�M���8l�ӧN�:t飧N�:t��Ӧ:t�ӧO��)ӧN�:t�ӥ:t�ӣ��N�:l�ӧN�:t�ӧ�N�:h�ӧN��u��,�%\c�(T�'n ����5�^5硚��<b�TW���j���yPc3S��s=�W�U��Ay�A��}�1w�!�LmIZebiWq��D]���EF�9uִ��c�K�C���]4!u�7�
��u�V�\�'S����e>
P'��J��=�c�{Af�(��b�TPA7��}�d�h��0�!JS�	�h,b��Hm�/y �𫒢@�v�̿��]�	R�GVs��> wni�U'��6��ju�j���K�M��� ��e��(l΁��y�*t MU�E�Gu��@[Λ�P�����f~˂V�.uw:x�[o���0����(a�ڄJX�P����o���=	�Ä�ڡ����	���5�+��*�^R�\����T@��(�s
�؄	ډ��pm�y�r�кE��{���5]v ���H�{~y��,�����A���u�{v흦C���UB�EӅ�ڽ�2����a�;@L*}ŏ��l9��Z�����hiet�0�b-���v��u��2�]%Zk�W����t���Tl&Gm��0�>�ᔳi��`�4Ό��>Xh�\�x^3�]T=�q3X��"��M���Ƕ�붯;%��yv�|��bG4[8�7�R�&���¬����aX�� �����@X�"%tH;y�m ���Z�$�-��n\;UÓ4�U�
��sF:��k�U묮+�Z񁇇JS����<:t��gN�:t�ӧN�<:t��GN�:t��ӧL:t�ӧN�:t�ӧON�:h�ӧGN�:t鳧N�:p�pl��g렚byƆ6��:E�y�����`c�}�-S ���HV���Y��b&���1�(w*�G)az6���y�{�]�,Ђ�a��Y݀o���Vp=)X��x�e��n� >�g$x��m��i��۾\.�
�2��e 4���r�D?k��֤��!�V��n��C�}^�''�l;�wt�,Q
Հ���X;�u
q�����Jˈ�V��Ǿh}���Z��ArW3v��x�������($h�z&AXx�r�D-�Y1є��x�k�-��Ҽ�|Rk�<�W�v�g��u�M�D���X�(������K�(+�xoWA��6l$�N������-g�� ���@�	ͷu��� 1�)�BJ+�yy��3�Y3��XrA2�X;$��`*��0�G�:X~��̖ڰ��)�㵵π����'��l	%���D;�Yż����0* ���1V�ͽ�On1�距\�R�؅�%�[�����Y�/w;�bg|体xM4o5殫
��'�q�߇h��}�:�"�ѷz��Vݳ��������\Mof� v�u�3��5U�:�X�l�k�!�:.L+��P�,�f���*�[��j��ӵ�+{B�|��U7X�4h��awK6}�Vڕ�]����n8:��<E����؝}a�܊;{����s�͜i�];{߾�Y����ke<8R�8t�ӧON�:h�ӧN�<:t��gN�:t�ӧN�<:t��GN�:t��ӥ:t�ӧN�:tçN�:t��ӧM:tt�ӧ�N�fpS1��kCh�����/����z	Ux�k��F�u[`)[*[�]�V���1�)��*L�\}�]�>ǘ�2�!��B6�!���/��nr��f ���+r���'��N�4�׋���nԂ�WF��\�,�r�< ̳Jq�D�Auk�㶖��V���X��0ش.7gx�B�[��M�����l�������[�I��+�*��O�b�P�v�Of���{�iw.�f�M=TZ�r�e����A�:�s8���4�>d��v�S\�w��M�l�0��n%�[���fWuS5��	$�k7�*��sXl`�Un���򊫔����sW�nt� <��L��yM|k_Wp噫��eK]7̭��V��y%��U���Eĺ�e���V��s�I1Rt�-�gamF1!x+{���u}(�����#�}x���{'.�y�6�f��*�j��eO�ZY���E�����x�TD�HN�C�`�}H�H�Ю'W\��<iF�`��ܰ�����r��h���(�g��-�Ux�r���-���6hN�*vNWW���Owq������]��X�]G��S���D@@4  8:t��Ӧ:t�ӧON�:h�ӧN�<:t��gN�:h�ӧN�=:t�N�:t�ӧ
t�ӧN�:t�ҝ:t�ӧN��I }�rU�"yJ\��,E!u���0ո3Jg�ⱋ 'H�B�~[�+�|*V��>=���4̪�+1ask�����	3��9�{���r�-��O��{�$P^����N�M��%��X�Giۄ��u�*��|땽W��7A�`tl-���>zn�kb��5�]vY�Ϝ���t
�Ո�8��CB��ɗ�&p0Z�a�Bλ��P$݋R�R�c�kZ�,��D��gGj��e�y�M��V�c��b(�x	,T�n�e�E>O�ò�N5ܹ��Y�Xz��%�3�XC�@�*l��}��Ψ�j�m���2�bS�v���-f�4z�oB����R��݅qx����静�N-���1YM�l�E�MI�W\/1�C�N=Gr�	F��84�l��I��E�m>��'U㜬e=��Jp���s:��<ɳOo�v^#3/T���y�u��l�f��׫�7|��S\�AƝ���i�N�k��}�F[p1Lf����`����g�kt�q����Uz�lw��%���&��k񚃖��X�����@��Y����R�к�f@�ڔ^�9�t�٪oj����x�����ݖX��Q�b�T���^$�Lת/q�-I�;3�.�@�]U�1�"%��p���:||p�ӧN)ӧN�:t��Ӧ:t�ӧON�:h�ӧN�:t�ӧ�N�:h�ӧN�=::t�ӧN�:t��ӧN���8	�Z5�,k�]���,�0S"���W^�Ar��
}fu�#d�˭A
�Ɗ�z�3y�⡤V�!j�v	x�Dus�����n,F9�jP�޾�>����\.,C5:"�"�E{����x	�l/_I2�W]o_�ܫ�����K�4ki����ԍ�cN��`I��J�:�f��\�����Z�R�{�3�᡻��k��Ii��/��3�$�� ��lC��9�q��\e��oT��-ڶji��B�G\���(�HJ�g�H�]U'[@U��.�F<�$�r]��v��xs\!�(]^\M^�a��c��8�n��:HA{�g��n-6��c�d��y��#֢׫*�9�7˯�������:r��b�ո�Ty�XM�x0'ɋ�qǩ�ݜ)�Amnu<��!�+�1��#N,|���!�;���+C�Cc�+:i���q\�r5PK�8e�U�e3y ��k4.���q�i$v�Jܼ�mR�~����չ��� �J�)��GT��Z�i	k�̤vkn�v�J"z�A��_kީ�U����aՕT+�j�hTSs�'*�,�%ٝAG���r�F�ܷ=���+�c2i�+9U�V8��Ñ�G����u�u#w��w�GS��{QΜ�tW����[ռ�����aM��㧧:t�ӣ�N�:t�ӧ��ӧN�:t�å:t�ӧO�:t�ӧN�:t�ӧON��:t�ӧN�::t�ӧN�:e]���}߷�������N�*�Z��#����e(���Lo6,]l�eN6fuح�}g�:�Ӱ��oCKb�j���I���_m��w��Ҭ�Ý�;7J�����}w����NV�'q1��Bõ�)����qh�+�a�x���M&.��� �y����x�9�+�#��p���޶���(���nL=g+��цǁU<�N�
���k*�_ou��:3�t2�W��*���\�)�5���)��������M��&����U�3-�珖:��UEWfK)+��o���5�Xs(W˧h�kL�G0>e��[��y|�+�DO�a�ln��՛��^]���h`ĩ������g*�5�����+gf�7�Y��!�u������έ��gV^C�h���%B�v�*�o,���i�e�'2�
%,�d$T7�\�iHGWB�+����R����v5q���bH��rW.���PJ��𙜪���brY�<�e�@��!u��H�׽Reݷ��"���ݜ�sNJ���:�6M'��J���W�sZ��]��V�'(6#��EeB8i�0a܃B�t�e�_G���s���,��Dٺ�w�3���WV��C&�S9�;�����k|��r�4>=:aÇN�:t���ӧN�:t�ӣ�N�:t�ӧN��:t�ӧ�N�4t�ӧM�:t��çJt�ӧN�:p�ҝ:t�ӧO���_o����\���ZyG[҅�%a���EeV��N�B��n�
I��=Uzv�����Y���Ǟ�n�m��~�9�! D�{\�;��,���''C�5�c��V�%���I֚�b���Ư3�ct�f�o�x'I÷C3��u�����E��f�y݌�
��&v��������o�P#wU�M��˝:���u`SI����%⭫�v4�o�.��W�$�xyMtb�R�b��')S�zV9k0�C��HĶ�m��Kh��Y}eݵn�hA �x�����j�xP}�M�B�OY0k&+��3EJ�{A2L�Qծ���;s���^aogtY�)�܃V������UmN�����N�'9<ל�˝����Ɩ3��`m>M=��D#�J�&��An�\��Xiu)�S�^�\��={3�l�f�۴Y�u�Ȱf�-�͝Y[R0���C��V�EUXw�jV�Ov�/{��z�W�!�ci�hp�m�SGoEƦb[αa�1��Dm�5vaU%/�>�8���-�C���z���Ł���h���N�u�vX�\�VEJ
ɻwd͆��Y�D�e$n��Uї%3��by�vdz1`��Y{]ѷ�	�گT"ֽR�h��̍u�p��Om����T�����hu)��!ϖ*N�Қ󞒈��]Z�Fc;"mG�7�t��9"�}��
�W3+S�t�4��P�9W�-��W'تȯ*E��z%��A$�С��D�Q���}+Ȝ�����^�iwP]e�N;�-��R�Y�s�#����h��C��w%��<!!�]ӝt�On�*,��������|��IJٙN�e;w]YR�ա�Ky�w{�-�q������`a��$&������ƻ����aY�S��Cٕ�dӕ�\:��Y��5�,�ȹ	�v�e�jgaX55R�S�*>Lw*Ѫ�2�K�t�V�TtLA��Y	G���Y�op��H0��3Ǚ�V��[;ef@W"K���g�����t��N�Yȴ�*t�ݛUo��фiQ�v����01b��=�fp��{84t�X�@�(���pV(;�)Hs,�nrNg*��!�7NG�}�R�9-��5�\�3��$e����NZ�a�kv��}�$!�c�Z��ti���H8J�ϩu��y*9G�)t5�͝����¢�����c��ԟ-v�=���s2�S���c�_eD ����	����R���ˆ�x�/j�ﭷ�/������I~���_V���>C������!�"d9��$�u��eB�A��`��P�P�[6�Q
�b���F$��4Q	�C(!l����"BDD#�aa��6*�O~����VΝ��[�P����y٧o2`+�˝hh��N���!�'�[�ɽ���u�r��Y��V�tj���!�Ӵb�������A��BH�N��Ũ�oe������U��G�L��8��d�ѓ�n����a:�"�b�������n��ʄ.�\���t�O:�T.��d�@���L���U��]ڜ����]�p�rK��C��22�h���Eܙ�Q���[y��ʮǛ�]��^�K;^^�T��9�U�G^�������g{@�7&i=�C���C����'����.�QuTX���c�ި����ڱ���3�x�y�[r=b����fΒ>9��Ƣ�U�]}��!���a�����Z����\�l�9��A´j�K/�.8�q�)7S�Ws��d'��&<�U�<�q)ʦ7�Wy���A�b����M���ҹ��n䢭�s+��ܝ��v����c9.�J����+�-^k\,>�l�6���L��{�i�c�I���Ww����*�T�D��oU��{���^�Y�'}˕��ݼ�u��ӟt�P ��8P�`�[M�եmSb��z��J�m�+ƞ�xي�ګ�xz�G��i��4ڱZi��1XĪ�S��m�V�M�ZLm�mZmU[TکX��ڶ�a��V0ҶҴ�Zm�V�V1M����m��S��bp2�e4���\*.�%��B ��B�m��L&���YD�𺔡��~��񐐙M��a��BA�AA�$��B$�� T�wA�VF�QLN�&���%��ʢ(+��tXJ`v��O�����ů+)l��M]Yz�*�VU�R��7���p3(��2+��(s0��Ř���c�f͟�8t�:���1_��U+X�c^Lƅ�UVV3�V����ZeH�I�eIk3�Ƴ�i�eNTeеh�!�2��6�.AB�Bfb�ʙBe*��RթKK*J�.c1p�˅ROǦ͞�?�_���-HeFUU�RLR�)i%��qU�.c
��)kR�'0\��8�[Xf`LDH�ʌ��ĪfcEU˄̘��X����b��eU.<�f�ی�:tѳ�:y�U������%,bԲ�Z�L���X��Y��a��5K��ȸ�?�4~?���\�U��k���QD[�E�X�UV�F��f1�cjն[��*��_4Ɨ-_�4xzt�ӯgعXZ�c&[V��h+�l,(��3ir���-��e��k�m_��-�:a�ç��:�e����Rխ*ohфX�F�a�TMSN�
3,�:t٣�O�<���R���**���6�Y�Q]�4l[Zc�kE�4�X\��a�F�Pu�9��H�MU]rf�������ѣ�.��-�C��l�I0�L��D3P��h7��Q��W�/Ǹ#��5є7y�w�{|▆���s���c3�52�LR�h�M�F�z�cf�a��`�� �  @��6�j4ۄITu@����dQ����c�F����^
�D�`�
���*�EF�r6�|i�n�P��LE{K���\3sh�Ɂ3@�q��|z^�0��$�CE�mvۡ+}0���8�ǲ�r�����V0�-����w�)�g�������;�ǢLv{�G�Y�헴1k��u��w�G��j�(��~���@
�ܩ4�fw�6��~�O��=��?w��uV���ٲ?��<��b��,��<�{ zJ�{���?e˝��{��s�����nP�u�S�q�8;���{Ր��KO����n�=X���J`x���}�:y�q�����a:-�YU�;����x�T+�/�s�}�sz�{f~Dwz�zOk��� )��v4�E�:3d��7�H#D1�b��Dm��
�A}�*�z
�]���-�=�S]�m�(M��� ��Rw}Jٕ�=�&�r3��h�*���VZ��nܝ���a�{Ntx�D�fTVH���9ϴzy��/ϵ�ưJ��ݗ	�	�SI�i�O.Uc�S�KTen[C�dn�����2I�/WW��/?�a�;�����v�QOƮ�s��ɾL b�ؾ��6}�Z��`?��0�����w�;��1U�uwun��+�>��������'`s�8�������N�<���=�]�xI/}�G�wB�\�{��_sC��Y�lV�	�d~k���ܽX�y��y�Q�f�k{p;Ӡd�hi����Lq����qx���NxD�I���憃CdPa����z�	Ȉ�'���y�N5�ϩ,f��#�"�@���½T ���p�W����G�����5<��{�f��� ���G��T�G T��1,X=� �����W݄H<��>=�X5u^�@�x��3l�K�8E*��}�h�xw��V��>�/׾�O/��׳}����KCv��f]l6���˩+9��j8oo=��)���_��Vx(g���ۡR�<��O��C޽bk��/��swW����xswpk�ԫ�ө�Ŭ������J�X] ̝������>W��G���͇���w�^o�e��1_:~���每b�~�BV����n�1��t�.����͚�ޮybN�����{���O	Vp�����t^�a^���)�j	ل�x��đ��+	ќ�v��_}q[�R�����7<||3;�3l;��zr���ʍW�sc>Z|C AA����U����N��1�pz�}~�p���t�hhyʓ^-�X��a{�����_����S܋z�nu�����	B����y���LwD�Hp����di�m뜳R7?P��8_��v=�)��ɳ���M�9��NѿsK�h*t�8}�vA�x]=w�}��R�c7�b���a:�U����wr�͊Ԁ�<�vwM����~��it�+ 5�+�'RL�\~ݣ�Ҍ��3I`�{U鹑2vV�������̛˹׽t�t��h8io����2�W<�*���~4 �PB�b@�ELbXP�����P���Jf[7�*�W�%�%Þ��I��lv�.�����j�Qtu~6=�H���9��z�w*���.����s���d
����;i�nj�q?13�e�%^}�d�~�y��UX���e히�۳�~ݕgM5߻�<*�4�c�=읹&�úf���ճ��r��\��ݢzz���}M{_pR��X��u�=�yz�0'S���5�dS��<�j���X�<����윍3�'v�{�r"�]a8K�gA��^@\t�R*�����5�w�޽���?yt��9�;U@Z��rС���ܚ�p���c��0;����"��˹R�#�L�wn�#���19��� VQy�w�;����ݔ�zr�����?g�����>�p�0�>la�����x?MznȈ���;|,���θ�ݛ�.���o��m�0����z��v�@��U���4#�ݣՁ%P�3��\�Ve��M�Y~*%�V�t�~uGBA��x �t���+ʙ�C�w�k�d)�Or��P|��(�W��j,�l��B�HZ�{%���یX�7�5o_��٦�ۘ|�F4Ӎ4��? ���5M�H�$

�JŖ�/b���c=lh "D0@��џ��w�!��
��#P�� N��>����~�mЀ
�����J�>����u��ĻVT^0���!Y�{_��r���|�>��}`���]`P#�n�����l?gz��]/J��-px�{KC��<��fWd�@�]�x��1�{���U�<׵�MgU��Ty�g��H����}I�3��r�X��;����x~��U��97�z���gǍ�^���4�'7�ޚ��/l��|k��R7{j'����|n�Ku��rrݧ>��+6�Z�q;��?g�b|(�c�<V6��W�S�G� hxϞ�U�������o� l{�}�OOK�G�8
"�6@�ho���~����� �6�6�P�h]�Vs[�w3Ǻ�?@��m�z8�x��o����O���e���5@A�S�Ǵ�	P����M̔��Z����Ֆ��`�ْm�>��(pmh#���"*��������i4�h�z��N��Һ���L�'[�[�[@�k�-����Eb���g���kv��S���>�]d)��&2�0�;N��W��_{����{(w�������;t�7-�3�]$s��ݓ���=��~��������׃���@F;�Ov��m�P*;N�����b�F�lc�~�1�(�'6G����r�NL�:��ɧo���p�X'�Gb�]d���I��� �T��|�rw�c�h������7Zc}ygoX�j�f5���0]5�}����+��ֶ�:��6l����S�u�� ����{��+�{a�h��7� ����1'8�)���ǫ�z.��܋����s��������=c�g|_�|��z�@{.��
��@�V���\ĳ��m�X"�脑���*��̰N9�@Mq�<y�fxܑ�٧'�`�O]zt��Uw�C�h��R�=�����+�V{�uꕷ�[�zL4E�ga���d)��X�~nj��W#8�pՆ�b����3�лv�8%dJ{j\:�ص�2�>]�=���@$�w�}��	){3.�ǣFT~b�XR�Ւ���gl�M8t�y|�^>g�6���-�cM�޴�����Qꝓ�st�>��i�R\�e�H��U>��W�Oz&n/�|vΨ&��vj;d�����"{sWy� ���e~V!*�h��ۼ�/�F�u߁��.jsO��ӯ����R�{g۠P�����쵟Q~�'�#c.hxۏ^�6	�� q=w���k��*�s�M����dM��I�W���`@�c B6�2?Pn0�.pq;c6�=�'s�5�uY��!ֽ鼅���O�~7~�\7�i�K �`y��u��D|��$��rt9�]��=<��>��CHMX+a�^�O��fF�9ky�-�R	7�Ih�����w̫P���:��L��so��x��3��M:��z�ފ�O)���>̫���`3�������ս�<���~y֮{Wy\kV�W=�~<"�:��SE8��,J-�**���<�NV!�4�{�^�;����rd��OwVon������ٛ�
��=A�mV��(/��5.Hxl�P+�V�uw��u����p�����k��@ve���=F�P�O��X�����s�����챀\�����۠(gS��>��XZ�+�"v�U��}�/=��^Nx0�C ����7�M���\���� ��C�=��{;}u�/Hz����~�묧�p�hcվE)��H�Jx$T�3G{�VN
����Ӑ���J������j��.��K����*y��%t¯4d����,oRcY��٠ǼS��]�,�K�	Iu�(�~r_�'�=V"�NDO��������E.�
��*�O�r_1*�J^�^u�0*�l�I�9�<|*���\�-�׎�g����3��l���x=���o�t{�P���<8ݭu����˪�J�8n�6���Z+D��������srIx#�-�u�y��5{Lt/�5���!��{2|�W�@�{ʻ�����!����2';E��u��&�:���g���y'V�^��n)-��	.�.o7ףH��U\4�nC��)��ZA���Sxy��{��Z��㻈�I���0���J��]�	\��}J]�t�<y?e� 4�`������*p)ēX��Y�����,?�t�<_o<S��W�\w�Y.M{�n��[����.X�t�G�������o�c��Á�:(ݞ�"3�ߜ�,�k�Y����[�؟{?w�k��=�7���Ck�9��t��x�c�د� [��uW��;�\^�V=�/��&���>�W�Zǟ���0��em>��o즂���z�u#.���3'��u�D�4��d:/؆ }�_!��	�� >9r�j{ƀ�t��㵇{Hr�oB���!~�_em��ϝ���I���S�%�O������0��AY�w�k,d.��&����{��]�y��
�'�����O�� �7�������Hc�{��k��gJ���'�,����L�N�#8�p3C�-L܍?:�򬱕c:N�6޴���=xF���ם��^6�Sg��C)�Y��r[y��M�S�$�~�>��3�G�;�-N��<A�r�4z��ɳ�_e�v�bO���-��ܼ�`I1мଡ�4�
���de���1%�'��TT�@7�����L[Ė��"��r_OI��sV���sC�g��bs�h�TO�g�������H���	��~Ȩ&�y���٩fΚ�$W�?=��ܮ���ޱ^���J~�9Մ�;���LYFo$wU�LSS�㥲�1 ���H�.+�k��sMq����W�GT��{�As���Җ�^�V�*�o� �1/pG�	`f_�N���=o_S�B^�=�Ky�Q�Y�[S}����BI��	���f����l=�bX�'�e��~�����=��+=�z�qo�����g�����[Ƴ���j��J��w]���ux�;�sƞ�|E�3�,���As�7��">����:��=���?��=��;���o�?��x��c����x`��R5P�N�,7p�Qў����]��f
b,B�ݲ�T������V�а��g_4�F9��[k�yl|W�"������'	�˟.&#de]t�ڮ���A��՛쵯�oiu*�Z�����Wݯ����rg7��o[�U�d���m^뼨�WjF��v���bpol��]�.���8��h"�=5}��A��S����쑃5(/�\���T
J�`�A�Y�U�{��,�J��X��ES�.���.���D=(u:����o8�1�n�
4��Jr��S{��Ul��obD��r���*��W�q,La��tC$C�,[�&����5�-�7:Nͪ)�ݝ��wK0�1�,Dq"9a��u�7n��jof��ew8H�e'7�n&��Ėx���m���p�ɞ��q��c�a�ǄʥqV�%MO�sG%���oBF���wO)�6��v�
�Or�f*�j��gt�yG��sOFP�[�[���G�^�,�e����D{	V�U��9NiM*�|N	K0в:}�˺c�mۼW���4^*�rO*Y3�񻕓qH ҷ�R{pwV��d+�@[�T�����J��4Чx���50�m��汧*�#hÒ���)�G��,�]x�KÏ�@jڭn���RQ2r�jS;��<.r$�U�lQ�K`�01pA9�Pc bŰ=A	@8�B��a���,X`z�1�P��`"��b�CF����xM	$�O	�+�"ة_`?04j/A��[�E����?2>y�+
Tǽ�ߌ댱�v���cR���
7={���#�)�ޕ7��U����[�+ږ�I��^<���S̵7�M��[t�ņ�1Lb���ʣ��q�Ns�:�MX�þ�R=B�����99�ɲw��.���9w.��u��Q����g%��m�u��b��YA\w�y�x'��ָGhF0�B�I����ŝ*��� �o��fV
,���5�t�8[����XX��eJ�+-%�s�	Y�ɼ���Cp��2-B��Y����|��Ղ����Wc�a��ظ����ڠ������{U��F�{y0)�3��җ�Y�t�k�P`��aO�T�*�ū��]X����h�Ȗe�X���n�h|�T�r��|K��N��̋'P��*���{.�9Ί����c.�^=8z�����s����\�"���=eʊ��Z"�]�j⭫�`[�29�4��w`�j��������.k�59��	Ƥ\�n��}j��e�N��hǱ���-Z�뮲��B�^q����+��>�e��cu=�g�l�wR���Vt˪t�:.2\����8�<X{rv�u������8A���&~�EB���T���:#"*�|6��6ݖۋiUm����F�M�!�vr�sEQSɉ��+y�f-����_>4���GN��O�3�jU�.-�j�F�ds�3F��Ŗٕ�aTT����=?�=ݟZnȩ�30c
���Q̠��V�sy��O<==>8t��vfQS5��AQQ]����c&6�k{&*��������l�ѳ�:{�Y�p�[e�r��)�
��h(��mZ�Y|�/O�6t��ӡ�LDGaŅCT�q��w8���2 ���]�?6p������ն�kʘMTIi�h(��H����>1>���qKm�gN�l��p�a�q��F�PSUEDQ�T5DY�IPZ�(9����$��!��� ��)�J���u9:���b��RgĞV����������[�L�gm\��I��]H�0��
��1�r:N��V$�>�! }q��:��y4�.����dl�����w���=_?O$��+��$g<Q;���9Y��^���a�;} |��G���ʎ�d�߼������p����K�+�F�󛒲<���tss��tëow�^w�������\��%N3mi��}��&���v�p���7s�
o
��NA�X���B�z�1�r'{�LN_�C���*���P��ޟ}���^�!�4���eN�ھ�<P����1�|�6����t����xX ����P�䍟�����w(����An0`;���s����p֫o���דLX�����+(z�b���������W"]̸�p^JśinOU�s@^@21�m�1�}Y]-��k�7��eFC��캚<�5�5��+�%��*����HnCK[
��60'_�Q�M�yB�ckPG'!��e*��[��n��|a��K�f����$�Z���b�q� �x��/hq�b��?� �=�׻��8�{R!������a)�x�����&�0��,_�n��7�7^�t�?9���r���\RS�h�ٕ�Fa�p����`��F�gJ9���Y_�4x��6nVz�potp�qR�Bꦝy�O�.�:p��ʣ'x�����i����
�}�Wj>�sq�z�
�c�FM� P`��� ��fA'7��;�b]	��%��[�
���qܑ<�j/��ˡ�b[e�4wb�5����vl�q���l��Ca�޹f��=6%�)�$[���R��=�`�̪�������(��-�?Y��������ͱ���`6��E6$�sBn�'�ɕt��K��1迄ƙ�S��M�u���b�	U� ��栝�k6Z>�^�݋!bfp�N��Hq����Ǌ[#[`n+�柹���fK8���J��e����ƫ�-�����|�(�+п��6z�?����g��C]��4�	�X�����B�c�-�_*���'9��	��0��[r{M��
yk�N#�#�V����Ѧ��`
L�����`�H�t�3O��߃5��q��+������TУ2�1�U�9�*崵<k��={�ɿ�}�?���x��z[B�b�|��
�8%S�,EX����;E��
_i�+�a"�)�i���pr�e�uxc
e�캬��עϬrK9�+]�͌;V4�k�a9Ů�dwNl�yPi8�J�%77�լaJ��]{;S#}yD\,�F$XW� �u׌`�_a������e�b\�Qn�ήV����ۅ��-�G�GO_CC9��zm��Ϯ�#�\a嗜~�F�0��[1H�22}� �@�]�N�B�V���,}�0����{
��_�LMȭ}O�㶞�L@'[��b���۴=�T�8�Q[���è����ʓ��`��;.����6�D9.'��4	�bӗ;B��|�e �:��kx������y�\+F)�@ӭ7�=A������A��G6��t�t <����V�JguK�E�]F>땰@�������VP0��.� �O���mi���_�5cUy1=�EmuÉor�R�~m�ފ����y��R�ç���f��%���<x0q#U84/ǹ�Z�f�}	�<�����z��Z�����Q<�|�)���]�C�f3�׭Iʣ���[<)o	^؎p�����H���6.�O�S�Q�:��И��:˹�:�,�0���O���N��35!6ޑ��ff�Ɲ�S���{�oXĕ��7f<Na���[�s�{���hq^�g���; ,�1b���h~Rk����|z4ŝ>5������س3��;��0�����JL��ϊ��{�m0Ny"qR���9ؤ-"`��\^��!V��v�%v���♔�f��m(4��c"m_&�d�ƻ���˕�=�����ԝ�4�j�(���P��f��nlu�v=qu�y&=ŷa�=%�ل��z��f�U4�̭��Ýx�T��.sk=��<@�� �y��T�<b6�'q��x�{\x�@FKs�4=x�3ۗ�#�@��8\k���	.އ[wj��T�Z]G���ѝ �_E��M%e���J ��E�sKV$���墯�+_�x�6�S��ԟ\�I��_u������ڸg����_X���^R"8]z�uU�j����S�m�xb�Y�c�B������ ?	��Ɔ�Ьt�O��3���*��^��@f��<�ӽ�lٵ����C3�w�}��Lב��_~�y쌕�ܭ��k�n�7��V��HKd��>j�@���+��㗌p�ϸ���1��r�{��5��@�vx=A�\8�����z�Fa6u�nN��J���Ne@�wU��B y64���Ͷ�����5�G!����l��ϠX���)���l�Z��g�L�>���~4����֫^W�=����d�'��TkV�"
��;_y��S�/�T0
㛥@vw)��㙶�T��x���Z�$����oD3�C������j���ȍ�:^���*����Ӭ�Z���C�zh�qLM���J��n�2j-��2^@�`|�P*����_`��9�4B��Ω���A��e�$�xӫ(��N��"�+a�󔘝*�8*�U�su��3��$:O�3/O��	 �+��p����ABԵ�޷ǐ"d��g��� &c�[z���&ԉi���l T�ݩp���+;�R�ym˄�v4���	�N��a~� x��B)��e�6�_1�5RԮ]w?l?p@irؓ�n�����-�AP#�a3����p�'�����|V�c��lܕ��y�-*��PO��S��zH"�d�j�jX��q4�������?��{�T{V̻�j����z��]����y��Mm)w���=Oޢ`�ܟZ����"�]���s��p�C�Ф>�v|�(��͔�������)���3|��y��A�:��b9n{P�_���L�kS?�������y>������#T�*��dZ�촚u���v�j��O�5}�<�m�	_����B��~t���Ϯ)�a�S�T�I�zN���s?�J�tO/��J;���v��Aʒ�*j�^�n�'hY͌_�c'��~���p�0M���ɴMı���{��<3�ƙ�1���Z�YL
��Rn��e�l��^���@t%Ʊ�a����)�|{OP!�R��d����$�Pmfc̎ X5�����J�����Z������LSsP��+�V,�ʈk;1��{pQew؞���
�f���Q��(� #�J)e<a�)R�5G￮}ߓ;�����`lk�����|Ϯ��YZ�*oʌhm�����܉]��(�(of=52����n�L,Y��:N��b�yV�k>jw=AOFU������>���u�_�="i?"���C2J5�k�F���=��,u�u`K'�����.%�eH*z�@����0qi��3�g���G�������)LGB��!����z����C}�/�BU]֐�t#�u#��p#��h�Z��m��ˌj�|�WO��]�}�<����\9\� ��`$��F���(�;����u�
z�����<�j�[|�v=zJ�w��Qo43w0}f�7��./J�!���=��P�1�<�4�J��zЩ��l�i��hI�o	b����g���V�і`��;�hmN��@�L���X��8�n�Ś5����	�}�=�$xS
���Ze�xY~`������fá�5��|���?/�~ �������y���|�Z�8��ԫ>4��;���0�V�m������e�y�����-om��J�maV�}~�d�I��`��00Xt�T�l)o�I��ΒjV�w�M���t�RZ�u��I�.����-VUMe����v\����0 0n*��U��m���i��k��Y��a�.V�R��R�K  ��#�T=�e�f�߷�����8pj	B����&��_1`�ˎy�_��K?RcI�v�K��J"|�ߞ�?�4�>H�d�Z�ʾ�n������-^�?�|O~���-�>??���jk����<�dI|z�Zv�;LS�e�f��;h�1�xzn��8��|r��XK�t�x 3
�U�W�����ہB_�`
��<4pq��1lSsv����W��7��Sb��r�V=}z�<Z���L��~U,
@����KU(�)�����%�S��z]����V���{/�-ܩk��]b��̇�%�!ݵ/��zod�7��O`
'�1�j1�M��9P	��;2#ŻŝJ
�K��
��n��+ k�v^�>��"�o��r��.��n����C{����ێ�[k�W�i�3�˟�>٤n�ܙ̘�/n��8�M����˟��g1��
���׭�#�X�BC�į
��Q0�����)=�Tsm@��,�~|���Ӝ��U��3].Nd��{^�q���yN@���@NS�4g�XT���V��a�"�|�Q{�{��m�w��hх�b�f��	)���]�B���t�f�T"����v�F���h�q�:�${P�q��lw�K6�W7UXý�X���n�v��{�9�eb<v�|�8L����i!\}]��4�-/9��:or>�F	$!�Wp�8��`�޳$�bV��o��e��"#yԿ�=v��w�)0�b�BQ��,%��h�nM7��B1<u�K���n�Z'�M?A� WKμ�G��K�*��o"�Q�Ñ��-�=�E2t�M�
��Ǟڙp�,�l�g�0�:� �Nvx	E�ï/��}֞��ݫ��z�9^�<����T�g�<��& z�0O�|�h�?��z��d�ZE�?���V>Oږ�T:{vK>HwhCT��qMr�O^��f�%��%E��ש�����%؟��z�T�[}����P�C�h�����Z7Zb�5�����}w�J��'�Y�6eh�om�Ab�����,#�o��J�K�����	V�Q���
��0{j���_�*�r�.�.=���;
�v�O�L�fij�%�4����;�S��Ɂ�U����iN¶?��`���̨
��Ǒ#:�#�V��o�G��Z��$�{�B���i�v��nR�]��������WB��_���e+�)�l�m/r�		�Ge�L����u���� ����.���&KY��cb�x��Q�vc9�ޅ��,�<˳��S�g3.��G X��,X��]X�2p+��H��H+��us�nV&PX��j�fp�v�Ǯ��7[��������N�OpB�#)���C�#����r�wA!8��O	��F��fX�!@V7d���|TY5"�a��X/����ևh��뎓����C�0��:�=]�%t.z��]R���
i�UͶP��"�!-_�s�3�3���	����r����Ш���2E@懺��w�R���1��Ǧm?6'���
����οq��ZA��j�f�<�ݱ�6<��xe4�����Њ�:^�F��QZ؜EN��fZ����l$Pq`�h.�@��~O,-7�y5�h:F��#[��Ԗ��KO�l�VG\ވ�pF%���K %�0N�8�n;���22�6Ʊ�������,?�֫�/Ƅ^��S�o�b�J���5�f"Yb�l�q���'�3�4ϻƦ hr �� ��}����&姛��)��;nP����Vg/��97�W���
�wI��T�Ƈ�Q$��;��r��+��q���>-�X()���ǆ)-�-��ߔ�Cop@ٚS4��Hha�	�$�ac��'�.�:�2�߁�l_�y�z\����W�(���ց��KG�y�>�(5nl��{�y�#VQ{�a`���j�Q���6�S�i+���uFn�O��<y/5?hJ��7�U-4�I�ѱ���c��,�RN&M�P�3b�Q�*�f��,������;��s�PG��h���� � %=B`H�B�B�B��0�{#	Z��)x��}�1���3������m�g�c��;v�u}���{�ʙ�����%�2�Ûz�����}ȝ��15@������~���T��Ix.V1���)�����\� A��T!��!O�}��O�x�T�i��G*HE�D��x� �����X�<�J��������I��{X�)��s�KU��z�Y1�q�F5��n�Ύ������|��C�_V��#�@f�q6�Zj��dέ�c����]>���Zʊ/ VWm-��}��m
�3&n�P"���Mp�@~�:W����\�v�bl��Jc@�㬜D�:�"��~A��s.뜇���K=��P8r�ٷ����5�
u���$J�5�=P�
(��Sĥ�^>�C��l��Ӗ!�7� ��d'�ف�L���`���B9~s�Λ��s'��:�d;u��-1[1���v���cO��jg\���:���t�1�������=�K�M#�Χ8Q<N�ɏ��UH9��X����+OU��I�j���Db꧹�΅��4��js�B�e�ǘ���ƛ˰�"��W	�WZ)�au�ee���l���Q��V�ޑ���'
�ԯ�s��3�vz�J����>��ˣ[�K�`H3����F��h��]:s���	3�9_>�:wp�B�J����wU��Mů�y���{8J�d��:�U��p�cz��ۓ�Ge�l)�H81=��ǯ�R��/336�p�����4�m�)�V���R�
��+��ԭ��@m`d^�v�֣W�՞Ь��Ӭ]Qг׮Ŋ:h���o�=y6�Չ��nʙ��m2�Nm��\�]���wwp$�3�,=r�ۑۻv�̱����t�Gr���jx��7�r��EU��n�M��`�I���]-�OJ(�
Z��J�w,��oQ�z��V�G��Ie��u!!����?,o	���hc���.f4��r]�(2ɝ��PW�;�YZ9���ɡ���,1�q�h��Z5��b�b�[G|6��D�1ߟ�Z�.5�2���|��e�j]f��N)�N�_w;���,�0��ٵ��!x��;����ĬR}k;pw'�bͥ٤Jw�,�)���]�f��Ѵ
�u��MEʹ'KR3�u]V/�����+�u"��qs��>��c��#%1�C>�A�� �4([����_!^�,Pv����A�	+i�����`"�� б���,b��q�: ��a��^�������g�X!����"��Y�h��__����4�.���9���}I;�핺��!%MaCs�Yo&a��-�ܮ��)[KK3���[׎��sZ���vd��("�끕�H��VZ�-FO.��-��B�0�kJ�;��(��v\��io	��Uki�{rn��e˺��w)'��y�]�״�;:�گQ�)V����tm�zńƜӏ��)[��+�K+�r�uv&�_N��M�T˕%	V�U�Uv�A��������H���]��W�q��d�Jw9�B�sf-W�
�f�&�Y�je}�B���!CD��]��og-����K{���6�r<}H�q�4GyeM��'
���1,�GR���r�a�5��Ml�f��B��b�!W:��/�!�C��wuޥ8����+�BU�3Q�5��n�Dù�i�����QD:r�.Nq/Of��
G���w��]�U[�	��"�qG�I\�K{Wj��棆N�S��vr�_a��ɨ��Q�k�eWm�Xƹ�9�Yu,�6�aoy�+V6���ʘ񽾳8����r(�Vm�W>̝ʮa�q��'e��3�_U������eJ����L���4�MxR״F]n,�uR�[����A\o*�Y3�I�b�G��9�ϧgwt"ƈ0hB�
b�l�Ҵ��J�Ui�X��m��Um[SmM��m��m��m����ѥi��Sm0ڂ(|B
&JJ�B�4(��D�F�T0�j\��&.?�	%���^�<��
��4���(�N�3(��f32�1""7=:|t�z�[RҬ�T��+BTUTQUĹPP�Æ6p�Ç��w��,��DIME-;�L\\Y�2����ZVWN�h���t��%Y���)*$��b�-�2&�Ģ�Z�:�A�g���[�--�*ڲ�m/S�������y�b�������=8t���l[�U����I����&����Im噇6zzp��n�2ǵ�5�5%��PU4S��UQir���8a�Ç����h*��j �L�"��ʫj��ڰ�N8p�����;FECAEPq��dT�q&J=F\NLQ�j4N�;�!����� 2��γP���2r� ��&���!ķIF@ZHZL �l����۸�}�Ȭ�::��e6�J��y���m]�yOї�Y�u�we:�܊"�Y���X#�h`�m�i6��UZ1T�dV�����l�Z�*�ձ��f{ ��Q�IJ"�
u�*I�RJPe�y��us����5����1��(�2�v���W�f���6�=��ז^��9�����v=Z	�-������o�Ws���CA�i�ѭ����%� �t�k㉌iN��vky3zY8��lF� �T �[�5�w0�W=�K�:p����ؾ,+h�3�XL�S hy�67ƴb��/�(P�4�gp���m��;�嶺"~y8���.$�3���� �x�@�Kd������^ͮ`�uf��]�b��"W<�R�$������C��� �p~��7qm��D��t�C�E�Ky��]�s�By~$������]7���s@���8���Ac��7T��G���������Y��E��Y��?A{b<A|������s�����:ho�X�ʜ[=O�{��n�!��A�H�����P�OL ���~a�u�&�E�]X^�z_)xPr���|5$;:���	Ȣ��Ѱl�?�}��p
���d�	�LC>���]�r��������ﮣ��\��6�'iP��Y	*���m�ڋ����	.�L���	��`��u�s��>wY��f�K����GJY��)��(w.�ụM*�^��;�An��gm�C]����=DZ��-�;\'q�6�j�1KYG�s�w%{�����
�4�%���m�e<�uUOF��� �N�����z�;�Q6�A`���$��
XH�7��������x�O���#am�ǫW�+ܲr^���#�����O+�DD8\���E)z9����}8�K�u��Ë�.}*=���o`�gvb�]�]<y���M�Ϙ4ps�=Y���@k@k�\嬘ze0�r��oLςe~Ҩ�Z�n&xsC><��m��m���[���0��؈�_`�^-,��N����V��'�b�Z���D<L���e�G��i/�4,�
��s~A����{)���F�P�=��W� �I��؛��zj����Z~�����CσZ`�O����cC~x�h"#�)#���0M�0�͈�[�]�Q��X��V����>y�� GlB�t�25�=1b]�o3�cR�@��_����>��u]��U�'9UkV�d���u\P�WN���	���\~���}b3j��+Y�_����z�L�nZμ<1�]0CC��/Ё�$(� w����zz�^q�{���cŅ�f�=�4�,OOs�'�H_>�AF�~[�6�h���t�.8w��`ӽ4�_@�.�	�T��̼�p��M�Zu`�_�尃bp�r�	��Õ��t+
�ӑkҮ�o
��,R�)�(��u�u�+������- ���T�H�\�kC6�&�r�y�R���M��o�7V�s#	΢�M]K�T����� G�� ň�,��RQ �C$U�<�;��= ��w�fv����zD9JMX��Ȍq�.4]�hiO���4�f��u��>Nr��������u�"}���S9�J��qz�����0�S��3���=8!Wb:������ӷѮ��!�z�^��̓f��Y�І���?��u��^u�uM���Pv1�;0��xc��[�U]
#�Cϭٗ;5�۽5����+���Z����`�nj�x�>d ��怀�2��cØ's�2�>f�m+�aK�r2�ȵ1C]À��8��D\�y9q��k�Q��@���+rD�(<�9�`� �L&��U�x���ͱ���(���k5w�ڄ1���"C0r d��+vt�	J.(�Q �Rk*9�v���A��NIyC��R��z��n0 ȹg�vlh�<1�Jy�M�4"�O3��jB&;'+m����ƺ�m��6�6�X��+@_���%7�?/f ��n�^H�c=Y�}O��|����	���v� �sr��0!cL�ey���v�Q�K>ެ7���eB��.�>g�'� ��XN���k*ܽ�[���z���mvJg`P��z�'tɫ"��ѹ�^pw�GG����匿{8s����ve)u�`��E6���8\�p�� �*�\�}G��:�j��>�!%��<���{�9�W�׹��
�}d0J���P�H� �J����.�������73��j��=Co#[�b��<�연T���D�`õǱ�z�k�cc�f�n�Ty����x�B]�~O8� ������������`7՞G5��/���	�
��p����j*'���'2|����7�e�5�a>aʊ�\؞����������#���:-9�
d�Z��Cm�40�wk�vg�`�DHv�GT�P�EEv���x �cv�v�e3�ښ[�K$pAU$�q�Sl�ܗ�P�R�`O0'��Q�o����3��q��6����M��'��eu��?� x
���ё��e�ި�p�N��F�=���)�G(�H;E�,���h�u�rq�i����P�Y7���%���-�z�$8�����{w��!��f�P��+�J���c��<qŵ)���\w<�[���,o���Ro�����6�k�~�ߤ  �uc��M��B��)@,c܁�6�/޼1�zX�z(�[��aUX�շ�߭�],�ڙ����2p�?�U���}�!�\H����g��V�Ď#����d''*%�L)�3n"*���Y؝S�HQ�\���[y�d�7N�=eR���]ߧ���7P�UA����ER3�0FXb$(���;��������ѳ�MrM����%��e�r�ˑ�L���el���r�y�5���.񐆽i�J�#Lb�q�Uc���m�5�5�wmH�X��P�,��$R��J$��
X@�`�2TG�ط��ͽz���8` ����"BRK�~�� �����_�
��~�E��e7��[!�Ju�Ә\��Z��f��$�<�;.Ȋ�[��֕f�{lI��#�Dpz��Ĩ֘~�)�<�V�KL�0��k9ݐ�d3� t8��T�>��G,W�ƻ�>0�����ι�o8�8�a�������>����;}X���:�j&�q`8�,�{V4Ke��D��ݱ.�ز���P�T�܅�R�n��?4^�Z��e��������������l�?�c�d��)õ�۝~Ĩo���<�~,��縫�}��N2�dSH��Af1�٫��Y�����h�ă���TUo�P?:���=x�D�Ӑ�2z�UCLT�Л���(���ψ�|��H��5�Ɗ�a���;>=�܇,��;�s&`;��<6�ood��y����|�� ���=�x����2�+�Y��`�K�����ua�0е�u�I�uN��\߃���"� �����'�Y�������\�!�:<�tN�;�ڜVS��yfd����}���O����p˥�����ͪ�lY�ʼ:���_�S�\D����rtu����[Exp@ t%W�-�k�m�T3�uμ5��̾���2��݆��D��;��<����f]�Ϲu?���* �E<�C�E�K�Qp$U��,�j�L)5b	C�f٨������/V�ڮ� o��Dp�,E`o�����x|3~]-�8�Ão@�<wgnU��^�ÿ9B#����&�_�1\
�OP�����j�Ƈ����QY���:3���~U�������"�f�E�!�o���yj�<ۇ�u�)�\�@A�r����H��O9Ǘ�k������<��c��[^�o">�x�@0�|gd�v9f�Qm��z�����gZ,�Ug@]K�2 2FVؼzz��6=��-�����HvC"э>d؂wAZ��x��P�0��\3Y|��~rލ�:��=��T2:<..(.�����RV8ʾ�Y��$@��r<�`����nc�t =�|� �Hy�8�}������,��h�Y�E�oJ�� w)��Y����y{����/�#+�8�Ӛ�BzF�G*6 q���b�bzC��\�ݙ˹���[+|w�!ųC;�u��ܧ�m#"O�O��)�*E�M���b���Ъy@��t({hf�$�}�1�|WK_��T�<42|�ov����
�4�:�:�lv�bF�{�\6��<S��`͕婼s.ԯ:�w�w{,?z���玎��$Mf�X���>�]����'2p�W,�7T�tZ3�n���c���zN��y�Nd�쬳,�	��yp<���H��@��AK!
YR�IJ�)Q,}�xYs$�ރ#��
;�4Q����n/M�y`D91���
|u�!��{�Ƌ�]sH^�M��`¦��^��?@#�_�CW���X�Uy�ނ�	`g�&�]�՜�ܠ�<��S�ԺN����xckH�k�z��g���g,;�v1�gzx�9�H�(#ɕ��t=���`���[d�=�҃^H����NG �k6�6I�^���A���;����K �*�A��ہ�4;^N�ި4����sx	��fv�k�a�I@�{7ô�Z�E�������~�؀'/��WU�f��-��ͺf�5�7�:g��-��3����{$���E@�)�������X�{;t���ʸ�
���c�������%d�6l.�,�B4
e�pͱܕ��n8��3�D��8���L��Ķ�����WV�	jfS$��}�Kt��Y�7��]l����Hݸ��4�C�MX�xmx��LrǑ�ܧ��M���=�ɛ��>9se�k�JɛY�А>�R-�{�c@���G$HJ=y.�x��ݼ($���߻&^RHG^g��_I���>�e�x�z��9Ӳk��a�����Xʝ|pqb���FY��� �΢M�M"�ޛ�� �	�暪a�V���g��G�91����ܯy����Kt��ͩ�i<�0e1�s�X���;7�G|n��)}�
���VD�j�0��H��L�&I,� ���� �5K��-�5�O��$T�[�(\��?�;�|fy�Z�gny�N^���~�Hc�r��-������aݭ�tC��xcP��`o�dB��F~?�t����~z��_��$Oy��?yF��6���i��):CY�#��[o��FΊ������\��}��B�r�i㊊cÛ��0�fƈ�$��s_�@Hz�� ����ۄ3Fb�,�3����C.�*yU��<��Ц{���VOd8=�~��A�-o����#{��gjhۇ�5�kЗM��y@��'yV� �3q������a<v)3pG	^�����@��Quu!0vH��HQx	��8T:��cPKߔ��<�6��s��fo^�.:���z���Y!Z�Y�c�>�~��X�;����:�c�	V6�{;U:V ��� ��
u�C�KL&rd,�?~���yN_��S�ݾ�z��4z'$^����#��|g{]q<x����RPXH(Z��f?���8:��?�5������i��O�Hr*a\�'����s;r}�ٲ�P%F/�F�.��F�_E�W���5Z��PuI4]�ƱAJ1(�@��-�M������Z�9�EZ��H�R�L��ܴ;,Ts���A�q���p�T&�a� �� � �ژ��mX�La��6�e�Fk��kXZ����o��}�"�U*A��ȉ�L(�R��J�%(�Y 5�q�߹�߷7?UK�|��ARE���#�??�qL6Gl�<:�;Dj��^��[(�� QQ�>.����ŽU�.X�"i�U\�B��ګElB2E5� T��e@���]�"�=�K7�j�l�*�)� D�+��k�ިCNC4�Ks����@ML0�g4��X��Ȣ���P�����b�;ì�/L�v�N�,g��Y�,�${���@�A��Z�X�� ȳ#`\�:�5Sv�\j���xԾR�B��B�^0��xi��z;<<¸��0�*|�ٲ�9�l�hR4��h�N���;��s��zf��o��eF�f	�PW����~	ׇجY���'-�}#�Q���xgZS������jne��(���2ak������5^P�sw�����dh4�XE����3K5Lu�F#
���7�*|nT6D��j
�=�r�h���Qx����[+��31�w�P*����j<���;�7�a�w�n���1������^��9�����gg�@���3yI)��&U��	]��u�������=`�9.Z����ڌHǤ�dn�N/{P0�{���J��6�������̋S�R���x��8��y��5�R����s��ω�̖ފV-��a�X#�Y�T��j�O8�k,>B��|ڬͺ�{�	�*����yF{#�:vq��|gV��κ9;�ԝÉ.�۽g|��;����#TI��D�X�)a�C
�,p���7���\O%��!S�D�:��r�c０��"�I�
�/�'?1p[�\x����U�k��Oz�Go-�2uO"J +�=�2X[���vl2kèϏ|�!�,i�I���Yn�MQf��)O�Q���y�i�*MaDKE��|ڸoH֗������0�軥�ӫ@�
ji{�U���{�b�&Ic��ߪ{����?��O���-��$��5�����}f���`<�a�ty�C@��="[EC��dr�$=�V�1�����g�0��jľ��AI_��z-��B~�����y��ǐ59�i�;&�6c�3:�70i(A*���ۘ����e�k���+��}^��{c�S�=��nE��zݲ��"�Ύ��:���U~B���E����P��,�6��]� NY���
��<����'����7�`@�>��Ǌ:ؼ{Ux(7,���|w���g(ƬJ���Sr��޾)K����4 ���j{+]ۜ7��k�*} m#v7��`6��8k|��x{��җ�����^k����Ȇ��܍��S�&p,T����	:��F��T��fU�!�Tʛ!v��k���#�،_�H��׫���������=]��4�v�H2"P�F��pr�G0
�/���f)�Y6 ۤ�s�(�F�vv�fЏ:�w}�C���=p�JnQ��Zp�/c�kUM=���ጉ_c�U��f��5s��Kjh�|�R�s)]�b۶���6�}/��j��5_(t��c�D=f���,嶧�<v.\��"��:�ugD�u�&P�v1%��*��.Κ*��q+u	}���]���p�����7+DF��UǮ^�\ı�|IgQ�`Յ(�J{hDJ�p�]Ppu�Ъc��g5Yz����{**l�G"��u܏N�Ϊ��Т�����{;�8�����e�Y��E�`�6�ٕ+i�k����r4'fwE��`r��N�����v-ۡ�X�����j��c����|�e��Ψ��O*�������0b\�*��Q�[�\���]ڮ���:�9d�\ؾX���J���mF�e㸃�F��	yҺ����������v���޷sT�:��p�f���}#�ʫ|��cX�Z����M�9�왍D�[���瓘2'�Ҳ�J�;z�p��c29��A�M3ՇvA^��
����	b�I�,4�*�(6����1��q��x�OsOt����z�y�ך=��
gff�>�i������[ӬyW�9�=x�ҕ�� �f�,���,+}c�ڰ*�����X,%�{��\�:�����]b��]�3�9V[:z�׊�i�����
m���5�^��4���]������γ[yL���x�������Rŉ]��Ke�et|�.ggVrZ����,��L\�77u�Ǔ�e;�p�Սj�[EO�;�[����I�AxQB�@���sڂ�Y��.n�Y��S�Wկ�\mT��i}֖EPf�$��ma�3U�ݡf�+��L���`Ӵ�M�W�w*iv++.�G|����pUR_{-��ҋb�غD��V.��1��
����Ŭ�Q����1'd@�kfWo�Z��FG�ʏe���.��t��A��9�Ϸ,�ٌ[Q�ڻܭ�)�Gyߘ�vb�[��1�s6W:��]������s��U)9��V���ݼ�L�k��Z���T���[�ʖK�JYƻo�/�Dj)�^�8y�ƅ�ia6�&a}1%b��m�9�^^�V�Y�2QS����u.(`�5q<�yS�9p���M�p�Ú������Vn�"��I�����d��4$�SVMC����i�/y>�C$[/��er�����B
1=�3R�=��$y������2��O�pHo��4�Stt6p�����X��d�b�l�K4���*����5�ﭡ�&�m��p���������VIA�8AK��30SBE��+,U�ץ:l��ӧO>�FEB�ӱKM!�8W�Kc�]bj���t�M�=>:�*q;�������Z�X˖UV�W0^p���Ӈ�R�e�l�Դ�hz��uU#ERQ�lt��pA�qR�!AKUAB��ذꋷ�qEFMZU&�~4~8z~?OjԵ�ah��o��)�%�{Mѻ*���4x|zp�����%J� .�44��4P�CkrB��UC�UC����V=���AS�����,���D�L�zԺ[p[��/K+OG��Z�:���[�ˌ�����3���y���B?�D�Y��
T�R��!��)R%(���x5�E2hdߡ���y�:h� 2"��a��-z#��2���)X�����p��_'[����Ɔr�ǔ����[5�Bwc#����teDk	'gY�{Q�V7�������1MƿkI?���$X��Ƒ�K�m�ߗ��ҁ7�x�ḡ�:�2�M)�Ts�:ޅ�2Ҙ��S� �7G@���7��n��^M���!�`�&.b�91wQy����(@` 7��
P��L�\�g�,{.lCZxűj.���>H�=�w��1w�B7��SV��u������
^+�	��T	�ky��/>�A0p�"AV$6��v�ˤͦ&qF>Xi�[�חl8	�\�%�>�,+>��|0�(ݔ7��q0~���(�SC�[�10��*[{�Bǰ��ξ������=��~Y�Z��h�������F�x0��L�EL�[�Fq�����Wލj�&r|
��+���T���x ��!��gc�dc�aUܵ�U��kcW�;���]x�D��L� W�F;�<hD}�1N���#[ߣL2�-����C�A����=U��M]��S���b0�&�_a�t֞���ٯT�'�Sz�f�r�'�٬���q�0��b�_h����[�?�cIPYp�׊��+��F�^�Z/0U�|��׾y��x�{��o;?�I�,�����*�`K�J��`� � B�Ԏ����^����=���օ���t+=�����+6O(��%��z#�W�Tե��\��L�;��U�mz׆G|8�7����`��ٙs�U:ܕt��5��[�sg `�:�� ���^� ��
F�K
؉c��S
!�����<��h/�l����;G�4�]�}���Z��c`����,�<��Q�^S�
T�����[l]��r�#������ΐ3U����̝�}�'� �n�t�k�� z#��q�!�ԩk���Ķ^)��ZzSu�R��O�|��c�I����|��_�>��~��Sz�;&y�R�s��^�="	��J�~�h�����.I��}��#���
C�#0������U�/�3b�H�����^*9��)�u�L��ۃ`hf[ٶ�ǦA�5b�$�.���JE���Њ+9Х����9������y��q�iZ�O��0ҝ�F�(͛Xڵ����Hy��ׇ��a�z��>ϣXX�����>�Bn��������+�]�G��\������)[{���L<[�D�z�N���zUj���8cTB*q}w�)��[4r>æV�`"�����`�`��]��X��5��a5���Yܷ75>Fgy�x/�R�s{�
~��ӱ6�2�ܣ�hf��8B���S��7��C�*
X�XabJT$\�!X!H W6�-u��u�~ݯ�
CE�j��V���b�I��� k=�P���g���@�鿠�y�8i.�a����U`���L��~'��Ykh߫���|�ȱ,�|F�s������ͬ�f�|�e&-�s�=�}�D�r��`���NB��Q�W(��Q�g�xia���j];���pVg]�A��'�ȵ�B��<��v�hئ'��R�&{*�J�N�6�h��O�Q5d>p�±��O[6�W�P��Rvo	�RY���N9�a�b�#�� 2%;�*�}�q�1ɰ+���UW�@g�ZՏ/���`�y^1=1���B7�n�-˶i=��bX1�Aݖ9�u^�	��9c�U�Z|}����JV���ո;Ke����&���-9-:G��R�R[>����r���,��rP�﯇��>u�=����W(0���3��!>7��z��� �'U���M�֐�ɇ:����8�*e+'p+�ƭ{���J���o��/�me�Fu��#�S�q��c]R1z运hE�{�zD ���w��3��ޫ�tt�'y�~��W1���տV'�����X_d^�Z��YRfI��h�[�z�@�Yю��r�>*nV�]�>b���fL�47�|��KD�
�a�oXK����JA���p仙os����*?��)��0$H%`�x�>�wǞ���
����'z��*��R6����<SyXS�Ӿ�� Y���>�^.����wѫ_��(<"�ő��֠KH���u��?�b�Đ-g������*܊�۩�@W<��4��}�]�}h�2*���^�ܞ�����|Ѝ�Ҿ�y������}�$��g �
� �406:-�H΁̎.3���§E��w�з���ˌ2V7��nj�������� �큲��7 f�V�W)���\�w}���8ֆ3�r� KydG=7 ʽ3%����׺ ;�7�D��d��Dd_Hz�b
�=RJ����/|�X����f!��;��Z��~���{[kq|��`��jJ)�'�"Z<���k��5��kU�+����B����� F����57�k�=q/�i�H|4w�]}�.^/�z&�s8#�<�2��]�IĈ��`D�4(�!�/�3�Q`o����DKe1�##�e=�$;��x�|بp���x��\�ߕ��n��������Ze�%�nCt>^Ul��
�}8qdH�˷�JJ5�Bꦣvn��{^���y2��a�K/;�o��q ޲p@�묕��+V���0���ǹn�W@��5��P4��O/^kw�_ob��J�=�*�<�&U����p��eB��K�z׽���_ሥ��4QJJY% 0 x��	Q)kf-i�ۡYΈg��� .H�%�ҳ`���֟A_���c�n��%�jkk�)�ZF�X� ����_جsc��LȀ���d(�����;05�!*��ߠς�ٸO���~~�X���1���X(��>(��V�(W*��N=�zw��D2�A�ze�sUF�-sxC�ٸ4
0�(:�6c��yeϥG�OUBL�LvA�<����)j��D��`�7��d���s;hc��9k&�ƙL&��~y�ˆ���Mҧ�ZoIv�T�F�44���f
��x D@�5��8q����;�"����e�,-�/�M�ѫԍ�!W�������k�F��ԟ�-l��ޡ>m�����h��.\B\-�Z���J�vq:�c�Ԇ	���0���*u���SO�=���|WK�~�>�BG���mS�v�t���y!��S��\�^��M�f��hkO�-^.��ʆ�ir�<Y�Fs�`�	�{�[*r�+2��4z#5o�&��oM+ʄ������f���9>������ݭ�ϓF������i�l���K/캘h��y��wZ�fW��*�㮥y8�hPN�c�={'T˕������,�A�e��r6������,�<flW�Ǯ���V����ٙZ�?�=� ��G��Ly0�$��#�u�;Mz6�����Z�~�y�p=#� �����"e�u�&~��v;�9~�4ww�m̀ak�>=Ј�C%"&L�B����	�0K�@Hw�Kŉ�������E�m��9]���xwzX��:�@�����J�uECTU."�D����Y��������,͏�b{L-(svC�,2�4���n<��׃"}��������O�N�~L�2�~�����Wv�F�I��,ϷC���	�{z�V+�Pg���*K��
H�3�6�W+��7PU���?���ͪ�>�^�i��5������7����w�j!�&ݛS��˖��W^+�M����ml�y���y�9������S��$�i�Vw����'N�������Yu\_�xED� �*�%�\�-m�CE���}���Sw{�Tˀ��{;�m� k�d[s ����5�,��%O��@ɨ�v��R��ƙ����Qt���&mWN�C��tĿ6�R���8G����`xSG��j8�����y}H4�3�!j�)Ȃ¤q溷:3;tj㔶�:-\�i;륐!+78ö#�K�:�V���ܗW٢�¦'�m6A��Z�b��B^��}�L�Gkv��&�б8.}�V�pv�KqeR��������}/���_m��x �� ������`(9��R���<�+E싅R�JZf0�KB��򘺥��V��4�1�K37�LG��y��˨E%:����*ʚ�~pSsQw�#ѐ:����������O�NV��ݶȗ��b���/S�d�H����<�1��?7,��"_detm���2{�0����ý'��o��[�+}��������ī�xk&ʸ��f|�88�u��T����� a��f���0aj�c6���%������gB����g�χ&�}�v?J����ɽ��������D���hO����ς��E�,"΢�t����x<��J&Ȕ���3�����pD������%p����@8�%�*(c�esz�o+%r��`��r6��=�:�8HFo�@�t�.-.8TY_52����x!!�ɹ;*�LY��5�۹d�Z�;Bޯ���~�"(�z�
��C�;�V�yi�xl��r�1��0E(����/��7��>~��A*�Xl�@W�#L3<R���i���a<b�"��/�#�6���K*�	P�������UE�H������.+�F�
}7��^ug��z$f�UV����,W�\Pv���ҭs��R�v�6�>���M��V�F�rO&�V�s\<���7���������������q��#Çtլ2T�w���,�X�'rϭ8�h,tLS:5{wmfT轟���a�k0�*���{���}��~')~{��lƙ���8�p�� K�AC�L��6}�ކ9c�3L���o9���������y�%"�(7�lVD6��}uQ�����$�m�4
{a��q'f���^>��V#.:6;	��b���zȇ�m��>���".�"�P~~��f�I�$_��wN����R��kf�(�w����ef�l�a�ⷀh��Z�gD>3�r4F�-�胫Yz�&�c��SƝ���+��gȨ���
�P`3�c����/�u6���t�y��"y�	���2�glj 9Q��Ů�s�/OV=Y��X{���`�w��� �Z	6D��S��Kͺ/t��W���(��m�д,��m��X�T�T/J��u�ݍR�vN⠑��~�/��dj����ʺ�ڄxv6#���ĺE�����*�V��v||H��4E`�O��O��0[��K�f�j�p[B��z%{�Ԩ-w�X�澰&��y�;Z+�f i�� �Y��s҆�@������D�D�c��xn������7�l�'�e��x2��st4Z5|Q�� �@��$Ah.�}�;�7��sw�[N���*�{߳V�[�Ե#�>�jt���z�܄c�,.���ŎW���@$` 3 �彉s�����lmټ-���gE�S?�pC$刢%Æi�t�<� #VH��%�#���lv!S�C���y��� q�����J�����ݷY�9���������Z;�0����ge�ӽ�q� �)�K�x8��.�tڗh�:gh=1�aG`��4Q�j�<���)��&"���8�OͲ~�% ������PS�J)�p�hRT�w(�U�]�qg$6[������A�Y~]X���!�ê�h{k�Aw�44�PSł�$tn�����m�c���p���G�*��q�7Hrl;"��0�־�o/��kqr�P5�4�[cNB�>�R[-i�qo&��*�}J��Y9/B��4Λҭ��=�����u�Uφ5d��3ϸd�\�'8�+[�<����$�}!x	pd�9c}s��| *�o�׵ÿ:���c��Qqx�p?��'P��04�`����t��Ϯ*q;�&�nd�����f��Y������3�� T�$>�c��U�Lַ�`��}��V*��o��UG>$�)"i�w'�ʐsg.]��y���@m����ܶSmU�eu��5W�qkC]LP�zaU�s��(0ӎW���R�����3t1�XVH��m+�k�H�1Ĭ��!oY�ÝR��[I�}L.�
����� � _ ���G��������+�1�⤲�1<�Bئ�C�Rm�����B�gߗE��������|�Q�u�6ل<T���@��q�⤰Z��]� ��i`�a�i}!K`I�jݲ͙���BF��$�:���zF"�e�0nE�RMi�h�w� �ʰ˫z}3��ԏ���4�	��zkP]Ct����W�O�ƈ7���@O0ǽ#��������b5%l�0��@�Q�i��d�~ �tX��*��}I�J��_����6X��g+����W�2*Zg��Ŗ������<��ck\���C>�n�o�/ፁk�m�Ssg��g
6�rh~���f�Q��j%�m��~��}���� ��Z�<�P�ߝ�H�'\��Y���@�oi�Ci�Y�����]2&�!a��L�?�6����L=�.j�7-.l�RQMk�ޱ�C��qh#7"qѷ�F+���sӽ�5�]3Z_���~��zC�|����h�3�؝�j��&� |ORR���X��U�~�[s� �=�􁽘�͟_�}U�"���wiY�� �T��#���$�uiٽع��'����c0�a FWp�BEt��N�;����20q��nh{��uI[��>��Ԓ��E�ɘL�+qf��x�V�<�
�}V�9�_p�yrlƩ��t�Z����(M/C#�BQ7גl���$�R���*yt�	h�y�n�ެ���g�%$!]RDn�%W��V��ّv:���U���U�yag��97�%�Koq[<&��<�k%�t`�ڻ�g��ܘ^E�`�fA�$�����tB�=��΋�V�ɏ[�U$�d���\��d��1=���wT�q2�N�'�l��5Uh��봠s��B%����4�ӻ���.Y-�Yt* �x�N˭$��2*���"��T,R:v�Y����Ʃ�u�.�̬oQ����0x�@���uP�9Ju��;�L�O\�����x�������r�8�>1-�����YLSOΜ�p��;���uxc�Q�vj��1�=����!z�yGr���I�3��Zܨk���M\�<�^z���uATB7�p=)ų:����E��֨F�b�hd��7(ud��&�Y���|+[���2���y�$v�Qa�>�&��}���i�+��^�יm�);��ˤ'l�B�f��qi��<RvZe_Hr���Dp��ӝ�0��4��p6����H~dX��ABCA���f�� d6�7z��o14�Qb2L�`��J�X�(X��?��b� �����9�c��L���)AP:ҁ(#ot1B(Xߴ]�a�e��lA��{Ś�f����)�+6�̮s�-�%��Rn���i]�\8S�P�]ci��إӇ
D��{�ҳ�gC�Uvt�S����8����/y�m��g6�l%��L���q�����N�,oc����	2�RX6漼hu�έs�q1��b�f9��伲��o���3$��kYތKmV��vO3{��N�w&JcGM�q��@����jӭ�(h��;+��g>��;��w��Z��w�x�XWܧ��R�Wk����$�1��7M��je��qTe��J�l�^�諭wZ}-��G}�
��[ns{�ņ:�h��n��ĩLhTÎ�:��Ps�u��OvsTe�4�Naɉ�3˓�1J��f{���k:�Z��̆�-5��S]��U���3�R]P.,~�\uo-��pV�1��b7(�G��]q�5�n�d�KZ�P]Qڳ�'Jwlo*�䮂���;Vr����G,�j�uZ�0���=�˵®�qv�sd���͚&��wWP�yq�YNv�����f�9n<�Z䱍�C�K��R���Ӷ'ϱ�&*�����k����(p`� !�1[M���iZi�)�4�G��x�J�1�+a�6���V�6�cF*����1�W�1ZSM��UV+m�i�l�����H��"E|���q[k⊇�՟���i�!��Ym8a� �
&�m��f���
�3	��MC
�Y2�Y\[cF�ON�>��,KK��%X�H���l[�çO:|O�߬Ci��.`u$@�a\˼���çN�8p���S�e�T{R=���jj��#�0�ç�>��Ų-��j���Z-�Iih�
aÇ����G%9�h@e���bE*��"e�ښ�M]S/Jaӧ��3�o�il%�qS�2�T��G��*�ʑ�M=<>;Ð:����5!AM--W��Ҥ�(���8|5Q��,�d��jH���&I���I�!h��rH���w���h��\��6e�*W�^,���\�V���۪���]���NhJ����aUt��Ž�|fH���ʾ�,mǭ4��1�j�&+Sma��0���Y�8�"fjܗ���i���e5���U����0 !0P!!M���.���W�%F�w+����c�⸇���}��HJ�6f��S�ٯ*��D��R�^Fcb�c���1�س���a%8�P��%�×L�]�xI���iO�<����4����;�UX?��,[	*} ?>��V쇮�:��w��'�{���p��3�����9�(V�М;�+i��0&!��Ѱ���mS*,L���UZ��7!jKzEY�b�r�l�s��z	E�5 z�=K������j�
�`�Cj�\�)m��Z�إ�-��e��H����5[�TW������
���|̱E�������B�v�M����Ѡ'����5�Ʀ��_�Pw��O��+;��~RFb
��o6Ԅ��$;G�(�B�Ϗ���>����GG���7�]�[Z���80��g���}���������C��!F���g����s}w��{���f�m�X�wZ��dR��_��ƀ�pD�h�Tg��S: 8v��~i��%D�op���=k8�6���5�Oe���Ts&�A��;~˱������;�%���)��T�f�Rus;/Mt��b�6ǄB��E���;0t�̡�,t ��԰�V2�]yJi�Ί�r������Q�l�uX�%z���'�5O��~������@���ΔX��l�3��C�b�8 H�z_��:��r�i�3������zȇ�{:�5��x{kՔy4��t��!��Hj��� �q瑽u�s�i��4��;x�l�uH<�z�M1���j=4���_;3�C�n�̟y�B9P��c��������o7Z�j�ߛo��-�����E�d���Lבz�r<�(����Ť���mh�7j-�ܶ�͜�w��^O�yW��U�1�g }�/�ݪ^�"�π��ރ��,(k��$�k��~W�_\t�5�O>��99Z�%Vk�b�v�we���Ҧ��d�n��0�F��Y]�����Ɂ���6?����\!Ӳ��t�s�Ԩ^P+kW+���}/ۆ����3ٮ8�j}�N�ӏs��f�r�=3��u�q�F(�Ry7���c��'�pIc���p]���v�g�6���i�!�&vMb���}|��i��ۣ�EE����R��(]��|8�8��wYwP�4��H�΋�LT��<�0���]���&L����!�m5�#�a�fͽ̞˺�Y+#��k��#k��w�)[��S�
4��Md���qЮ��n��jqY�/�d��Y����U��U秅�n=]��]֤�Ĺ`��Y�k�]�T�t�ϊʠ)Wd�x(_���f���v 3�O��~ߧw��SD��y�A�����g����yXU���c ���5}�S0��'�_����r�u?��3�J9��=?�36��CG�����a�>��җ��cSK�D�":;$��9n��'c�E�����^�i�;��D-"m����_�v��O���&B�z#����CY��yռ�1���z�H���������M�g��T�¿8�vj+HB��V~�}��U�}.e���Q�SX���\Д��hO \�p�N��Z&h��m��wX|�=���O��;=�\��t��]�~<I�����UmQ�U���Zg�Ft�L�>8���MG?1o�&e�F�1�/��Z�Tf�[Yf�5kF(��D�۾����a�3�[K�Gߠ��y������ibXF)|����niZ�5��78�]2�q��e��aM��!�w��w�E`�>��^�]xW~�G	�X����r�wE��K�qѵ)�2e�;qI�g8=�Eۊ1�n ���֩����Cve�����<�UVc�f�}�@qW4�Ƚ�GjE�b�v8ɮ���b���c
�����=�z�[ה���b�"0,x�ι�r�+V^���V�+6VʮS�ާr�Prb4�r�kVk�N8��n��ΐv]�p�o�� H��`0����V����C��q�4��k����
؊O��J���sP�7W=.Ӝ��k*vWV'��3E�" &m�q6T�P�M�.�]�':���b�s�Q�b��s��^�4�qռ�83���?��������֑�A;64�49פ�Y�#zS	0[y�8��<�q��Q�r�� vSm%+P�`^Z��1�~ 8>ԇ���?x�M�jR%Q¢xj�Qîi^�I��)���+���)������̙��;k�a7�h�p��LE�H�_�b�%��ot?8�~.�1ύ��}�/Od��� ���L�<���vQ�t'�b�/���cd��43�� 78y �?P�����ă�g~�Z��Yw�XB�b�=䇟s�c	����>��E�C~B�_���yO���a��)%�3.�=�RP�8���MO�ނ ٜ���H�
�K��(I�#�D#)ѕ~��}R�C���V�_����O�ɦk��52�~�����T�qBr
z�lq���� ��5��
�����c?':�독��J"�A�S��n�^�����z�0r��s�W�.&o^�C;q%w+�[L���Bp�qU�CQլ��gr�T䏏>ڍ!+%q�qw;'��B�}�v�)�L^!�ă�5@ ���� Ҙ�5n�{kY��f����i*���,w������@�@��YkOߧ�$��(p�~����@{��/�	3���T���Y�Ru�`�n�]˩�i^���@��=ρ�w.o������Pهc>���Κ�����D�Qћ���F��l�hq����L�!��d&'�Ь}��j"��N��i���ݎ���-vy֟�ax|Q��~\^�N��w�Z���oa*��� �=�b,��2h�����x*%+*��E�>�h .5<ǏD9�O��U���پʦ,�d�>;yEWp��Z�u�V0���ƽN��At�-h,W�O��ϷUs��숇Z�z�x2�}l���gz��g��3Y\~ ��g������K��2ۢ!�� U���Q����o��U�>=I�k����J��0�ǠV��_[xk�M�ɣɟ=���,g�V��'Ā��U�����hES����`�Ǣ�ۘ�;�l r][K7l�C�r�ڃ�r�*�^��P�a7��3ݖdKM-�e��(���; �τdb�*N�{ɡ�KpJ
��S��4�q��f�qA��f�>�="	�ɷYݙ���T�vh�����s�f�u�*�������4���-�����t���.���2�6�c��5���V�fZ�\O4���;E�4��y?���9��Z-53�}���?{z&��o�/˹|?�N_�,��oJ47���џK��������i��\��E�D����=���X�O͆ �g`TdkmOG0�"�fsU��$B�5w@~Bz��!���3�f���v��=j�?�������E�ԝ�j��}}��9|���w%�.�
��g �@haCn�'X?X�w�Π)/�G��S����d�,vbP����\�q����p��/����~U��&`�
��ח~)���kn��l��x�=�M吉�d�d�v�wނ�����DFCǠ�U�\�s��a��V�h��ڭ�h�� �0�B����(=������N?��*)�JS��f}P[�����[4
��w^y��&������#���Z���$縴��Rށ��jQM�"܆-Ӗ��_Ö��Ͼ)��é�MH�=�VU�~��3� V�t�q �V�>� K�BⓌl��~Ȼ�Db�W��5M���\��s�@�Ru~["@���9�V�*k[�-@FC���l�K�[X*F4�= �O�=�M��wsBk �()���F��YD���uS�jcV�Sn|�^�w�VѺ�I�:%Y��d�X��
�]��%�XuK�a.8僶���.�cHkT�2�}C�\�R[]�*ꖇ+
=#���}�_}� � ����@�մ8�K����(ư¸{����Jx�^P+kr��|����Pg�m7\L�J*�v�Z��1k�.�R�;*��9)�q��w�����*�P�P)����I���EK�a_�V?�_�ߔd>��Ҿ<����+�#0/U
م���Ȩ�ʧ��)�t�G��n�d"B�T;�a�Oq�@d��xjn75ͨ�+�y��&d��h�կ�o�]���Ђ����'�e�|�PF��g�Yߞ�ʢ�_�����P��Q��J��XbPX�����w���5K���M?O��Y��|j!�Cj�F;�Ȅx�"�P�D��e��Fu���Nw���ȃ����}��vd�L��-'�^�u�98j�4����g�* j��F�cPd��&9����T���ֹ�p�]�òhǼ��Kd������G(��˹ �I��B\�#����9�oR���]�Υ�~��
����ÿ�����]у�Ɖ1�{@�²b�r�uZ�<�x�X�U��kvpS��s�*ƌ��ga�z����^��n���W���9`Ёl�s;���p���LQ�]N�8�U�O+�rY\��u�O.u��T2�s���C�5������l�ĩVtgRS=��  ���Á �K8��j�0@w��nP0oJk�_����@�Y��A<OB^�ŵ]�پ�*������\'�i}��}޽D���ˣ �LC^�#7u�д����C����*��["�>�B�n�=;��(��Y�����	�����k�e5�ZAn7B����hg덩�SGaVn����j�~^��s���ҽ�V~t���~u���o�E͌;Ck�Nc�œ(X!��r��C.���Уn�D�V��S�;,p��h�����2 ��c�r�oF�Gբs���y�-�K����ip3�cd9m�����4%^�c����\��T���b�ں�ۣvt���3g.�A�ީ��,:��D�lgn���M��x؋���|f�b �T�����\]�se����e��6IRq�BR���
�fb^L@-��y.�kB�9����w�A��O����#������x����eD@ �.��ݨ��v���޻`�k�W�T(s�qM����k�RX-i�k.��6	 ��>�hώUH7�j�ꗸ~�x߷(���6�����e/s����g�t��j��u�m�R�F0K�Y���`� �Zc���\���,f5?L��&Ix���+�Uy��}�C}���tFJ�>�٭�>���:��8��%n�M13��=B�(!  Pb ��8RE����8��$ H ���:�]�}�;�@E\G���e��PK��bz����xJ��ѧ �cT�C[�G����`;�U !9��q�I�]��d)�t� ?6�mn��&� W3r�`�i�3��3B�w�\��EWM�%��W ��#���^Pb�p����"?��,+= ���S[��cy�s���s!")���Y�p���uZQV�����?�'�A��1�����ѯrUNVY����Y�6"� ׷~h��ʱ�WG�����Z�Z�Zp�	O�����w���;�¾����{4��_�hF�QgƎ�/�����s}- ��/���3�����.�
[U1Q���`�C(��B��Z�����?~���9�v�ЬV=أg�p�k��^�n��s�-�<)C�2�5�agF����~�\��/�p� ����p��Mc{i=��
g�Ii�L�4@p������.6�k@K�@�ډQ���Uj0M ^��g�q�dAci�*�ɐô����˕����սS�Q�/�TBxO� ��6.��~����!���{*��L���V���v�%��mF9&dl�B˱v��D��8k�^R��S�<�]�SE`9�R�ye�; �1@�b� �U n��i,G�C6��vT�).YV���/1Ǣd��ذ�u�K���B��meN�r�>+E�i� R���H��-�b��ԭ�G�ѧ��K�8�ք�5M6Ҋl=l���x�(���C~�N�fI?�b�#�	��z��6�˸\��	O��BԬ~k�O��N�2�0�z�q�4*�홥ҹ�P����<2�Fy�|���S�i���f$n=L��<����e��綶&f���w��wc̡�3�
F�&�[zbi@��[<�-�:��`�,}{����:e⹄R7�})�R�@�1��85�͑ce�gߥ�j���?�b(o_�_p����Ҿk�:�V�������,~� ���*�`P����]>;�CU~P>c�V_��N�3^r~Pw������!�	��ɲx� �kF�_���g�a�υ����L5Py����q')
[b�a���ol��<g���&����'��pA�)̶����o端���O�]���n�� �(x��X�?���WELC���^�0`j �m)�H��8?4Ex�JѠ^�=�_է��259���[O��Hw�@���,��2x8k�GE��9��Ig��q�z�1�׌V>S*��nu&2Ė�Cӈ��I9y���Ě�����\��m�w	��m�����wDn\9�w$�"'����'�X���sR�y�6�gcf!����kE��o�;hX��eu���j>b�BE��xmN�����8��O�"�*�'w\wsz�������=ʬT�nM�H�ɷ��:�	�kNWn^g��������Ɂ�����+İ���C�4�%���ws�����=��Rf��[/�;\Ь����]ǵUh��$���Йt�X·��[��;�����f����VJ61�@�v�Y��N�eYB����)�X��,i�wXwzbԜ[D��U�<4�5�`m�u����Wͤ�_V�a�sg���#��Ղ��BU�s1\�,�{�3���Sr��a��S����y�B
��8fU�D�uT��j�`�EaZ�GNG��q����d:��6�;j�N�}λ;i��ժf�c�2"��<��'M*m�8VU���K��U�S\3�c���*����*N}}J��q�˶z
�aY�wɵT��C���-B�ț�l�S���5��۽��śV����.C�+��Z�\��PҼq:�\Ԓ����;@/�<��+�2��S�D]��M��B@�F�B����4n3��!��	oٱ�Dm���hCH>�,���EBhB��CVNj�M�|>l!T5B���V��tt��u�=4ޡע��>��NuJ��t�`Y��s	�5c�6���s���0�9;��*�A}��h=�eq�ہ�W:p�F�e�SkVb��9&������o��"ڪoG:b�i]^0E�̬��X�VV���.�ay'v��R�D��C�r�L@�f����@:UٖՃ��MⷭS��Z�*̕�'3nƎ��[�{�ɰώbV��-�ef'�Z:�Rʒ�5uok8�β�Ac2L���w�f�b�r6u6�>[��:�Θ�Ӧ�ݝ)�a�E��<�&]�y{Z��a��f�.!��%nVj5��y����,�ce�.������u�paEX^fDF�����t�vfuK|s��t�)�V���,��/6P�sd���օ�Ē�N�a���֚�
��&gwM8'}����8"�u�y�yܪ� v�v�S(vmŎr�8�x0��W�]٬���A7oo^0Q��k8E�P˱����&�8�*u���0��ѥOWvb�Z���d'32�+1gv㾿#7���ګ�}kH{`�w�v����oi�r��9�;��&;��{�;���(p!#A��������O� U�d0�;f!I�dP�Ѡ2\���l���ñ����9d,���N�j^y�	R�!�������RxQ�Y�Z��X�HnځԔ�B�Ce4p���Ç8�7Q�bN��:�2h5�ʐȂ�CV2�r�iL:t�����!:�!��b�H&�NJ`A�ç�N�>��dʏ)2ƪ9�kX-(�؝nbl2�sM�'�0�������'Զ-���mqm#�)7�U �m�م0������꛳|�8�{�6�x�8����6���$�]\��7���ç��A�b�2-���(R��9��k�L���j�+PQ�<C�@�@���A���b�]T�7�shT��|���Ǝ���qM̾C.��XDȔ�u�΋8��n��(�� �[�28xcd��Zm�9�3o3�����o�|��z���{Q�^t3?��,���f5�fyH�ٚ�w�cݢҨ{����1RW�SVX^�p��,�C�ү@�4��P�N��b��Qh�m��̸ؕ|�r�W�P#�}Ma���ma\c$�Mn��jV��^�V�-hռ�tf\��+�z<�"���Y�����7��;����E5�;T�#�ͭܫ��B�0���?��A	r�c	���9��zxr�����ki�$ ^�ͬ�}<[_&�5*��~�6�{�}���O�u���~�u���XV��qi�_���*�P��͕��]:2%veB�����1��J�i�6�����0�ePv�~�Hżf�'z���\Q��mHj�a�lw�S�h�:|��y��]7�H�{N!���Ѽ�օ;A��ݳwX����56i�n(��<��s�$>ư�����Yf�μ�ye+4���"�v��v[��1�-z��г���>>���A';rt |����"y]uu�ܒ��D�u1f�-�C�TŃ�v%��<�w�t�)��X���t��hQ�eNt �� Kˋ��"��u%�d�)�/���ҹ�FE�kØ��[js&����+9K/~x�5������~?�é�~�)����v��W�&&&��\�G��#��q{�!��0_��C��g�ă	$�ѭ��7)^�3O�'p�>��%���\�r�CY��c/����'X��H��B�lz<n|�Uk���:��a@���r���e�XWɃ�G�"�����FFPg<��cF߳���UJ�h��\���.hj�g�����8'�G{��Nܟ4?���}O�ƛ���M���e~�1�P�ڀ�k߇?�����j�̇�J �i��w �V4g.��a3!���H��z5��w�3p�þ9���H��� ܏���.�6T��y饂�M6�2��WBc\n�Y���덩���Fv�*��'��܏&��G_�9�j��g=[���KP�-��;#��6���P%V���.�:�Hm��/K�F}������?=�S��~Bσ�h�ŷ6?�3�i��\@[b򺰓�u��5���lA����x�uC�oO��~�b��~����_!��/�⺮���&��V��kj�S?��f.����t.���仳5�ą���2����s+�_�����ߩ���J�(W�k���^wWD�uW�u6p3s�{�����A��,:��q��W!���Zɣ)�sjsR��cb|:��f�d0� C B1����iw�۫���)h���Wifz����l` D�$l�L0N��u?|]H���۰�T^�O8��,���ӂ�Ґ��6��!d��dҫY�yd<�,,t�6k�����`�g)��6�_����u������������$������Eգ"E���ԧXq��I ^y�ז�,��Ŷ;z|�k���fO9G�(����i��G�Y4*�Oy= Tw=��T	��g�j	ٹ$�g;&�猏9��A �|B����Ǜ�'��O���z1��K�)��oN"�e��5�=0��Bj�cN�W�?���?����-W����BM�8HZ�����j�W=��3�+���/<'�ˡ<�݂��0N~S������(P��%��Xd�E��Ə)�[]F�P��ږ��Y��k�8,��k&ZAxg�5 ��@��~C'�ؿ*��T��Ģ�����.01��'ѱ#2�ߟ!�訽[�a����X��K ���_��j�%��<��8s�)�'N6.݀��n�x�$�*�}F||h��_�ܾ����T+�e�Ë(�\R���X�s�S�N���h��0fJ��(��l�.>��R�1�Nb�(�maxD�vt�̎AR=�v3eFΗ�nU3�Vlt��
�4��.+�,�ٜ���������ɵ����|_��88p'� ����� Y��yli�S�B\&�ydr�z�'zc�R&ߏcȫ6�66t���{�V/�|Oͯ֩-0UD���Q;��Ƅ5?1����_ߪJ5�z�U�~�8��j��Hb�\�|����/�=toT�.�G��S��Qf��7�������X%�@~;xm�g�N����\ի���=�3m��0�%@t����֘H-�At��p�Z^r�Ҏ�A����<���(��E�aET��Ī�~�3��Z�f-�| ş0f~j�����6��EӂV���6i�̆��Z+�C��o����&���<�mx��(��X��������C�f�r�a!��Ky�1�/(��r�^��lҞoM�4"�N�.��q��EE�|�,鳞�d�[����;���2a���n7S-����MB�g��"��Q�ؠ����(M��m�:cw�\�d �'�����6�>���7J���	�m�nS�I ����A�sm�t���IV� S\��u����E�xE`
�{lm׶��g�MT��h1^ؗ�jd���Ƃ����qD)���nv!j�e�������Yީ67"� �覫��+���wѥ��l<�M�N�N�иEd���9Tk����S�������Qr&jk3ڮ�����; � ��3 �(۾D�x�1�u��X�Q�q����ސ�4q4��!��K
�>.�r;ʪ�ﴲ��q�J%��1�p��;5;�y����-&"�C	b�מ��g�u(ܛq�����h����S�R�%��t8̯a����g��/Ţ�GT)�纗�\��,?�_n�re�x�q��`d��.��,��i�am�b�5�W[�ɡ��g-�� hfg���������CR	o�v�U��,Ǐ�'Ҁ�L6Q�@4�:�Qj�
%D����<.}�����T;�2'����yg�|����T.�&�d8��ua����U+��{U��>�֡�X��c`��U�q�`��̛6=Lb]@}L|�����;��+'oVu�e���`g����X���%Յ�)��Sx�Td= �n췚=S׹�D�������nsk]<V9�.5��Qz�V�iBbo�h^P`G.f���\d��YǄ�C�DlD3Z���Lպ��3��D%>���EF�V��2J1�\r1@����f�'k`��d�/���?g��Ѻ�T�ۺ���L��3N�ьbE+ZʡQ�j럯~/��6ee@��Ve��c	��B*cX�Yqcݝd;i�i������c`p�A���ړ,���	�ί�E�<��)q�7yrrг����L���U3_���}�y���t!���ь2�ݞo2�gbr{li�wK��f�.mmA�B�][7f�ʥ뺅�0��hrð�{������ι�q��E�؊p�b�u��r�p�(H��m���:�e�1o=}����S7�x�G0�䰆?~}����|�g.L��ɯ3�%���=T	�a���nO��զ5�+��8�3����f;�c��0�cPa���uoM�J�ze�q���E���M
��N.�d�i��Nd;��l��7�A� ��/�v͵��xo����*����0��W�����@��y�<]�����_=���~Y����5���_��P:��eb�W��M�5�H�U��cm}��s�l��Z�m�dj�g���ǅC���O�9�,�v{�'ى���w3�)�kd�R\cS5����̼M�i{��$}\�;���
�,�ߕEV��D0�)[����D!HY�h/��ЃN��=7��nH��xsC#̓@t̮����	]���]l�%P_��y�|��W���^�b�嚒���<��k{;���v�a6�A��5��\7.���}.�'%�Wd�:�ټ�]�뗼T�_ �p�o2ȍ�oay�@��`C�( Bc�<1����bcu��[�(��n@�������h � $�D� ��d�y��_���C�	7 B��ǵ�P�*#���^��:c�n��Fq��W1e�#���;���cr��c3���M��k�^6Es��1�7k8��-n�� �a�<u�'W�(jQv␇am� J���~<�& *��my�����,?���	Ӏ�.[[���ȅi��Z5�lݦ� ؘ���H=JN� ����������q->{��F6C���pj��9�{2��u�d��k=����S�>��rư^�c9�Ҙ���i8;> ���*��]􋗼_�5Ç�̴���_ �Ԗf9���*S+Ҩ�Z�n&sCH���q��/$|ʁny)�o3y�;v�~`�a��{`���B���0�*�����>���[��]݅�\4�uL���.���������M
��x���)��#��YS�5�6��2tE��,��l���9���XS�nKr�G�a��=�b�������O�b�����f⅘�,?[d��f�NE���	cM�� e�u��$k@|2[!0x�[���X��5�����G*��w��_��t�*��ȣ�_H�Y��I�5�ǧ�eeC�j���c��f�h�:�ӝ��-��L1�2���:NZ�g�4j�f���(�#��u��h<zv�=���v���2$V�Q�����jT�g����P 8���ka2���_Ox3���`��s�O���=yʢ?��H�p2��GD ��=��G̯Y��1��!ǐaAр((���>&:x>����et�T�fGK^E٠��<��(p�(pNU���]g��9�zٳ�6�a��nx���n�)7:z͟ ��uc������D�j�IԤ�W���/�a��B#!�a�%��]����C>ox@o_��C�S~Ĕ'T��*�e|��7��
�X�֟By�#��{mm1Ոi���}6�vg�|���^M\�Ŏ�(b�=T7U˞�	=_]�^�m���t�u���f�.����r	�^VdH�oR͆i�d����<|�V�Ï<h�8�wgc��%K�Ҭ�Y����a��sL�f���q�b�H�@]!a-#@Ӛ�wfV�]�*p7%#
$��Sa�b���7gǸzcԲ�>#�V�S��gp�~�nۺ7��j��}���6r��������nu�R9�ͫ�B�ʴ�VIӱP�͋f������n�;�s����C�����x�[�߀�P�@�;���J9!�����%�'��X�oZ/��y��g05�l�Q$�ߘ���nC0|P�Ȉ[�1�HO�1�~ك��06�Ce�7\���r{�,V�.��m�\֦ܝ`����71�{��:�fq�ri����kFi}��7۽wvL�~ӰKLw�;+����:�4CI+~��ۦ��v}��>cAI�~����{~j 5h	�Ֆ������@C�@���Wuǡts�Ϊ�:��
����<��VCb�(��[�#a�-ޘ��,A���zarT0d���/d���-4�Њ��S[vt�s7��"�?����;@���vU޻���u��B/Y�L�5S(��d3iwp}���̵��:�U��� �?/%��:2��8�ox4�;�rө���M �hp���4��\�!�u$���nTr����ٿU;ׇ����W�S��~	bxggo1'7��f��o�����^��)�W;�L�ȏ#��P��0���EG�=׻v8q�-c�R81��wXWL<�W;�L)ڋg^���黏t���#�%�N��P���S߀���K�  ��Շp?zzn�}�ҏ$�\� �YuN���l���뵥�05Tl�j���ӹ����NXFokYL^�fk�\�ئ�V�hycE[b	ꌽ>�D��&�!���^oM�6+��m��s )R&�lԬ��:�d��}���~�X_�[�y^a@�[�����R�+u��ᨚ\z�;�m���Z7�Gf\�OCy"p�o���R��Y NP��X�[�wE>�� �6,�k�$5��c������ۥ�<��6/��	��#�����3y�4�Pѱ9�ѸM��Vt�O)㻀rȅcNs(ReP�|N�����-.�S��M��)�#��4gj��F����j�G{\n	�r�[�
Y�����������*<���wU�P�;9���q��{�ǫ��~����3�<�pq.h85�\�����7�h�����8m�X��᫛���ǯIKy,�����c3]F�"�S�~Mo/kGJn���J�k���\h�X���R���2Ҙ���z��R[s6�r�Q��w2`���ZU�ʣܹ�]��.z�R�g�l��듈������g31�Ζ����������9n��s^I�4:;7λVc�����'?am���n�7*W��v9�Q+t�&��re�n��8;�	pѭn��uO�n]�[����԰^KM+J^�=���,;��=ڪ-���%�y�Q:�����U��Z���a_P����{3�I��͓�Tb�>X�������p���:'�X���lE�j�9Cg*ۙæ�j�uu�G2��2�nu	��*W����5�,��T&��o9�1:6Ԙ8oY�BR(nAKk�	#�ʴ��|tbk���GA�&s�u��ds>}9n�
;i	|F�2�׸�dXj:��{W�µ�2[7�X��X�m��t�nC�5gHP�7F�:��/NU#����g[��r�'�d�̋;� Eݙj�]K�k*�J��z_ݼ|h�Ƕ�ݽ;�Y��-iW���U��3;���p��4+ճ�j����*���!�YH!jgS/��6�F4�|�w��z6\��"`�^�)�wXy+u��no�<W�;��W�p����%��W���y�Mo�_q�꥕�~cOT�@�@�T*� D��r��2�~����ぅD|����95�2;\<(��Ǎ�OL�?0�h�A�5���H
!x:HBc�~a^��MC����8m_Q��/�`��Mh�T�����h���։uL/���VY�8��Y��u�D�ñ����<�j\�x�lWS���q�AE+&�-�ø%���J�N���Α�^�̚����F{{U�4�*IF[�.<��b��[��{��1w��ޛ0ӥ����Tw�T������O�ow���u'����ֆ����,��fV9N�n;��Ep�-S8��"��W���fv�{Ul��j�)ĩ�4k{ƨ�E\�����qu*��T��af��6��%��Xq9�fv�in>a���Y�r�Ll@���H]��۝���6,�,���6�ZV�*巯(�H��D�NQ��3�q&���N�sIW[�]�\)9�.����J�<÷����w$n1x2}��3�'�0A�vINc[�Y�SS�L�2W	T��z��,N�fu�`�זk��JFLֲ����;J�SyxS����M�xl�]�5��w-K,T5�����\Z�fu�s�YJVC�v��[|�%�k�U�s
��񘂢1��po!�����_�wb�8�C�#8Iݛ�6���N�d�Ҹrs�w3c�� C(V6b��<Sl�b�14�M�x��u�����b��cOi��M�i6i[S��ٵi�ZM4Ѧ�ٳ�Sz�kU�G�)A����PA���$M�F(�M�Ab�)�E^enj599FkI�c�@1��M�H�P�\� �f����t�}�l��Ֆ�Tj��=��X�V����<=8p��%��M�LGmd}�Ho2Km�ؖ�SN�=:t��A"R�/s��G-�>_,e�݂�����ӇN@�j�
S��Zz��u!�S�eKb�R�6t�ӧM�u�"uY��9 q�N��L���t���ӧ�G,�H��;Z��r��=���S�G�N�>�Q���~��f�{{[��C�fP�&[G`�U4S�:z|t�r�(r��S��Ŷ�1cI3[$)C�"����J��!"B�0��[�f�֭e�]f�l�A�Ka����׺�c6�]W][c����,�n����[�Vu���[�)њ�U�T|A����܍�Ǫ�Uh��1Za�h�h C0�#�P�i?�I���	a(�����@?��e����=슘X@�"E'��	������0�Ǟ#/�������y h2Uv�I��z��i��/w-@1�
�a�6��/����Y�6�&�1��.�.������ZE��p�#D4�4�������k6��OQ�{{ {ۙ(�7���z�́�[�#q� o�M���M��l9ʉ+�xe�b=Ӳ�g�|�|��^�L�|�v�Qrګ�Q�$7(��J��p}�h����R�5!W���&=PQom�RT-^M3O6e�u��zNk�9��}xǥ� �/X?���� �Eb|~��|�iO��N���r��Y4��՛ÏU7�sy����pSx�]2���;"A����������A`� �ː?���:����s�������Pj�GpR��)p�py�Έ6��*f�E!ӯ�ћ��n� /aٙ	8��b%;�˷k��oqU���3�;Wp^�Wp���/��|qU����9mQ�;���#�n��Z�T���sf��L����W�p# qĹ���)�鲪�#rj�ql=|�`�Gr�1����4�̗�fv�WZ)>8%WN��v]����~���,��©e-*�@�f'9#�K����5] L�T
:v.;��5=ԧX�ʜ��e4��l�{�-:�� 8�,��3�w(Г�/�ϵq�+xQ���>d�5w]���mN���=�,�
��%�ܧ�˛2�aA=Ub�� ����]�j�}��qi�b2 m������3��g�ƺ�#��3�2��S�<�_�H8�13-�
�Tf��ژW|](�N@�B��a��np�I,�Ek����2��+{%C���Mv�,XQnP�M�|-O��/�>��0
�� #Z� s��ZK;d皲pl������p��mO�;�
V��GG�����x��4�=����W8�ѧ��!�9<`Q!��� ��p��Foڶ31z�"w��{[��;��X� \���SG�w`X}^A�k��>��<눗�����|�D���Hs{�)�&p� �a\�/�%�;��ְ\����o5����gz�h�f�eU�Q� G��!E	�7f;"�R\�R����V9M[���,uk6��i�M�>.��L�u!�6���ӾU��s5?��Rҩ٘��0`�o_'Ύ)��}�س���e{Vǃpa���4���&2�kz��>Ue뾎��%���x��Ad����U�U���Y��mE�`��-�2p������BO)���J��@'�{Cr��@�R��s��Za��1ا3s)�-�vd!�"%u�V�@4���q�"�V++�@)_I(f�R=�YT2g�8��@vq�R�<��̙z�}~��`��%vM�/>��/���D�^{O[�]Or�$s����l�/���{=1�+�"Vj�B�s�Vl���h^�u.+�XP��.t���l 댈�'�&u��}���nvf��c�WeMg\����������@(Y0�}y��?UYWCtP�����@&�������#�������em�M�?gva:��؞φ!a��0�S\��{I~�yƽƧ���r~WnyFn�;3f'��%��GsvkS���l&:`��w���i� ��.}O
vGJˎ� a����ɠ�ĄX �UiU��S�� �c8M�=rUl�t�&�S�Yל��݃!��B����~�n��8��N��?-���[e*�R�--:���.��C6_������nW��m�Hm1��-r��7n�b�gxWtm�@��2*�n^2�� <W*�Y�M�x��]�Tk�ݱ��Y�(Čf��X̱�X曺���5sr�����E��b{��T�5�����β�b��'7��=+i�\q� �o`i��Z�z@�5S�C��0ֳnfn�����(	]]r�؞�kM��\nj�y�+Q8=x�ߔ��5a�7�րn�NuÆl4�ϕ6�J��^8U�y2U�8y�/+Q����n6ad��HQ�=|Ee���'+��@�3���O��Ü��j�}�qU�{�7[���"F��ϳ��⽢pH	,����sl�\��Mo\�w鬉���]Y����<��v���D�m�`.����Ek��n)���ʝ*U�Ԋ���6�90$X���ú���;�t���c���U�\J��ctZM㹙�z��W���٣���A�]�a��?$ի� ��:���B5چ.�����E�Z�"҇�T��8D/�p�.�kU��r.��`g�`G5I.D�ι���}%��=�SYn���stWr"�V1�0���m[c��۽M[�]�[��t��iT�3y�ZY���g���I��h`�3�pX?� �����3R��;��:Xќ,W���X#��7Y��ћ�1�^��������^r��[Ǡi��{Zwj!�e�y7��3�,`C@S�t��Ͻr�>�^����<gC����$�ig�I�}l׭D�x��,SG����\L����	�O���_n��mt����F�k�u>�i�Hd]����Z(WE* �J���ƫ�%^vl��� 52��@H�9�\�|����&�D�,���o+kڭ�vWY��������P���J�a͍-��h5�g"D��90��1ỻ��$Y~̸�hZ��:}�f��be�w/�q��AM-�%�S���g$s�$P�4CE����w!�����5߃�ZG �9�׺�v����Vl>=^�������d6 �PJ����T���h��r�;���/ڮU��fO]��1�d�����+�_ n�u�+����	G���uvw���]N<_�����j��k�$? @�B�{֏p}wܺ����U�x���呰OZiT��N*��[�ޣ�CnJ}
�,J�k�]�6wk߷����)S�3�d/�&M9��}�,Su�g�
^5X~��龌}�3Y��/@��O�˅�����gW�Wq���^q�����6C�]:�v�%��cg�^$����q���vς���j/�i�����,�:mƌp/-b��6�����Nl���{�F�\������B~�Ne�o7T3�/p�҃zo#"���G��8�����}��Yh��r��Ɨ�>u~����r���э\XMr\smU
�D�Y��KMS5��vlc�4�D ҉~  .���ߧ�d@h��mhȈ�1
 ����*�d�:���Zi�1��nI�n ����*�7n3qh�b2 e��P6��e���"����}�Or�ƽ�����k�Z �N0$�}.C��w�ܮ��n��xs�=��;��V�����+�����{MXhH#y������[��J�t�R��ӱ���F<�9�l4굌\���o3�\����ȯiH�t�
[�h�a��fd��U$���<���5�կ)_k~D�Cx��k&�5�z�|�,��o�!�h�I���Q ��?������D�m�rbɺj.����b�������`�A�}�7=J�g�\iϜ�l�Ү�k-���T�JDM���ׯ��=�z��/65�A�$�Wci�����6��=����}eDSUܨ ���h����1�E8��%s�r�ʪ��)g� �ߑw�Q�	����UղY����暳�i���sEοv�,!�W�����jz�k�,�>S�iR�)t���V@8ڳb�[bL�K&�A.��X�@^2�l�z-^��ӛY�:̑zM�8���:g0�&2�f̩g��霉�;;w�i����G?���Z�]�{y�b��_��y�+p,͗���c�g�N�@�[>jP%�F0�����h��1�!��]����X���*�sQ�*��Ŝ>���?-�����~y��y�ɔ���Q�&��w-Ě���&n��m�x�K5���������l��<��x��tu�7�h�ŀ]uS�
�'R��a;&v�����X�l�<����sy���UKK�D�Z��|z�U���]Ik��J�Fb�́� y >�
�&WE$3�,�H����pkV�y��>H�D�!�î2"1vma��W�
�%I���E��n�>�ۚ�3��O�x�o����y���ATvՉ��0�����g;�(��TlV�t�y��O���Л���/���ϗ����;�o{綸X���ƥ0���d�o�&���lWޞ@�1����wT�v\�\ޗ�Aƻ[8s]@G"�n閭�ciu5�]t̘�l��3��A�Tuxt6�x�e�ЋrVa۶,��|���6�'/L���>Ͳ����$��u<1@x�G ���T�P�N��}�'W&��՘4�^ދ����3����-fCӱSn���u�7�8�A#:��_!R����`~��x�*��;�56�6�ڵ�tT�M�}��,
a�C>L�o7X��8�9i�Y^*�җ�!���ٷ~�{�~��
;��V3s�������k�Z����{I�Gv�C9�Y�}��ڭz��x�	=��;b� �{�� �V�GlS��k���Ѯ�l�r3aƥ�^��]]��y��	�a.Ԡ���R�Sz�,B��΄и(D@`�@�a
@F ,ʍ#M�DC� ՠ=�����ڝ��{s��,CXD��")T���V{�.긽����lz�썂r�����G%���e���ޞ�T����6�͚U÷���:�BY\]��[n���̺@�^����`���7�L����2=+!�f�P����[�����^�˟����u�P'77<ړ���F�[Lq��5�'\���0v+�����8p��l�� N �O*���%F������	��@DߢMde<��D၍oOu6:��@Dr�:�Ea��Z��Iq�����u�X*=�������L��%C�E:`�K ��P�ىVٞ�h<7zr��z�
"Nnq�θ�`�D�e�89�]Wm�&���7m��G�:*�ޘ��m�C������j
���#�3q��@@16G�Ǿ��.��#9�XW.�ok���M� ����R�@�lS���L�Gw){)��S����ꗻ��<f��5T��ʂ����Ά.���ص3�Eb��C|����^9��P��5�n�7��q�D�y���:� ����)ǀ�+"h+0a�re�`�dD���z��?�� "����Z�@��ϰ*��W\7[�����Kih36���lSjW��}���һ� �&|,� hn���ؙgx{���e����yXx[�{Ø�[�/S�U��;	T�\O8v�	���͑]�����F��;�~�l���~@�g���5!]�X��\{C-JLb�����/Xy���f����ٻ1�E7�o��3��ɹD=_n��Sb��[z�5�a��y�����Ҿ��UVƤ5�r�D`m�������G_�� @����k]�葦V�`�B�͠ ���@�S�qZ�/���J�㌭-@���KFr[{}�)V-�F����x��=Z��f�썾���m��sٵ����,K�K5��8�ÏqVw%]�E0���K�𧜦��[Ʉ�0���,��Fh\x^��=�����w�;�b����j���35�U���s��f�c�bw=i���!�Ivc�4h�݄�r�,�,�.�K��ms�	u���#XM��V��3jtuF�Y���"��f���� �b��4ػ�J�������a.v+lS�=����ٛ�����s�w�-V�f,�wR�`�[��N�8�f��0����[�t���%X���c׺8�"_ڵ��a9������k��,�Wx^�l�Y�ˇ���*�'�yLX��lf�K�'Y�<���`���VuC�k�e���b��f�}:�+�kG������>ᮦyW�q��g`G�-�(��K���>{�GwW��eel�"g��(̷��ܘܝ�)n+�E�s޲�<��QC'��#��2e��A�0���Z������*l:�cv:��"�-�c3A����)��J�c���N�zV����Sz����!�b�x.�M�J�jr���˹kr򶱬t��P�]CB��B1JG6d����A�xf��2��,e��Zٝ݁N���<��lPC�G���%�����	VD2���Ӑ��󗁑�I�у^\�̖���9����S2��l{w�;��]�Fz�j}�tV��Ŏ�|pW �A��S��T�hv,uQC�2��HȆ�%���h��UC~�4P�cE@��(87��4�����F��pB
w�L���u��չ~��[��֯5��cs�j��FE�9u�0�kk��֭�ꔷϸ�j,=�[��=�A^뽒�e�����Y7ǳ�L��QZܶ����7�1��,R��bC��Z7L�ޝT�ҷ}H�/J�e�R$��kv�zy��Pܗu3:6��,�Uc�����
�8��+��Ϊ-'�s�:Mbb�1]�*Ⱥ�T�4�gpapr�u.��]�T3p�������b����q�,�dǝybT}h̻E��>E��\���:��2Dj��W�m��7��>�ơ���O[�74�P�_f��B�Y�Ǧ�C9�d��hWr���mu�Z]J���mvF.N�bl=��#��8SQ�ԼC3�6��[�j��ͮw�a�)�HJ|{j���d��03���!P���m�D�$%�ˤ��w�X�N����ڕ�c���,^��Z뎋�k;e+b7P�$��*�q��=1�J�
D-��4wH�K9�U�=:�č�B���o>���1Y{�����D8�Q��%���|����eh"�;H�+*J�[ݡ���ü	��ϛWc���W\�^	�<3e�톧W@�!Y�c�b�Y�>�3M�g�FE��,���~�1��$�\�w+�I�ݧ9Ν�(pcA��i����s�Z��!������Ha4�r����JB8ώ��>���%�MT�3;r�Pw.J&�˹��� �F͝=:t�[+/l�m��� JT�
����<��:�
F���D���!)����Ja�'�m�� �p���~?��ybs3*Ke�k"v�e�Jh����O��K[�3OP�B1/vE-@Œ�y�C��ښ�H`��9Ð�;@�z,%�
h�rV��jV����e-E���Fώ8}��-n��["�a����0ه�8y�O���*��\�$�5&�:��	��R�N�C�\N�(iJ59's�Ps���m?<�V�zt�u.��9ˁWL�wUnwE���9{qEKr������.�IY\���@���	 2 ��爉�����N��n{y�2�>"`	�~Rޟ�*0��8�KSN[&��y�xf�Z@�z";�7�q>�m��Xb.6��^�u�Z���KLixn�g@��>��`n�á�<��.��c��ʺ�u���3Ѥ@�V,圆ʱ�c6 �<^ǀ.Յ���J#���y�Խ�]��,g�2H%�$֚�ߊ�0NGM���Xa|rC�nQa5f&{��Qesj�{Vz�l?�0�q�5��^�*DM���hm|^����ֲ�*��u�{��p�oi��_�X�l2�@d�@^
�5"3�}J�!5e/�jp��1ռ�g �`Y#:�ɨ�%��{����=�HP<8Ɗ��"�cH#��^iqvzz�F �eV+w�S7�����KM�jS+�����Z�1y;>�](�#%Qɹ	U�
���z���a�	}�^d�����?Mv�|��ױys�f����x�����B�>R��TyL2�Rh�F��'���k�`�.ҡÅE?A4h��(�ұ�6+��[�J������+�S1nJSg�;�\w+CM�pަ�UM��c�=b����f�>��0�?�«:}�Q�Qw�����)��+�]% �>_|��m��j�x���k�J\�.F)��ƀ�""p���_�m��j����n��i9�:�s{�sL�7Ͳ�|�7�:������P� �T��'�0%wM�lR]��D]Hc�.2�)��J�6�|G@vښ�f��F?��S��-�}U�39}�=	�KE��x�]�"�)�ҭC�[Et53������i"�X�Β7�b�u���P�YW�h��Ŧ;���ǎ}�B�Di�A�[{�}�I�9>����'3���V�������Ce�T��{����@V�8u]4���1��Fѽ���fE�-h����m��t�a�l���}1�M�1FD[�m�Tlċ����{���8V�ҧ�����xh}v��&oH��ʽ}&���OƮ�4�z"����FM�tM]+�X��싖%�3�P�6�h��G/���Q�$��X��SnE�_��?^��M���A�zxbų�q�~yU������yF�5n�cӼ�����m�WS�C���ܾr	K���G\y�W_lF��uR��@`@��1R�jܷW3������⺧���i#���p�g�v\gn��W<�F�9��<dy��{��4�����Y����Wq����Qw���9���@�t�9c�浀ޛ�l棓�%�S�7���Mp����٘� ���ƽ�����+ή��i�o��2+��3"�����X�<�WjzJ;�c���x����5�py٦����z.wDf��Q޾7��9@�^캖��W.��F�9bD�	�*�ʼCNt�j$�[�!'�k
��{����]�1��m�,���;����f�)����1���ԕr�"l���2+>;_����j���k?w7�|4	��a���E񛌀(��Ӳ����� -YU#��Ɣ����̭�EN[a��`_,w9ѷ�Fg�-7�P��<wo�_Hp���r1S'��0YU��]�Zn�}��#��ܻ��*m�6-敫�P��(q��I��������޲.9M,�T��f\wL[O��s�֓{X�ZOf/i���˾\^�YJu�<��wr��˶J�wG��R�^I��%�#kE��%� ;��V�;rSmG�@��(1$纴Tz���#WG��;�;�[w�C�%��}��uw�5�m-lP*�����;>Ôl:�O2�:�'jw�-��5 �R ���`� �,.@db�3n� ��˶[o�7��ъw�ρ^��7(�	�����F�~�ɓ^���Ub���դ�_Z^�ΟE����I0�� ��w3��5@��yW�Ø�z���E5n�4��u�xP0������
�z���	(�����������$:�e1碤GL�ԥ��cx�u$��H`�Z�}�w=$vڜ�wY���#]�
ϻ��� ����ys����f�@�+��~o7XW�6��ذ����X|T�Im�����q�y5un����1��ȪY@U�W���ߣ2�p�c^��s-LTϢM8��Ice�p���;������o�gkc48E�Qƫ*�=�!��]�5��.$���]w:j���`�wg�Q�H<��šjἻ���`����V��\����v�U�R�X�ă�6��ۂ��;`�����`>`-�FQ?�ﵡ������~��6}��}�~ݰJ��Wy �ޫ~�!�<D����l��}D�oVz,�p��]�F$�N�y��VWm�H�J���"���?^ :�e�@axr��J6+Q���ኇI����cH��wNuW�Z����`s�2�eL��}v7�׏�W�!�LNi�ٙٿ4X��=.�}�ue��64����`p˓���	�a�	4���YYx����%՝�kӀ"%�r'�VM�����@|d@�"P�4�'���y�Vwrۮ^Y�*%�;�LrW�X�8�-w���ȕW�uY�6Z;z�gF����ZS?f�"O��}��Ͷz�󊌉��f�����	}gu�c
��t,��x�^����k.�4��̈́J���mb���*āg,g8�j�%���HFW�~��N!�~�ح�:���Σ����}��SԴW�)}1ڷN��۽�U�m�\�^p� �H�PA�eG�f4޻=��D-��uW����:p��ZD�s�g[�:��U^E���xzX?��\]șB55^K7�M?ӥ���3�e4����'�>���U��rn���u��/8 L8�tc����RO톼j�=�@�S�tN����"%�G4@`���ׂ���zv��gh���n��W}S�ዽ\�K�VL+Ҁ�M��:��O��(��g&�c��9uvv2n��h�>�f��Ht��<+��dl$� '�*����n��K�~%��Ѱ7^����t0�Eǧ6ht��iF�u�E�Un�Nټ�H�����{���緅��b��i[�'�t�F�yLNY��f�z��w��EU��p.���[͑9=�Z��'��$6��"�x��Ԉ	�ۍ� ��g�j�h�K#��ț���Y�k~YՋy/�W�}�+Ft�
;Z`W{���
X,��o>nh�����~�je�=�ۂ�{��a�fZ�ǩ�)��
=U�jW��_�C�T�V�_],�z1��@j��l0���o��(3G��z��RԦ�>�o&�x�q5���U7�F���
bv3�9-k�uVP�Z�ڮR����ţU���h!�F(`�A�b�/�e���>q0�HP��o��ȸ�Dj�\0`�g��f8��Y"���F�FV?O���vkgmT�B4�E͑~�U!���
�ׇi��n<4oP�f�L))���=�y꿓s8c���[��D���vU�#J�b�)7 �z��L���^�������, �����4u�}�Y�Cㆾx����8��0r�:�ݬy�G6��!����{Ml�c���^@�X{95@m�tu��'2�r��R�܌-��cz.A�s#��t5��1����9i���&���~��-@�*&��'G�*�1R���[F���l��`L�Zn���V6 ���d)��e�^����u�)��L��%.�0L�"�U|��JvՄ���»u��p�΋<Ff�	�tJ��p�}<7�����+@�-H*�d���i}�5�4}�l���uِ<�~:�Mv������Ȏ��V���
y�D�쨍\Z_f���\x�Eo3-��p6#?\ �O�>�QZ�j���f��W	��v�Ւn�E���̶�����2f�n���E�.a�U;��&s:�����y� =�	Z�YN�,}�=�5r�2�o�D��옵 W�!a2��Ӿ3+ڼm�/�Eq�s{^�����.r]m��#§d6���Kmdd7a��v���l�u'{��)����/,�12Sbǆ��7Ʋ�#���z��F��m������ݳ�B�mRɌ��h+B}���� U^�]���Q���WU���1���jG�M��;�z�{�M��� y�0Vl
�(���������G��`�n����#�f濲�K=%�������� �Vݮ���&�]�3:�
}�`v�s�����5�^�/һ/�9]�x�f���nđ��>�*DZR.�fqU���޲ln��·!�Z����h{�����oI��>h�Rx�𫽢�E�g#t�[u��έ��euX��-�>�R���]�Ql}��٘&y��nwG��䪻I���3��g�`��c|��7x��f���|����	[yb�̚��V�S��]j��r�ֺbv��b:���_VfZ�߀�`=�8 ջ�I[.�v�mS@�o"���	w�ϣ��~�w���Ev�7d����Aʷ2��?��T��)0%�K<H�k����m�wvwvn�6M]]�]��y/�S��|l���Xކ�)��W���=YǴ�"�o ov/ �l���,��&�%Wʞ���y��.�T��4S���޺��g��5��x��pIa�0���i�]��UVx�˦�uS&;2/v��{��k��Fۖ��n�J4�ι�ׁDҳaE�ٙ<����΀��x>��d�����W"��\�--w2�̚�]��4�ڮsHU�t3���g����s�wbr�0�}C�^!��tM7*�3���@ ;�a��d�h�1ǳ��E�yi��]:�e�o��Ξ\qt8�$􁛜����MX����`8۸T�t�����un��:����ZEҾޫ��U̫��C�_���l�2�j�kxR����x7�+�� �@ˣβC�_M���6����c'�Sf�7�ղ�����aO�X�3i#[4���������@o`>o; �K�$�7(9�	�W��>N[�3�	a�[�����c�:dX�z��_-S>��<*N�c��|6��ø��o�HVF�۸S,�f5,9�r:%���F3U�@ �|�/��M�EC4Y��sw�w�$hxF�ٕ�{�Y���K�x����&����SS3<˺�|�Z��X2y�9S4�s#F�N��#g�Db5	���M���+�N7�>jW``<k���Y�w� S�5P���
�E�XJ�6�;��Q�en��GN��p��V�zޱKhm��q���Ks�щ��;S�^�c��a9��]�P9W)q�A�@E�!�3�6_H����USW,3a�e����y%���4[#��*�{8N��Oa���k�P*l��e��]�5��� �=��	��5�'8����0D�L+�Skde_+[��eE);��Wd j���w�c/����5S��5�ꓔ�Y<7��tJ�I`C&]fQK���l؏���W(�M�� �ҺgI��.]M�{�8�`[��^8���*c�g'��R�WLڦ)>T�j�s33���Ƣ�J��utUĞ2�f�����������.j6��wA1:�R�c)�a]�Tq�E��Uhrk��u�IZ�zu�<���>Y�^�̩j�21�BѾթN)��5T����r��T���ޤ��#�������U���
�;�j���ۡm��:��Zb|�W�Hq\\�H[�*�7q�W�j�5��S6��+�n��YΈ�z���(�y:fJ��Ƕ$�t��a[�Q��Y�M<Tľ{q>ק^��ӚV֙���泜|6����v�����喽�ԃ�_�Y���T�b�(��fe�>��i(��6�0�J��p�hf��֍($��&����YqT���77(dy+��W�v�Zk/z��R��	\7nռy�e�����L�U�	IS�uք�N��,b�����qب֌����0ar�6s-�k[Λ&��W�R����W2�;z
�U�G�������K�;3fZ��ъH;�X�hTϬ)l���VYN�:=hj=B�T�q1g��4m�k�|�����$\� u������}c�+�,\�\@��ꅚ���]�;�o����pg�3�LP�:	BrT�����+b
"
f�:�~*���.
�� ��G<�6���S�s��W��r��rh�8�%�[r��W6�% �xH����`�!7�/~fD��Uw6��_�ޙ,��=[ө�����T�H��F�\�c�W±�k�j�[Tj�=IX����3;z�*,L�i�T�#�h��9o��4�+5�u��xl�V"V�n�l�Y��5'[��J|[�E*B�U_+�z�k�A�kq:)@����{���(]�ᘇAk��
f�v�^7�B�[�˿��R��+9�����1|N�G�����	^S�+���zv���ҷUՌ��L���:�E��A�=[ƬX����p�`���s�-�GSޥp%�^os/7���톍I�i�l�e�z�e<I�e!El��t�\�%�t9ٻ�j��T
��@�"+������JLI��]������k��l[-qY�Z�f�g1���W�
��90�ɖ�L�h�Yέ�$۝09Cp�ͩ9u9����ShZ7�5���ۚ9�NP��ι�i�u�'w�ma�4�eƮťs\t���W�*^�����y�mm�W�.�����s��s�t���Jڶ�ei��m�1��1�i�i�1[*���iZm��ұU���Llĭ��Lh��cm1[i��+Jm�1)��( H@i�R�}mQ@�`�-� P��&B��D`�\!��!�$!
E��N������AK�9��JQ@s&Rէ�-��l����?�ǩZN�%����X��C#$���+��=?�ǥ�����
i
Bd
��me8h�g8{>�m�S2�^�˸2�l!�V��õ嚲�j��0��ӧN�
��SC@PӒ�AAT1�C�eUP�G0v:l��ӧ��E����V,��MP��0�F����:a�Ξ:t��ʶZ��=��B��$(j"���a�<:t��便�kY�[#HD`D4CF�L��lOΚ4l�Ӈ����~�	�j������iH�� Nl��L�l�����Jn�)�y�3��l*&',��3��ɲ�	$�3'Ĵ����ʞL�ྐྵ/�@�K�V�E�I,�5'>F\}�ż�V�.�C+��NU��T���*)}U��fɭ���B�-1�1_0�6QM��՚��4m�T)��m�LG�� t6��m`5+y��@a �`�)��f|�
��l��Q�sσ��C_���0�ϑ	^�Y��=/�9���>�;G:*�c,�Xu�>X���@Mpr���m�{p_�h@r�Q��=�5�O��aE	�.F��ah���[����zn���;g(ɽ��\��3�@���V�6�%D4��h���O��j�	�����n��{)G�T�7:��86��N����lu�QS����R�3�
�{7��a�
�E�-�pڮ�G3>l�̔A�����>
o8`��=�왓�Y�K�ţA>Q�(𶘼5�x�����|�`��3�<� k�-�!��_<)ѬY�I�.�cU��9flO�7\0p�3�}�G���U��Çs]�{��Q��I�E�d��?N�{�m�[�j��������V���CY|��Ng�j����V~ݣ�pn,?�b���<R�i��f�W~�1K�L�'���˝^�y�R����eӑ(R#ln��*�xA�'�T��]�ޘE�eO�G-N����;��j���jǎ̼��'opB��Ni�2������d�  �4����;o5��D���� �N���C0`���d�4YaQ�Y�ߐ7��tw�5PJ��d.QW�S��ׁ웹��p�@l¯E�V���	��eK����KlTyю�L@fx�/��7�Ļ�Kwmߪ�Sw�Ԏ�`gP���I���ʐל���/�m��q5����=p�4H���eb�3�P��۝��l�D��Ŋ�n*�]p���G%���gPYkX�%�p����%0��]�a4�U����v�ɋ��N�8Q3Y
 �^��6R�;��ׅ���xm��ۇ�K���V�^���`4�	a��pfqoU�Q]1��-
Yv��u���\���2P������_�S�s
��8fu��aɫ�w?Y:�U�@�N��>�o�ţ&�Bq}Taݓhp�`�sf]���$vS��V
�:�7��P�T"�:$c`ꝯ���:��s���ς��y�k��T�աr�H^ަ���7f
I`�cs)V�e��ʩT�1v�S�F�Oo���w���q�s�:�Xf@{��"�7;�(��R���1{&��n8(�Qp��y�XG�3q�2S����ڝ�����(W1]�+�̵�H7��wF��p$�Y~Cf��=�т�mtAj�{q���țo5ՁA�^u�O���x�{��g�c���5o7^C�
c- CG��15�^�`Qg��u�gm��9�2�.ݯg�b p�@��Il�U����6 �ݸ@1EH�3\�[c���U(3��i�c��z�����[��}-���f5R�1��d�xU�T�W	܌}��ph1� R��1&�8�IUx�î�"�U��j����jcv�\�~�K�\O�6F��{7^\��v���r����χD˴�/SN�`܉�:�۸nT�f^���$u��[���Ia���
�5	���Yal�ny�.��`!�Y %]�X��iޟ8�a�I��B�l1�l��k��n���NH��rWwq���[���;��ulRQ%ޢ	d�v1*������,R��=���/�q���}|b3]U�:]�Gjs���Z�v��-A[-ZǷi��K�
�}엍}���� �`"7l%��4�T��H
5�꜑���f0��\��%t\��>dM��`_��`��Fni/�k��T�y�>�΄���;dȍM�p4L�����i�O��y���x�C�s�ue� Bƭ��� ��_Ov���I߯ ��s�������}+9Vnr�Q@�/�p���Ʈlw�ٰ��&r��kJ�D?oc�Tµ-m�2\5r`�f�X�Pޑ���h�ַdĦ��l�@sp	^X�����ߍhpΰ�劥A��6��ѫ�u�:��_O�d73�_:+4j;�M C� �<F�~�9D�*��aϝ�"f���j�S,�g��]�P,~���sՎ���%i��l|��i>:�.$;q�Y�>KtǞ�r}�v^�w��N��ժ`	��"4j�hoFI�L�@.6���4��P���pW{���j���$vˡU�U�>⵵�L²M�jN���K����Rҫ޼�c#W���lM��C(�H�$�xh�D;���+"P۸���wc��(s*���<G�J�]��U*Qõ#at�|���*�A��Ю���6����i�զ�cM4Un�Y�f���L���{� ����{kfS��u^? A�D���A)����uk�ސ	^Z�:�b�R*f;�\�-�nen��.��6M��jS�O�PaL���d�O���8�����ɰM�`Y M���[�V"�+l���6%+�Pޑ��bv@�"�L	����%�;	&�,��\�q���/8~�e9��X���gw�s@��A�157�!��'צ �	�V���T>V�WOY�͞y8��#��ϝ�k3�o6`3��dQ����[>gn����y�j��H��s�*����&��g�ȇT�*7�U�����YIEi�pk������¶|st�����0�}��:9��I�x;V֠0&��e�˲v���+�{�^�<r��8�ϟ�����T3��M�e>*\	��-���MF�7)��̀9^�Sya,�:)��u[�2��� vʑ��)����_X�m@sC�.s�&j�`�{�mWSN�H�,w"��ܕ��m��^tM�/�!DKͮH��W�c�"��6�B�g������"��̐ƴb�DCtxC�WG�]60u�2l#���(K�gfsJ�
C��8�ox{����:�f�3�ٽ��),<H�c0��N��J����Z/�>��Nd��`gQ��2ds˝vÏ���5�[5M*�73��������U�(9�4;�]}߬%������{-�537�l��ac<W�y�x���s��G� A<�z\�޴�`˜������jz^�h�\j�����q������]V��0�~C��6�y��Fm���3�訯7�+���Pb���'��b�h Ig�o�ٓ�ۊ��^U���w��ڸ�.�➛�[;5ú��I
KF�3 ,��Ed�R�+�o6dׇnԵ�;2���0�h���{��@Y��G.�Wf�iA��WsQl��͊�;K�� U�� ܄�Å� }�c�7X�ڸ��XӌF]]4�A�#��0`3P�Z��Z#�HQuժwk6Ĵ¼eC�ay���d�_/yo���f_%�����}���~���iD��5-.)��b�7YnqY��-:�b�8����h�7X�`�q��jR����,�wV�:c�������]��KY[�φH\'�Z�{.%=���X?��݆jهCtP㟢���N���j�ok���p�����*�.�L�͍�'f@���Nl�p}C���U��4�X`@f~�t0�-��/���<���{X{H��� �[j�m��ޮﲀ�<`0�ŝ��E=��qDq��g������G!"�-���`KU�`]��aQ�`f�x��`?H�f02LvCwDJ�3y��>�OF��	���= eXH� ;<@��)�t��I��:��$�o��f��C���w<�ژ�V.���E���5˼�q��o���rpȬxN�x�{~��A�U���U�W�E�Qe���au��f���p���u;-Ca�̈�
(�eὲ�ɘ��G��U�ڎh����#z�����;�n�K�Ŧ��	��ﲹL�^��8�J:J�\d]g1��7�;��gt}{()�c���C|F߲�����b�������5b6����T�B�t�s�w&�)�5���28�e�c��YW,q�Q��b�0+b�EX75�h�(b�CF����� ��?0���vq*�oՎ�&j�4����wr&
�ݗ���
��S+�L���y�v�Tn�V�>�iM���dj�p	��s��ܮ�fq�SP�V�/=%���<�cG|�������YZ&{���c��x�����ϓ�VxXp��`)3&/	M��1#*%�/H�D���)7��6�N�k7pgh1�͢p�������n=i�-�j��wƓ����ʳ���S�]�n��ob�D�M��*�x� ��b��>�(�[��t6f�n�W��g[�{S�toH�T�ݵ~I���; m�Zހ4K,WX��b�s~���n{�uF ��gP�1�§\� Z7�@��5 w�YL�M�3E�p��w��5k�-z�G_F�� �I��]���������w��]����e:�\&�Q�=c��p��Ȼ����o(7���Іs�3;ș'��
p��
�g0�[R�xѫ�a!ˏ*�ˢ��8�Z�)�F%R����د�l8~iM ���R��w���IȮ��q�t��i*Õm�G%GLќ�^\�xi�ˤ���G;���F��`A��A@�� �( �|Rq8�UR$��@��@�nvUA���"�g�p�� O����8�<�j����f8p��(���z�	5���r磙ٽs�$ �߫��:��<�.ޡ9^i� �z(V<S����6��qi���e����-�d����O��<d2�P�d�`��ڽ�;�7v�)�L=`@����A��Ͷ�}�w�-F3��6y��++��wE��1+ܼ�y�1�DX"�	��{�\�����΃��!�y�]̎����ʒ���v� n���[�o?U=�VD�ʻ�Z��q?�vզ}0?]
�%'�h�}�R.�.��]�.2j��F���˟�6�罜`�l^�n�Q9*�B�̊0�iYP�.'�8������gU>��aA��%���٫������]�v�`+��g� ��f����,����Ѹ±��n��گ��Xײ�<��Ĭ�x+<����2P�ar~4���B������-*d���,뙍�I�k���M�L��/���X�T*.;Ok;$.8�� Q ��F��z�]�v��xrp�eoL�)t�-Y���Dd^�n���i%�z$��S�ީ#b���`��-�.�T>6�� -�\m�,���VǸ�r��]MC�f�j��Ӟ��v��a)b����J�\Vw���/T�|9}WGui���i>�����]7>
C{J����O��2�\��M����2��Gf����쑘݇
�ޚ)6ske�`���5�o�7`��wY�j�h4h�c 3� ��]r��n�̽u�#�6�b���j ��6���p,tC��z,���z�xlt3=��!����������~�R�T����
��y��	.��,���ޟvS�kr��g!��29�Z7U"�"%8p�q�]"�躔�=;W�=��zf7>k^;�4�a���%��Ѧ&��	U�:e-�[4y��l|�O1�g����J3���j�3���w\�a
��[-�S�j���0�媷Mh�M���$�Uu�cZ�#I�B�Ǆ�i�:���:͸f�U��8�h0��Iat��e�]n��+�pk���EC�4�w�[���1j��%�Q�F*K��W����ں�۫y��M6q,�R�.eR�֩_y4��"��BR���=�p�$g:X26��o�^�l_\��}��l�r�����p�}��F1RLl��J��g��	����hjƠ`c}�3��mdR2����-K�T{yz�P�[�ݷt�+t��i�:taKꦮ�Wy�N��N{|�5o.�zQq:Tc��f7�lvzuU�IzGH8h�'5�W��7wE�C#x�����2ˇ�2���^�"ȋ�,昖f�<�c.���{�Гr� �c.�����̉O[]�R�K�]�3�Y�Z��j�r�s��9�b����w�>��T����u�ț%h�j:�:Z����̽io>X+"U�=�V�fv.mY2YY�͑I7��d��YKݞ�v��5Ã/Qh�^LR��;9����wz�֩
��S�7M��@��(�|��t&pJ�9[g�y E�+�e��5��yܲ#35��%5ݼ�Gu�Ȑ��N���۳�7o8�짢�͒�̷o���4]i�u&��Ae��ʭ�٫{_}V��Z����[1!���P��e
A01C&,F��D5fp�Åy��8��Yc�%@��X�41�b�`�bPC<�$�b�
>�/D��~��Bzܸ�=�o���i���{�	�jUoR��E��W�����g�A�m��/r޺���u}�{�fJ���Y�%��Ȯ�#��=ȋ�����]���֌�-Z�7��*�e�S����{^��UjWw,�U�OZ�o{3"��]��{R�_R��]
y�vcO��)DQb���ի�Iu�fɤ�U�w��.�nƼӡ��;w5w9����/�I�����\y`�+�%�¯ya����X����z��o�2�^۬���N��C6ye>S٘U���+ndG�\��O0�����y��	.��XO,����-ksu��M��t4�����X��:i��Yf7J���ݸ1L��RM�.;�o4��3:�`i�¸k;�V��Nu�Ɓ�RY�%-��RJ�=G����,�q��c/DA��T(�9�=ʅ�u�O!甭��(�n���b٭P���g���Ưm�s�v�V���q=�è�o�:���x���+�1=�J�>b;�{M����0*�9��rYm�Ir��lܣr4X���7;V�+��Es1vJ�N��t�Nŝ���B
Q���䢆�(((6̤x�
+��:�$)��<�OO���Ԝ{���K��V�ZZ[-�e���0çON�a�pq�B��5�e14�A�E�@P��>!�x!�p�s%uMQE%�IJDLQ]@�;fΝ8t��y��Vصm��i���S�Iy�AT%QE[m�����r�Ja�ç�N'��;��DSI0Py��ե�ImxS�����<ۭ%�d�EADV�j�#����9�,F���-U����[o�M<:zp�nqU4P������)����v�!9�"�a)��t�FΝ:p�{V�fg�n���E-�SAT������������w�����")")��f�����	�'ĔΙ�aBX�؉ş�-���1t�3����զ����;����rm!���o<���s��N�������@f ߟ���Y�a�&���nL������Th�|�e��u�L��3�Q}��.%�h1�,�c�u�J�Rep�orfH����9H��S6��B�C��g��lTan��+��B��`��f���G�'>�w�+�_CûBU�՜�d,��)j���hT������9g#� A��!E���o�:�p#�c�u�zn
�@ OP�"�Ԗ����=�D���ș��Р�䎰1��;]@��^�]b��Fkw�!�϶ݭ�'��H.ݠ9lV�ǎ4e����ݾ�~efc�%�EP�V�^����"�- �Ъ<���κ���� �6އ�g�ҳt�G,�/���a�[Vb�@l�8f3s�-��:�XSݿM��,��#SdC�����R,��6���{���e�E�����L����1t=j
:O��k������ɗΰ:�c�nѢo�7�{x`����g���<g.{=+<,�Vm5,I]��&�����%���ڨ4��Δs{���ݖ�j
B�`��� � a�����/,��+��~��^�C$�*[�v�f�-�S=v�!�N[`[�bR�Z��:�z����g�] �b�+�����+�Z�+�~��=�נP;3vo7���_`Gk�v&X�Q����`=r�GHYJ�fg_�u�rD��C/��4��-�"�?�2a��@c��l�p��� �l�:i����8��˞K����|�B������&S�䅛���YT��B���bmr+�97)U�^��Ztn.��/�Q$tTz锠͜�G��
�'�#� ܨƖ�z��\Is{���ڕ�{z��4����h2z���7��M<D�����^��@#"�('��Z'�S�㲺[�C߃�4��oK�lj��ɞMӍ'����o*�n�*�A�p������{zfw�E`�A��>���~v����69М���X��Tj�)�~��C�S�k.ܘ���Q���l���\F���D�Do╷9�x��U����(=����	#veح�]�_f�(�%�5I9�W�go+jbq�f��A%����*�� ��a��i�Z�gA��ݙ���M�=�bO`pp� 4���)E��ޒV�b�c��J֝�,c�@h�����b*�@�=<�܄��A�v����Z�����DF��2��cZ��g̼e�]���o�ţ�
�h_U�et֧!/f�}�A�db����ܝ�\����Ձ��>�Y���k!��뻐�E«1���'�5tw�<j��[&:���.z�[������QM[����M�r�~��ʌ�;t�}OǶX���P���ϟ�J���#����s���e���̍a�)�D�ʜ�rldS��f}
be d0D_1���Cy��Lw� {��!����|����w�!8}a��Q�a�.��刣2���@�)4-T��qŽ���{k뼧��Q:����^��%����d�S{x�e�TԼUHe��5NNz�X�y���}ָh���itG	��������霮x^�Q%�++�Q��U�EU'��I��
�;v�*��^a�Cն��-�w�c�-��Ud��Z<k2��-���v���M�IHݻ�,>ǭo\R�g��Sgs��'��?v��j&j�%ޱy�~iV�V�����W}kE�����fl��OەS�u�L\9�wI����(ݼ��j��7b.9�^����E��\���w|'�WO<�V
�	�=',G�͑��9�5&�^l_t��#���'�_*�f���]|U@�}�Kq��m�|���t�9��R{�_�#��OnerS�t�
�J�X)�}&�gwN���߷��WoLAJ�PzjFڹz�L]�Kn�<A�4�W ���D��9s�����D{��Cp	*�hf�@�!�rӶ��t�y>��]T��`G\���c���y�`��!�;rٰyo��������ۙ'�Q��*R�@{� �@z����Ai�7Yzo��ٮB>�_͏����m0/�}�^�x23�U{詽�WZ^�o�GS{�;�,��'�oY�ʗ�3�&�9]S���wDtp8v3ԡ�WT,����0h�A(@\pPl}�0�:�U����ْڱنA��9t�T���G{�S�V(��ĽZ�����eZN���1�9��ՖL��Ş�Xv�7�,�ޑ���C\���P�s��9��}h)�i����	i���7)N����5�E<�0�Ykx���N����p�`,�7�9[b������ wJ�<�z�ݜ�gl��	�ΐ���p���uN�8Cܱ�&|$:���e�\��,h�3h�h������7KD�Òi���� myTX�X��x�a�^���&���ٺ���`)�Q���D���$Æ���S�Wq �V]'��j��k�����tR�:��p���Z�f�)��+��,��r �v�m׏���Ǟ��w���5�B]�y�@"z<���Z=��!f��>	v��8���j��[�M�r����M�#�ζD-�
�7�z�z��s7	�^�OP�W���Ê/���٤sV@)���N���Hy���U�NC)pỐO+N*�N��=�E��	���<be��(־�.�#YF昣۹�U��'�TMQ��F�� !�}�,�������S�7�VTC��1���s��Υ�GJ�.�v퐕����^s*������>�����̲��>̻����"O�?���x�I�f�p����?�ʹ�ع��a��{p�9�0��[��U�h���'��>�`��$۠���2Q� J����>��40�-����m�ph�% ��F���7
����^��U�3��a��;D�WX�-�e�6����C��⭼5}��+;O:����e��W�t��`Ǫg�6�z0�˗X�REQZ� ٭��P�sSty� f���)<V���*ⷢF��ޛv\.m��ur�|�m t6d�ds��ht��8S�6�L���]y�=��8�:m����T���7�U���g�L�<��p�^\�&xB�b��M�2�vV�48��U�W�c�}��]כ��D�Z7��ؔ�$;Z|D���A��bh��F
��l�E�@{��M�4���-�w6���Z���t��yS����.Y�������3���=����c���e���������TGA����v!b�w��"��D�����FH�ڃ&?X���E�M���(6LE�|��FsRV\�<��ɚ*1cE@X���4�V�\oy�[�c���*OZ�(з��p᠈ [L�[�@_�6�*���X��C��\'y#���Y�pWJ�n�=r��4@�[&�'����T��CA�V��s<>8y�J�[�;�"w�sg�l���+4!3���nqp�q,ür25ݔT��F����>���3�ţ��[wJ������ik�Q�n��c0∾���:��`U���QR7�V_���痪��;�!�k����my�� �_t�WLB���*p�S\&�p�1 6��&�u�mT���
A�4y�����FIjMB�R6e[��`g�[����ᐋƃ���A�Z��A.�����]k�UC�/�>���/c�"Ƈ��<X�9�<<��^��j2�&p�}0Jؗp̖f���AJ�K'���24�L3�C=���c��{��O�`,���z���b��h��z�k��%Hd��oVC�M��u����5�.�szۺ�3��n
[�i�r�Q|�����T3������$��h�˭-�
SU�;\lX�q>��(t�9�me_v�Se;��u��#zH�����QI[n��w�e�S|s �G����aTͦ]^�>~w�� ���nVe���L� �
"d�0��}VwA1���U��~�/��]K�y}p�U�w�
���M-3D	�3?��h��$���0��H߉{���_ߜuPz2��i���M�1��홪C˼W��av���N ٲ��y?�$
��A�l��|��}���5�D���w?�.��(]b���q�jqel�t�M���ى5d���Ɔ�3��B5Za�����T�RՊ�#X����:��r����x����Lb] d �s��"�4j�ΟWB��Oum���w�UU�_7�����k�.�M0���`R��k���u-�y�O���\!�7ݻ�;��Ϥw ��d>oH�J�����\��z>��^��Z�;_W,ذ�0�;p�]���*���1�R\3�������s]�gQq�^u���Z���pp"	 f���Vw�*xr�v(!�M☎�4VcM��Ҳj���ą�3(f���� ��]�ǒO��a$_���q�H6��)�q��&��c�7!�8b�����T�wջwo{��EG��-HvxTmc�������K���q,��U��6s�~�qTձ�a���8L{{���h8�>��s�܇�YIo3���nD$fƁ�6�.�Co��0
ޑ
�����S��]���)7�}|�p������7��H��G@.�]!d�"&�Vs� ɞ3y�b�#5�\(��O�F��Os�f��({�15SU��r/k�I�=&�!��gF���nF�ݧS޵ �oؐ���*��:��,f<4p΢u�筴
;�T�Zj�U�b��.���)�*�tMa��,�Q{:wb����k�(��r�x��*����������3�WWMz*L��F/b����D�H���:�Ԭ�ɨ��S��!s�-
i��4�Խ���S���B�wXVA�1ʴPy�+2�ְ_v��[w��y�.��,�1�F�(���A�h ��.5�u�T�ga��Zi\˫5��C��$'Z����V �Zڷ�{�_%�qz"Yz�H�s����<�gx�4Yߛ)�q�n�`p�(�j�t�ޕ�U�W��O�P�˩9�lǆ�Q>��r!\>���"����H
���;#'#��D�g�7����ī�u怅�N	R@�W��t�A��K�ez!oO�	E�ǎhq��yV�=��Ga�ov�4;�WР,��n3�j�	l;���2fzi�¯S؀�ݳ V�8���q�/��{}ľ��\-��FVoUɨp(	�:���l������.k��NǸ�w��\ջ�C֜�Z��8Ŧ�fלml�+2�g-��k{}�0�M����K�:�����F����8'}��)xl{*�4��������ȴ��j�s#Lk4}��o�1.�5�
;b�U7?'����y��IM�P/� }�t����ۻ�=�����;��k}��������UEs�  �?��h}������Lt������1)B�0�{��,�\IPT�(,�	

���I

�E$"����z6�"(,�$PPn�FĄPX�B��E

B()o 2D�E���B�

BI ��!AQ ��!Ad�
E��!�hAARA�A��!Ad�
��!AR@���$�y�!IiH������AAb���PT���$�hYf��%�%����$�$PT%-�P��IbDQ-!��ȅ�a%D����J	)hZJ$��$�����J-EBf�PY���(,��I��A`�XH��I%��!��`�  ����~dǋ��
*�B �A��D������������O��}O��޿���?��'5�/��c�	�>���>?��������������'��?_/���|5����g�z���DUE{����?���P_���qUU�_�_�M�MI��/ޯ��`�)�"*�����������C=���:�O���{�L��ޟ��CD��P�R�Z@)@fA) �Q�X�hbB�Afb�X��F�b�V�ZE�I$FIV$X�bQ�dX�`�f�E�$Z�iHVaZA��VV$!�e�a�i�E��X�d$!�aaZ�YE��VE� XBQ�E� ���fDaaX$ZA��a!X Y!YYdX$V�bE� YU�$X�dFE�aHV$X	�a!�b�Y	E�($X�`aZE��d$X�a�hVdYa�h	��b�ZE�Q�ZE�)�@Z�F�hE�Zh(Vd� ��bQiE& Z�ZY�Y�i@�D���ZPB  b A�T�@�hT�e�U �F�P(T)�ThE� �T"@bD(D����Y�
P�Y�Zd�P��UZfAbQp�Rm��~NS��!��H�	�"� � �>��M}�����JO?���������}��z��UEq7��������v=}"^BW#��b������??{�6�R��+ǲ"�+�T�������XE��=�k�	EU�IL��8�v˸KNG��l>.A�l�a6UEoe?����"�+���t4'??��Ҝ�Mr�����C�_4���\UEx���dETW�'��3���$>��l~�,NG�s���O��v'�I?�Q]��	%�����B���'qԝl�״:C��	E����&�}�(����y��?��LS�?�b��L�����Nk� � ���{ϻ`���Ó=� �/���UV���5�KY&�m�I"%��("��M[dګm�[ffڭJ�5��ki�&��)������m�lb٫-U���)���$є��̋MJ�!-�����J1���I��Z
P�Rم��=E�p�@��d�S	&l5��FVY�,�d��6Ԫ����9+�Z��-5���[b�kX5i�5@�|��Of���^   {���ݵ�n�����T�շ]�m�s�kj���5�VfZ�ck������k�+�N�n�ݻ���(��tH�n-\�@��z�zԥZ��pN�9J�o� �)UJ)I���".��w��:�� ;m���UvΆ�[]����Nnu 2�S: ���)R�OwZ%�Mx ��F�SڵP���p
kj����������6�A���@;p 	�t4���B��(��� g�h ��@��]F�n�ң�c` w,րW`j�p�;V(WF��P�s�5��ڪ����°�h� |P({9� Wje*�ͨ��8 �8(�s@�`�۫�P#f�$]jTEf�� {݀(G������띎��ѻnʀS��J&����ĖU
�
uT����V�F�����l��;��Ͷ�ka� {�J�
�7��s���@w@)!u�:���8 5�8*U��B��Gs��:�s�JSV�3�Z�� 	��N�Ӣ�h��UUEStgv� 3s����i�ٸhk�;:�������( ��u��
��G��U&m�m��L�� �؊�<��ٮ��gr������m�:��P�j�BWq�)B�굶�Gwr�% ����h
�"��P�U֬�T< ��(:jܙª���`]m0�[�!u���E�\:]�ENu���s�m�]�m�] ֛�   �
�@ R�����#��#F F�����i�RUP 2h     ���%*�       *�	*�F       �#L�y�LI=�1�@ �	I"4�FSF�52 ё��z��>��_f��{;��c�i�|ݛ͸o7�D�ocW��7�AP=<���I���O���^�TD@��N+��G*
�F�_/�g�����c�]��I� �{
����!�xP��8���]�r�/ J
��x7���o~ݞ�?�۾���|����pZ�<`�N�U���k�37����J$ě�2Ҩh���%q�e�w����!��ʐ��i���n4���&UU��Q�-�9pC��Pd����M�4X�i�aqT��4T��*�V�&�LN��jU���;jR+dMQѴ+�PD���Դ��me��+D�L�GEM�6Ԫ��lBLn�[�9Pi"�I\�*��.gw]R=���ӹ[��5+����s㠔wSa��ubҡ���L��!�F��"��NS�p�IKoi��)h)�j���� �`ղֲꂣZ��T��ݹ��v� r8>Sn�@��(�U-S:
:�\kqI�|h�s6f�+���愯nV���eT-Rk�-"�n��.5a��P�����64V�w������;7��8^`1$����U�^�#�j�;f!qn��mfcP�f���e�K 	�w!��{����K ��VX��i20�ɑ��)�fd��J5��lv���'�J�+6ޛ�2��E��m�e�B�"���i���V2��[�j�JK[1��"�;
�*�)�	����mJI"y{��F70lh&�jV�4j��h�WY�<Ԥ�kX�(�O*�U�)c.��̦�	���"]��[X7G�Jw/�H�P�Ы��(�nҊ~ڲ��	�ha��5&h�h�A��{5+jóq�s���G��yv�F�jC��`Ԗ
M'.`��g�^�f��@!2�Kʹ�n�+l�!(�`݄���l���Y�=�Y�����r�ýZ���t��͊J�z�t���*
x�6�9��p�kr��mVue�۩q".��("P0�)~Le�	3sv�FX�kᒶ'�hn���<��kD�2�ք�>p� +��r�����Z�/%�q[%+`��K۰X,��l[��q�YW(���Eւ�Մٓ0է6�%V�ǗY�l@4-��
�iVJ�vΕA5�%��l*����G]Muv7BQ��n�fՊ�RI�i��0$�ǛP��hqMD��`�+QYa�@���4���Wn�p��8�%*i(X�w2e��5+pTm�&�x4x2	J�K��SNV]���kD�Kr%X��qMF:_^ �M�0mV^8U�j��&�쭛I;IZ'(mP�z��*M:H�F2�Րn��z(2=�){6�FVs���*a�j�lo�	_k;�T-��R��F�l��Yn�-Z2r`)�	t�Jfe�O�������K�4�ɺ�\�˛��������St�cP�)Qd-Ȳ�=J4�]�r���Fډ��,F/fXϝ�Z�	f$�11[�9%e�w���6-�m��A��T���cj�R&����fW���v�k�����݋C�r���á�ԧVC�!��7�ӹY0L�EPe`8RǧhF����nZs�*�,�r��,I��Ä�P�/(�:Z`u���K�Xi��7�*�L��ܰ�i�h�X�UL��YщcmU�f���l�l M�;e�m)SC?�hk���3m��۩[��3t�c�T��$��	�++j8�*fa�y�L2������zdk �b$�+�
ǋ#�`t)�����n��l�J�x�a͚T#W��6Ac@�6
7n��f�:A�:*�hܧD݁5�75`�3KҘ'Y2h�oN($@Z'5�9FMwLTLA ���ԯ鋚ve�.�`M��(S��Yj��R��eg�SMn�&�k��������5+��d��O]咉�d�� ����E6N�S(V�V����H@�FC��.��/.6a���tFPrIP��S�ؘEK�t��=���Ҙ�*&슕�5kb��%� �E��F9Jʿ�]"��z)��[87�ww#b�eZK	�
d�ɎR-ncP�x�nk�7]Z�]\�զN^���Zb��f�å��R��N��ti���&��ט�]�4�;��!�ӵF�.,�3Ga�nլ"�6�È|�#��hA�,��
��%�� ���BJW�H�Tkn5$�xkG�^�Υ�6��񌙷%'.���͓6���dy�eY$��.���藨�Y2L�H"`yYt\iF�Z\%Evq��i�L�WbKJ�mc�,F2�yfe˨.������QR`?nd�
��^Ył��2� T٤(�:���
�̫ҚǱ�ُN�F*zjYF�ŋ�S
��b�D�i�!%�jXq�լ]�%��)L�PI)�4���fķPK{����$�J�aWs4X�)J۸��f >�\����j�*[V���[���U�*���;�9vN2� �Z.��%e9YV��.,8�$���Y,n��,��#����hy6#�LnJF��v�c�6S�	wa2�/��Y���p��b�Hcb��M�E�[��,�C���(�f�Y�R��e��o	�V�Ekm��̀���
��ZZw%!��m��T
�J�x�&�vz�ǥm�2 ��π��:�qV�
��i��n���x���F�Ԗ��-5�R^}�fH�`�I�sB��X�Vm��f��Ht�Ǭm�8Y�T!7Mښ�I`�\����F�jF�ǓM�0��6�X6\�A�xI����U*nF�V\�)�JH���ʅPpU�;�,� �#�����+6��V�-ԬM<8��Y'�Sʓ��J`��ӈ�B���لژ
�����|�)U��ܛ�2�s˨,K(�)�����KY4��
��Z��Lű�R�f���8�B)q���쇃*��V���ܧ`��P9���ѩW��$�)޷��۶�!�1��&%^�7J"	W�����qZy�Dǫe��C����З�Ρ2��	�Ŵ�:����0�@�Fn[h�:�v��U�QM5��u���U��^��d���[��Old0Re!V��6��͙ot�C6/�s]H���bǬ���(Խ��7��5��-�ט)]<cR[�<�K2�Y�f����6T�Zl������d��He<gMӽ�̎��RV�=F�RZ���"��m(�����JQK[4�x��&dV���6��K��;F�˴"-�T�Y�H8���V6+]�ƴ���H���+�+n�TfH7�v��-�l4�nɭƵ������e�x^i�xৄ'E���W�Q(;R��.�V\W+sa2+u �6���FZ�d������`�2��m=����iPP3�k^��
��K+td�	���eG%[�(*��Q8�c�&��	���E�*�6�m���Q�5\7�X��@�U,�ִ$*���Yf��Q�D��R"G��gP�Q*(U�Æn*G//b5�2)men*f�jl u�RV[u.�m�Un�nFT{a�$E]Mi���fܛu &a�
Q��O<#cJ�<[b�_��\�[%n)%��&�N�8��4v+�
���3��Bm�.��ٺ�ړ �I�����{O>�ѽ̉:*6���<e�
^eFHM��]���k�z�V��&�TIk����ׁ�TE]��;�F㩪�-���nZV�
�ne���tlO�����Lb�0�YI�<�(�ցʑ��itV7%��nU�J�
;��c��ZG&}�>�*�:���or�	6��$[I��0��KLR����Xrƻ�*���԰�\֨�V tq�܉:L�ޭ)X�ʔƥv
!�E�x�c0�c�J6����X*�d�t�X'ζGu��R�&��i%�1�y��7Sp`�dYۉ۩���2��8�� Y���]��Mf�r^��ԫ�l���:�8v����RƩ`� j2���T�-�ؙ�"���m�m�JT"��)��*�m�*�,�S��Sluo�4��nb��NC`V�{��X�ڃ˕3mg%����TsKI0t�����c4W�XN��譲�[������,G{A,b-ʔˤ�к� 1"��M�.C�Z�A��f�ѺX���s��Cͨ�����2�(�$�ۢw7> ˓$�߳B�,�[����bC7(���;�-��2j
�z��1�WV3-��ɠ�����orڅ7q�e[�f�y�� 	DQ�Xp�Ү�P9��E
"�8�F��a#n��c�g��B�j���Ոe;yVAqA���T��H�	�I�(2
o~��ff<��`�wr;�����1�6��Lb=hVF����x�{��;�A��-l@ޗ`���f��FT�OR�4��u�g�"1����BV-Z����BWB훙���t�j&Χ�r#h����蝫�%�բ��Mh�1`�Tݛ��D[����v�)0K��[��wPV�Sl�ǋѲ�xC�Y�`�����C�+�lk5�1��r� �w)kZ��K��/$'&�77 �L��I7�md2*�L�vu��bۢq��8���l��^�Y�!x�0c��3V~�<�W��*~���md���ШV�آ[�ziA�7���(�x�"mZJ��n�p���&-,�)��Lܔ���&2����-7�$���9/^hOv���kгL�]&A?�a��n��w4 Ҧ�)j���[N�Z6f�䳏Zk^���Cytܴ0�F�K��pS��t��ڙ/p�q
�`��55'آ�ŭhY�9�mA� m�y�b���Un�FJ+QՀm'�Ф*ʕ��[tr���j�pӲ�ӈ+�bR�Oڲ&����?!�c�J�(|V݊Vw@�kTخf�r^���u=B�e�*����j�3��(l�����S!�-h��b�6��u���3VIf��-���9t4o׮:@4�I�d�!Vl��2�v��ܕ���)T� I��yXJ���Ie�UP۬�*�e�8�Qn�;�"�f�,�Y�����R!��)jV=˨i4�%f�zEܑ�(=P̩t+XA�N2��k��t�nIt��e7wu�������z7���xEj(c��-�GaWY%�f�Lϡc6e�BR��w��%摪8� c����&�1�Y-�Z�VMٰ;ѨkN�-mJ�5:e\�
�8��@KA��~�u���r[�C���N��eB)����/�6��NLV-,�i�i��k!2�Ǧ��VoT�X ưff:-��]�]$&�i+��u+��T4��vF�53H=$'P�:1&6���D�Xt7�,�U���~������w ��T͟va���27ܱ%f�8�em  NQ4��fĘ�����C]:�FAb0�;�[���[���p�u{3�r���  �e/�k��2�e�L}+q�Q�$_��yZ%��]M��[����e>�O&ޫ��b�A �ݭ���i���Y�q6멺ĄY��VDJ���Ldq��%+cJ�&F�LV��G#U2�V�i��ҪY,��U,cqBZӊ��)�i��cs.&�T���=4Q,4�T��T�mZ�%��D�Eb�\ ��q�r4��*�(6�BeNJ6Z�#u�+]��P�U�۵&"��J(�N�Q�!�)v��w����:��7};�U�x&���:39�Y&���^�݌�=�ǻ�*���K���m�k��ܫB���tL��$:���G'\1eo�+o�s��%�0�]yD�2�wROZ��X::7ڻ:M/�L]Wsz�cV0\���W(:M7ذκ]Ʉӵ�u �]Czck�Ųv��F{FԹ���N�ݕg��鳴1	��[�.���a)7z�U�.�N�`'�F�8�a�wK;Rq9�՘�����䫋;�]l�ݤ�6�B}��4IPN4X��b�#�IP%�c���+V�ǧ�N�t⠓���G�����H\㡱\�Y�W��g�(q?ki��X+v���>�:���=p&喐Sz����/�mF8�ү��j���=N�Pd�s��68v�IgL��s��Cp�Y@u�v�-�F�L1��d#r�;}�����]Gs2�r�����|sN���M�Xҥf�6�V�����Zה�Ҝ?�V_���o@���ȥ��V�t�˜1�R���aN"� *�E��ܖ{��o��hR9���&��7����4s�b����]�xm���J�MU7e��6�Al�i	�����T�Ѭ�S��;�Ң(Xo s�	����i����㩏��bix#r����
��*e�1�;fs�Z�{�)o3��}�S��vaV�
�{u��f4��="w,�QI7������Rh�E
\b������ l�=n�1fr�[��*�.Y��������#WϜ=�rd�1�zh�N��%�R��������x�j���P�)�v�\��3�|�oi��n�G>3���r3AY�*9e�F�ڶ�KR<��+�*�vL��t���������h�v��� :�U��s�Z�-fV���m���#"��m��Q��i�Z� ]9��E�2��[S+�T���z��1��m��`�tF�Mۡt�ۢ���V\�w5���6Lʖ�-�%�[��R�R��8�A�4�Em�&�EZ.D{`X�˛Z��<�H9����3����R<����������H?��-���dHy)�{G�xz��&W2.=}.�M�#����j�j�t�n�ُ5��C�z�)k9A�B�-}%v��}�m���Ĝ�r�]��+&����C���|�Б��d/��%p�j�2V����i���#[�-�Η�,���T}�[J`U���Ѭ��^���i�����[.���p�e� |k���qD�d9y#-���둁�[����"צ���G�bZ����£9ԫ��t���4���q��P��R��l��ۭ��{`��V�^�}{�u3W����&1����VHE�Fj��4#��.���01��e�A�,��Ufg>�uˉhU�I4�"{&'�.��6ł��Th㒦�|����uev����k���^��ʵ8&��_h岘��;(��wx�v=�(2�x�������X:2]�J>P�`v���[�����4�m�Y&l��NJ)x��.�kF��8�/d<GQ�q/j�y�P�tl�@dA��h�pT�
|`κ���GFy���鲵#Zw�u�ꏲ��r��78	*�EW�H�c�gkޒ�Ӯ1�k�e���$����W3!��k�e5�Q�j!��m�5��]x0���}5+]���F�.c���@t�
0m�#dy{.��PGz
�T�eB�Mmg�]jd�ڹ t^���l/H�9ccG`��:�2+n&�^��;;�A���������&T�K�u{ Z��uf�ּ<�i[�4�]��I���:3:� �l��X2`W\F��M�K��'j���W�nin��u��������ǜd��y���h�ni��S��� :���u��ft�FA]��1�չJ�� �dZ�:����X��m_��� P��|��WR�B�ȓ�sV�Eٺ��髽�sU椹n���gv�����3u�so�m׼���Y{f�(�AW0�hÆ�٨FZ�\����/H��u\�o%7�ш���;6�q\��|�h�5������oqN���7�C��̖���R���Ҟ�H��|{��8((��v�-tH�ko`:�H����w�Û�
N�RC0;�QJѣj`�Xŋ�W��G�v�ͭ�j�y�I��h����K��]�$=ʥp�;m�nj��]�)lf�ʙc��7T*��
��Q���Ԯ�`}�h#��cm("��� p������9��6�b��*)bk��i���0����el�{slf�+����e�r�b�H�I���ܨ�Zie6��+~�44��ۂ���u02a扭.�(��ԝ�T��`.�`��ϒvFR�F�̭6&"�Hr���-�����h�Www��lY�X�����Q�{��;�El���<�^�E\��0`���9R�7"�I�;��1�u��[G3(�pbrԆ�͹�V���We�%R/�P��#�.�������jl�,]:8�`,�l�y��� �;j�mP�]̵���Jӓ�kOd�9ـeH�u�գ�B���i��{���E��@v���n�w��/�Ж�Tzxe3"�ر�Py�����mAX3,$�K�HNѥ9�6=�3s�ۈ"�Tz^*Y�ƅ�0���c��}�����K��&K�hV[��~ٜo�`�W�uz�tN+���bͮ�D��5�ȴ8��}���=]�(��{y(1؛�Ԯ �����6NXD��b�7��IݢЖ��Lg {D��y�Y�xs�U���k_���n� v���\��q鉎�L�7������zP#�1�R]3�ʩ}��S�\��:��d���ב
u�M�DlV�{��fq��2L��s�-��7	�f� r������D/M&��n��QC�ռ�#/؁�o9����6���S����*�e�(�b#.�^�̾�Ů�	|��w���.l����Z�[���b���XB�L��;����}V7#���\){���]���er�E�l��6-��`w�y�,�O`�S��K嘩\����6f�B�R���*r)S^����Ć.1��NS�[q��%�<0�5_,��Xox�+�@�>���pQso'f�؝3���:�2�U���h�ٽj�#�� ̺�R9���Bs�����a�	�N�v�`��w�����Φ+�]�P<��H�G���ܮ��7+[�9�Lri�S;��ݔ,E�8fi�X��]B�g7�m9}�����;#[��<��w���Wɩ�J�eN�� �@ý�*X���4F�w�+�k��{�G��YK]�ڸ;[+��))Q�-l�z��u�cR�`�^6a�X<������1�]�J��/�f�e����N����䔩�a��r�Du5��5x���{���3]��q����j>�K�\P򺷹0*�YRsHTyw]���#d�Gu�h��,\־���U �(;�$�v��4Y��U��m�֪����C�%�����4���gm�K�,$Ӯ�)�򸳝)L�:�����.f���*im^m&�D1-+qh�J��e�dv�v�����3�D���2`Ü�n�Č�m`��; �rq/�lǫ����w����p,ڢ�>�#7��h*mI�ͻ���1pW�3nر�-���ߜ��⬺�e�^j�5�#^��!�&=�Y2_#�	o��<�D�WO�gK�O����˭��>�j2N��Nᬃ�u�(�SJ,���t�A�- ,��b+:u�=�����]o���K�2dSv�d����]Z��Q�9YlR�xub�)4����}Ϲ��
��id�p#�3//NG�et��y�ty�@��6�$��١��/��.+�,'k�Wm*���^I���.�!�	�^�v�Q���M��{����99U�,��� P�P~=�:R�W6�n��ob��T������z^��8T?[��9��	r�Z�D9m��ά�3����줺N+æ֜W�ֱ��(��[�ϸJhr�2�ee��ٖ���aa�ՙ�v����V�crڮ=}�	<eT�i	���|�r���[l�}�u9\Fwp��1��ռ��6�ն�у�N�r���7��E�e��0��cn�+B!nMQ��%]7��'�۬n���8��P�IJ�@�frʾ��gi����v��o�Q��B؇�6��yl�ʬ�].Ҹ*9N�Vmñ�it�r��NS�ҕ|h�R��v��y(��q��[����m���1�g�]s����}�Kˊo��7Ah;z��okL��)�*��F�AAo�Zf�vJ�}l��>��yO-����1nZK%´f�&���׳A�5�s��D;�����`O2��w�L�f��݋ߞ>���}�Rl�y@���IW7w*+�99��2t�9à�x"ݡ�
��A�C�S1�0��e��f�m��Q!Rں���"�����|���<Ϸ�����%ZK�r{�o�
m6��\�����&�ʐ���.����h�n4�/ ���.aޜON!��ү6i�u�۟�v�?�����d�jrFvN�T��Ps�F�[9R!h�c�;:ķ�0�K�G�;�*n�|&�����,K��N#݅\Of�S�és�t�n�]���RٲgrY[���p�a�ib�5�˅�S��Arsr����lS�$d���Y�;��)Nқ}\֪!�q��U�6�s8V�n�F���e^3� �T���|r�N·��m����ԨaeJ6.L,9 ���=t�T�D�\E�ZWr������܀s��Y�pMU�FW�ޗO��|w��e��d��X�u�P��d�@����x@w���Js�[��6�N��EwI��u��n�Y�Ǘsj�U>���dv���;x�4�\%�C�'��bf�1�{˪+�d�2�<�#�Kޭf")��s�iA�ql�'1�x�I'I$�I$�I$�I$�wL17g+N=FY=]��Q��1>ϐR�����L����:
o���d�3��f̛��ӧ�C�ME��s���߫0ß 8�!7��~?Y��1�F .��1j�@���%��5���[Deo�HI�d�����Cl��J])�M��NV�g�dbݤ�${�S�z2�vfڛF�,��W��X�Z7m����d������N�"�n�#2ۊ��B�<��/Z9B)@rf��a�KW"�=ܑ�tO�p�[���&�Z�0�Ǩ�w��C*�/c��a~���tEU��ߊ�����>�=
���p:q]��|��ץKI��i��}8p{L׋��ͥ8ͻ�{`vn�U�3��>;.���VOm]�"��22�=V��9W�j�▢��&��2�h4�oiR��[R�AC	*�[���1�An%�T2�ry|֚OI�6bA3T�t��2���E��>�hh'�W^�m\�rQ�x[\1��ց�������=e}�������k�oݦ� ������u���IZ��&��5�3��b.�� n�I��Q%�.͚CW���f��h�u�(��oC��Xr�⦆�6v@��q�kH�o^���2t�C�O45��A��:q�\��.+pTư�u`]��)��	V6����J�[̣��b�kl�F�/��!I�c,]-ue��5�Q.3�X@f�mW_Ɓfn:��k'm]�4������uʸ��u�ɕ}�J�8�ޕ���O2�:��)�{)�!��^���J�7���&$J�h�p��j�RU��Sh�m��X�Iv����޶۝�X�\cE�}k�{D�
�@L��\�\�vvH8�� �RrI>��5�Q짬��ED���r뙣�h�\sU����B����΍�8�,��'�<ĸ�Ë 
\��!����o\�z�wY��Aƌ��R}����oN����:5V��e^�p�@_�i� ��O���7P�K���g^Sg�Gd+}$�ot�t��#�*�L� �\�F�Gy]�u:A��!�*���S0*3�y��C�HfvѼ{@8*o=����j+�N�8.��r8����k��>��8k�[N]-`��i�ц��'��QzFK%�S t�������	黴����։#*;�Ȱû�q\�I��	�q7�e�ݾRt�V9nt,����ud��%{����б�T��1��դ��:�`
wCvq1���v]^�E@�8�;�W��:-	y9>|�#Bv7x�oWvmuoY�)��\��L�����$W��)�+7�����7���w�a7���5��q�K�����Z�r��Rј��>��Jw���h�N��#F����ng:X���X�dӜ��IV(�cD�{���ڷ�M�.+���Y�Z0��A�(����%�xu�_*2�e�mIA�&]��+c5�e�t���rxxՙ1B��V0W<��Eh-�ŧd�G�t�981�s9�(oB�(�Hj�&������2��Xon�$�^t�6D��� R�KVR��z��wM%����I�}r
�����\sqJ�.��|���A�*�#=5����C��|b��}|&B-nmF�E��v��i�vkf���;�m6���#S7bmPw1db�K4w��2���KN7[�j�؋���V�,��]@�-,�q.�F����d�]�C����iP��8�g ݀K���t�7r�n���&*�X6���o��d�tjR�I�#�5�[R�U��d�.�a`L8���ѫ])��f�1���Otei}}ch�A�����w�#��(j�[[���,Fq�x���i�����*�j|�m9�qJ���Byv��Fu`��]�t;vq[�\��?9�l��@�I��,K�Ž�C|���y���n�w��L��U���������,��j�ۉJY'tv������:J�(͂�Ҵ���ǵO���J����m
T�Rv,]ۜ\�܋�EC{��+B<��ѹ��@���I�Sv���Z�[�"nL�ź8(\SXvZЪb��a�K�bb��5@�UaX	���]t�P�
�vau	xW0@�7�S&p����pݡ��Z��R���9�V���.B<��C�Qf���1Ԑĵ��0ֻ̫v8�Y"���}6�ZZ�� x��V�ƶ���KX8�t��w�����)���ݟ�N�6���H�)�<��jk�r��Èڔ��|i�Nf�
��[U�0�t��,�L�����>�;¯8���W���VL{�Ր��p�(U�M75���nӋ8�d'ی�Ӗ��Hp��c����M&�uF�Г��.I.���w���B�[�ჳ&򇄖��ǐ��{��Y��l�L`����!�c�"���͜��*�Q�ׇmS��5w9���5�t��rcܧ;���J���2]8x��jk�9��n�0K�rP��A�[����[����F��wZ���/���/�����,u��TT��Ox�a��\�1v�K���)�1���"Qå�%j�)<7H%(�k{h���
+�D&Bw_P-��Y�2�K�V8�ؘ�0R��N��{:b<�)7l�Z�퀨s�[�Xl�rr-��<�1a�}�ïV1��Y�e��*.n�t��V��7��g<��<
�U��u��8�Pc����\�Q��:�������e��ѫ�O8�
�Y���/�.��'F�fu�ԫ��?}�SyյU���1�ˆ����8�B��+�"�n��Һ��W@A��}@����RѠ��fS}z&nnVN<���.�i��]'c��U�b� ( F�a]2��~4��
G$��T@h:�d�����K^
�wH���=pa
��x- �}
uur^�*�WM�*
�C�6UX����ԇXQSP�j�t�_Q�Z�P�i��\�w[c+9��wҁuB��ȏq6��Yy$���c$)j��F6Y��0]��7vܩAbZm��G*�65�3)��*]�~��껩�4��f����9n�W�ғZBڝA�)�(��w�M���3颳tr��k��K�}l�������Ԝ�uk[�K���ٛ�"J�.EU�m=���U�Vvg�DG��oFQ��|�����t6��U�"Ѯ�}۵�%��������^|�޴�P-U�C�r�(���2�I����������\�=Z���%浟 ��5��H���y�_)b�Ey+�Ww1��x�zU�V?ڞ�V�1A-���(4��1hYme��� f�Y��A��Sb�����v'����P�l�֖4IP%�X�@���5r�&�(c'�\�u4F.��c���ElU���Jh�pr�=tE��@L�c��f������5뿀b���fE_�u�hqw�=�S�eٛ�K�r���Sy|�z.�a��r�tk���%u�Vj�@�GaP�:��z��f�&��!��ٜ��#rC�X!S7�pۧ "���#�".?�7�6�]ʉ΋7��;UK�ZwP��|8�Vwym ���~���b�J]n���C6����(��Ϛĺ�R��T�;�(l8�^4`�"���`oc��Y��R�C�Q���<wU5�Bq�V2}bbٙSͦ�|8�ԀEυ��R��Ɣyٶ��wWƻLW�2��!_�GHJ`�[wOao�}��*ϭ
��)�W,Qfwq�]7��c�
�;&ۨ�&�uX�t5�6��Y>�mT�w�ԹNyf�S�g��t�2�6B�xs�����[����7��I�۴�
���w�4"�
״%�u�kj�7��	�WK��$+#ݧpo�
Bn�vZ���a3�>����Fr
��̝mìU9[�0��yu�٩ݵv��:����`�z�R;��Ŝ՟֧f�u����������Z���3�C3v���S�S�Zk���ߟ]��./��6��ѹ��R�-�Y'�).�S���C���������lvP{��UōW_R8Z��w>��_}��GW�,�˧��:�Ca�2غ�U��y��i��-�>Ă�t�lQ�P���X��ň��'ʷ�Hp\����K�AᚥN56G���+B�AH%=ƺ^��z��+	EY�U�-(�k�����d6�����֌�
�z�\N��w%mҢI�Y6�Q ���Gqm'�8(S��8.J��
���i7O�=����������7{�^�7l�@ �R��n�N�T�&2�%�X[�|��z����U<R��#@o~��>ʕoI�Ī��]�0�t�����XX>U,��llV�Ֆ�@'�,��N�ARu��6Vؓ7��YRIdL�f\]�[�57�Z�����Lf�R���V�Nu�a�%v�(�q��:R�!��R�V!0�k� ���5k��2L�5S��Ȁ��`Hp��e���8v�Gnb�R���XZs��VAH���B]��5��'m�(�+`1Rf|6�חi0��.�R�N��8n��<s.�&7���9�WF����)z�)P4��o�عΕ�Uj�b�Gw	��L4�m�K�6r-R�fA�/�n5$*�(^��O��,>[Ӆv	_K2�<.����i���>5U�<a�8\���8.=Gy_�Œ�:*���Z��!��k��>�j�l*�:���������k�� ��%�N��vɊ��:��Tķ�R��Z9��V�Y	V؋F.Q1�=� F䬲j�Q�/9_q�3���Au@��LÕӏw,�2>pc�F�g5}��Jрg �˵��f�4q�"�j�">�r[І�δ����9���i7m�{l�k�����4>�]
�o(�5�_�|���������<bl��</Mnɢ�����{���p|^M&�8������Y0��ȓ �.��u�otn��WHPN�IӾ�&�����Q�ĄW�LUpGE�i=���'[WN+#�Lx	wL��'�wZ
�-��M���d��p�]���n��˱�G0�c謫2>���Ń��r�;3�9&�L�Mh�
���E�X���S�ĝ�P{�d����:��U&{1W9�"O�.�9e��Suh�;\_$���� ́�>+%��k˕ ���u��%�D� �#�,-��ݖ�j�3�A&r����n�,�Y;�ͭ۽v�i9]a���Ɯ9WX�	�^)�9�Y9��g��\FJ��{�+AkiG���������"�x�ٌ1�{o�2me+oа�����N߇h*���K�#k������h��ҊT&\�k^k�蕁[]�+N�-�M�b�XNZ�ψ�#R�4�ë�o)���t�|b��޺�M�5.�2��Yը�ϳ�a{�L}/[93r��,D�˱to9��=y+l��2ܲ�A��"Ou������������s���u�����q�+�"�.��X0�[�����]:W7)�՛����Σٔ��{���a$K�5+,T��V:��m��=��('E�/k-�o�+���㼆��n���pM2�i��kw�t�J�m���ף'#X���9
ɲ��BKW��x`y�u[��t�ń p�D�����Rl�ͺ&�6������'��&S�}���o^�cf��:��\D��������<y�����Q� KQ���&R���'�nv۞�u��8I\R(�YdU�\po���V�
8ޙ�[jW��R(B��PiҶ��eb��U,��4�b����U���?X�­���4�E�/[;rI�f�ŋ��p�Ƌ�ׄ��-0Utݡ���-��f�>R����ũ���צ�ܒFܩ # y�*U�����Y<��;�KAS�q�+��j�=��A��RM>/W�[�D�]������(����c%7/S 4�g�ԗ�6�a�f-Ȼ�-��u`���wv%�y)e��{����*���ާ6N�f�P�}] �
���J�5�wf�(nEumL4��R
�s�$E��T���ɠ��M��Ja�+Oƅ&��Zzpކ�����{D��T�K:#0���uk�����/���l�0mns��J[���`����ƱY��2�u2�<,f�:ʈd'd����Ӛ��t�#E
î+=r�L�v'*�!�vެ�qv�&���.�oR�s�t�8��0@p���z�*l��;T���r�.{"�S=�u�v~��� >�>#�4�(+A�l`=Jh)��dյ:��k��NHuP�^��h]��Ɉuu�i4��Q�h]kBhth"A��4$W,:M��
4i����9�r]͢�r�3EE,�QT���%Ԙ���A�QE��)�4P��D�1,T����ll�F��B�t1�m��t;X��"���t�$�3S0�h��]8�j�Tf�*6�HR�4<��!�9bmY�4DkMm�օ�i�4�\�'��#n@��a�s&�f�#l�� r4q$DDF��\���[d�h��#lTT��W.A1QM=��d��*:� �Z�$r�=��-���<b�m��l��U�
�6�N\ �<�:+�F�nb�9����r�sA��m�ACC21-�-�$t)"mMPR�CF5�ګ�����KkJ˕FLL��z*��~"��gPy;`U�����>�6!{v���k������P;� ۼ���R5�X66sS������ŝ�4��E'�@�����  �Z�Yh�+��N��oc�@��N�˄.��x�A]xK�� �J��s,e��B����I�����b�Te�Gɓ^ w��H��4<5��>�SI{e���3�:\;!�Ă>j��J ����Aa$��V6��K�=�n_��;�Ձ8�s�^A�<|�
�́(l&�ϓ���[�Si)m���ǅ0��/�h
�?y�~�Q�=��%��Y������ɍ�4��VfP�V�ar����lR /H�y���j2�����3�*g3W�ɮ1��8q�~�T��	;�b��IM뱰蚿œN�fY���KHt买�T7L��O�V��^0we�ϴ��?��j���=%���Q���[`Lu6U�9���{'ԣ5�ly�������W���ɒ�v��/��T��{Fd���4
��|�YĭE	Xhj��j��9ZDF�f9�%��f����A�� ��]1�6���b�C�aa��bT;\��l>�Ā�O:�����Y�٧(��&-���1�假������q�^#��Å@����n��z*eo$� ޥ�N��vmN]���cO c�t-�1冴��-'��J��Ƚ2Ѩ��JqA��Cqؾ�=�32�ױ Ə��U�8�u�D:bM�F\8C��w�;_��?��ļi��i��5�0�_�f�� �g�v�"��$���Q�Ka5���4�v��!��F®(����a��W��i"yy7��M�R��&i#� gyxz�^����[�QႥu[7������Zc7��sz�W�C�jɬ��R=A{������hd�]2�-'$�y賻̪�8�!�{�
3Õ/�+�i�v��t1@B��D��<�{˽��	8�����q~9��h�]�. /Z|O�z�S�z�Z�d�=�+ת�P��ϼ��x�C6]&P��& Q���K���^+aS�5�,�M$1R���m糷:��y�u�����q`5zz�EpN �	]+��9Vwk���H�7�
o�E��d�mC�0l����Վ�{�Y��)������>��tR����0q����6���i�'ְ�m�4�+u�CvK��	��8�,�Ы�QU��V��Z�gn ,��o/��gm˞��E���Vi"��`fQ��6
wf.���P.��ZX��U�/�=�I#ۺ}9��j�V���&�q��ӹ|��ja@�6�r�X	q�Lȋ�U��{���(w��r�'�}.�Oi��SL���n���?��T�ݑ����\�*1��?F�}�g0ݚ�����V^�ꆅ53�W����u�~�&�yK7�6�������:���+�k�V[�2��+Z��맷���$L�+tށ!D�O��LKwm��Ɠ�i
��B�`��?<���aCp�ެ�4Ac�-w]S\��<4��(��>V�yt-�ޱ'�0}�4��%顧��������(n �����b�rtp��'��O:6������W�0��R.^o�}�fF��g�l��-G�YMp��wię�5+�I7��F�o��VS�4�^��6v�a�G��
�S �[���Է�H
[��ǃ�>���ȸY>^X8�*�W��˃�hξ��sh��nda~���F�g�*�C���\���ub��B��̫�N�&���^�2�"��������f��0�v����x���m-OCc3��e4R���⏆8�A:(XXo�R�m�&aޅ�Ϊ�����D����^3L��1b�lqٱ�Ҕ���*}�7%�j��A턽�e�W�|i/�;�W��0��U��u���ڜ��yW+�\�V{{w4V	��Ã���#���x�� pC��K���]{�Cs+�_-��8�`��V6-t,��<e�^$<.g��i3�/-�������Uib&�\�b���ztO�~i�)�׀��ˏ�3��.�|r��@n�r���m�Gհ�����i�\U[n���@.����r����(�D�Y�P�o
F�_�!�c���d�����w-�[JŇR=E�D���B����ة�٩��!G�nʛ�j��.�_Z�TV�؎4�u>In�T���2��K�%ə1�q�<pE��B��)�����,�{1hP�aW�
��#��B
��`n�T�^�'_�y������Ƌ�׊
��;^�[���֖�{�n��w>�0>�n,���|!<�y��;ь��5�ǭp�w�Ɲ˄T�Ypz������3:�G���2�Ӯ0��ݠ���ޖ1k�:��q�w�U��H�d(Ϡk�P�FY�Th�ǂ���V߼�ʭ����r���g{ڷ�n��Z ��O�~����^���"�ĢP<�H��~��ƅ
Z��ǫH����H|{�Y����<$�n�W�B�sz�j�-(c��d� cN$!6��x��6��W�Ob$�� K�ik��۶��м`�8��b�7J�f��������}�&���z���hL�&�N]\�n��Z3�a��9p.�hS��5��!�B��L��,��f�p���OxPgt{5�4�T?�������R���縺��]�o-����茛�H7����Nړ8�����U���ƹ�s�<Yf��b��ӆ�S�IGK�����s��YҨ�)��]�9��H%��ٰ��mIaa�$�H�*`�7�>��^f�q�����t�V`<%<.ax���q�
gw��$8�T��<ix���+����
�n:Uye6����~d��6��+w|��}i��0n`�u�K�u�u3[n
����+'�E3Q+u3$g	V�v��^NS�_i5/���U�_}n�^Y�xcf��t��͊���H<�S�+�^�f�w�K�L ���=ƞ4:��J���Pyg��m�ѱ����"aS�'�l!Uv�'�f����ʩ����q������K~����`���u�s��LY�U��'���`�n�i~G/~N�R���5�q�N񆖻�ߺq���^���3c|X���P����������;zC����v�l�5~<�ȁ<H���y�QxkGi9�X��;/���^��{Mà�Y���nc8�.BD<OZ!SΙ
�Ё�έQR�n0��O�b���Ю���u�YIBKvd�u>��ebxwB_t�k{+�j�e-�.^�¶�+�P����nK�w]؆�Z^�gs	� [8��U{�;�mgd�m=˫S��55xS�V�fX�I�'t�'g����u5��x!,A��R�S���1�i�h�ɠ�&��\�wD�뱖ؤ�������S�u�YS�dO���Y��T�
�q.�pP^>
G�-/2�[�7-��(�2��}t��0�u����G�t�u�Ӛ"�5[�^�ԦĀX�n{���v +B�&��?Wk��tX�¬i0=6{��ԅ�2������lq8��܅A�ZHT)���0J����kLr�Zp,�I�y�!��x�^%�1�"�M��^�OR�һ~XU9ء
9�s�Rs�z^��J��ܔ;�|�ѯ��l��F���ӯ�p�ZؗI*�t1��<*-��2������PH�o�4�F\��c�W��}���J9d�e)3~;�*yeZYZ�k= �ыm�*RF�o�HfET�z^���$�^z�Z�Ԯ�\��; ��>٦�8L9g�a��ut���"l?��u	;{;�
o��a$ӊ�N��]3On�,`�{6d'u޽'�ӨfӽbZ�p�i��W!�튓3)_*dO��9G%�хi�R�G�����MA���,|teoZ���,��8����P�o���͹^��
/WE����Tz^��e#���~�����z�;X�7ӵ���Y!�IW�A��=>|`�W���(�m��h��������fClǕ������olr{�}y�N[U�	@��О�H�#A�qL)�U�.���m���,%2�c읁)�;䆑9�H�MhH�h�f���:2#	ؼ�@�� ��G�Qn{���y;�1���5�B�E�cT��E�ѧf/Q�cM==3����<�ʭ���P/VN�!���=��7H�� ��MC:����ں%̩��e;�m<�[a*L�p��A%K��^od�����Y٩��m��?�[�
e��Bh�Ԯ5�v�]�%��]��	��>�������v?v�s2�V�5�r�����>��k\�s�}�:-k�%6��j�����W
��K���m��*|��;"�>!sYTkc�kH𠢽s��2�X<��L�~�!7|�t�-8��y��ț�U�:w�F�~H_�V�~�2m�n�.ཊ��T���*���C2���A�B{8*���{�8�kG,������Dc�Q��+Ɵ�=�=nY�����qS�c��_;�Ȁ|n?gK2h������*�%����@{���kNb��N�{���d�wq
�@ڂ��)�5����^�L#pόυa+Nk��mx�$��O�u�x�<��zګ�p�Y��@P���
�p��wķY���,���j��c����B�[�m�{{"0wPgm\�d�:�sx��;'Po���P�z�C��J��|
}#�Vz�{�!(�5}&q���H�ѕ�ʘ�� #Ɍc�ffޑ���$0�r �V趇3C�T�a���U�Vlb/�����yv��b�+��AH����X���}�U������5{OS*��2]�eV�F�3	���'
��K��#D�G��l��!$�+XD�כ*�,����;#+��بq�Sv��f�O�{z���^�2S�+�wO�/݊Olם�:p�;WeCjh�����=u�DqQ}�=;��>tk�b&f8��d�O �6SX{���\�˚�o�|=��9����t�0߃�K۵�{�򄀓�sZniά�'|c	��q��]�ɔ��H��ݙ��[��p���ӊ�b�W��dǴ��o�;;�VzB�v�i\]�6>\Vf�#m���L�k��W��S�mg���p�ȣd�Š}Oo{ '[J��`���)�S�N�X}�n ��N��/���}x��^�[U�-쫀rA�F+��*n������tQ��e��V��N�FֻS��\c�\�݉v2�h �33l:q�!y�i`T���b��Gh�����B�C't�5关6�g^�n��iw��сR�V1�,7�M�#ގ7YN�֪�x�����w�M�
��V{��}�:�M��_^���Ir��t9t���A��c�qv�7�\x ʈ��p� qg(�HB�:�I]B]	���$�ں�P���Rq����0Ԯ�܄�t�NF�`�4X=�lt�ۘ.#܉�z��5h����5��Q紎CZE �g����v���C;����nn�co����4�!2L�1��ُfQ�zk��=�.}+5�]�碳�t�أ����*Io#���h���$jov��κ=��}Q��i!�ƤO98f��eX�=��˳�sޭ2(����V��A��h�nu�`�X���F�V8M��g���}�W�i �����1Q`����6���� ���u=�He�Qφ�ݹZ�@�@u��++����L��j����Һ�D�@:��Whޔ:�=%3�[��-4�e	B��O_MW��7�P�e^�k85MN�MB�/�� ��អ�aZ\ϰC"BQL�i��pk��݁-���qrج�u��A]�Pɗ;#k�t��:,,h��\�lt�5u�]���C��zދ|T{ �z��HCǘ��W)���&��0x+QI�<Q�5^"/u�c1r6��/����)��ND�sn�\��w�^�v�6�R���{�3xp�+1�
�Q�ٳ�{����]�y�-L����[�+W>ucK�;�}�:�Y�
ki�w�u�i���;q�yA�����¦���M�3,���=	Q�6�=[v4�p�[�&����/"?e�����9{:wh�mZ�Qбݕ��,Sf�dݻ�Om���S�5���}����3�)��u�
BP[����m�u׎R��td�[�f!{w\���@${��4��*����3�%]��W��n�9s��U��{�5��D���k�j8�d�ޖ�QNA-��/��I�S�"`���,'�߳���v���R��kV,a�TE3Xڨ�h�t�S�1i-����N!�)Ji��mC0V������Bb&��mbJ����j"*جEL�r�:ረ�mZSA֌MΚ���SAa��c%�(
Z����h�b�(�l���)"4i֊
t��r�h�mAIlDP�AUO3�*��h���t�")�t��ZZ�UTTUuh9:��A��1�U�T
�M~�@|>|~�F����YwKز�[��j�	���7
)��y�'h����=���<ˡ���/|�`){ǣ�\�N�ۘ�=�hz{ċ�����|���v⇘:����Ç]�R��jj﹏,=�����ҧ�Ͽ����y��C���}I�g��n	�'x�̝�:���7�`�0�j]��1O�����^�{�dN>��y}C���z��C�+FT�����dC� Bz��7�	�x�=A�g�'h�u���)�^vs�rO"UM���������kc {�N�<��;�d=��y��!C��۷B�AI�e�O|���G��78��`1�DE`�䥻�A�u'kuz��^;x�B���$�z��OhN��9�Ҿ�����oc!C����0�� �=��	꽰{ψ�汸�:�t�C���7��q �S�O1�u��CHz�������w��n4�Ý�������{��������|�׌Uܓ��0����'h{2`�!�=J#̽@����9(s�P�9Gl���o	���L9����yxS��}
�bw�X��v���;{[���v��7�xM_|8���>�!�ڼЦп��{3�3����t�]Q����y�ٛ}5Y�2�v+Z�'�
�i=�Y��#.{�ʖu����3�8d�����L���qp-<`ps�9���N5	�-��d��3KB��r�^X��5��ˍ���>�{\�>dY�v�2J��f�2�+yQ�,{Rr�=�7���Z*v��7��mņ����N5ٍis�-���z��,�p�Ԑ��:���Sri�OG�%hz��YŎ������6���j~�����S^3��}ӊ5U���;��a�Y�W+ɗ��U���C����_�l��W`�b�$���8�{���x���0U����>�Ӗ�s�י�uK��XI��73�Q���N�k�s�c#z�MF�6h��l����ո��~8������EUo��kls��b��nf�r/����'6�yQ�᪜�Ӥ�1��#kbv�պ�'�ơs��F��h.zG*�5���o-��0�������i#2��u Ŷ�4�9#��G��T.P����]�ii�jk���ㅜՐ�uϩ]٩]�;�G�E]x����.f����j�G��\�˕��C_Y���I�$�[[��lef@������V�+AKg�⺩K�V��������:�,��7{�3Y���2�(�h�!�یۭ����wS��9~��9�g�V�S��d�B���^H"ȄT��b�u����S=Zˋ����#g`��u�	׶�R�&\��yq�k�[F����{i��V����������k����b���|	�+�1=���f�b�ч=��yi�^��μHN��W���|DX�]{u��R2��Ґ���l�Tg^���S뾒�,K?C������l�`�K��S$ڥ��oQzT�K��ݛ�|���e�pϷN�Ѹ�HPc�Y��B�$7o��������)I���n:���q�ּ�mQziL�W�-��o	u7}]��΂V�ȢdF�,w��)s�[�����tS-��L��JH���W� Uդ���YPnI\G	�>��ϼ8��ïkW��2�c�����q���&��<�^��M��V�kGp$�G\��
�u^�����	!�S��5<�3�/3����=�c?&Ͻ2���Q�$��ęʌ"Q-e�kN�N�k>k�a>���vߚ�ZCm<�_G���q���.0��yf�od����VC����ٸ��j���F�;Gn����	QH2��C۔�qM�����.�]E�./���l>��Ɩp9�pRR��ٜ��So�E�9�-��i����p3�L��n)�8o�w2.�2���+]�5R�vUfۡDvbUM��{4�$�Io�0v�)�K��x��J��r�2�Z��g}�I�Q6:�Rű�0�+�|ґeZѶ�1�����)����]k��J���{��3�+$��oT1�Pe,�]���ǂ�{���`���uM�0�IWma�8y,��V�mf7�m� s�.f))�h�+��%м�*��4W�K좟sM\<;>�2:T��Ǭv�Y��u��%)��:��ս��¯��/�8e)	��WO��|t?�SoN٧�Y#M㇑���T���qu�A��
f��^1�:t1Ɵ�z�*t������gd�:[���e� 6,D��:v�F��cv�l��l���ME�2�Y\�x��Ҵn�	��,Gj��q��z��-�oz�I�۽<�yTN�����E6��������/׋���{�vZ��z#"g��3���|%JZt����g�����a?_oY�p�PP>qww�����ߔt�J����-�����͔h����Pְ���`�����L�1B��D�M qE��`�@��N�J�:��1b2to^���LC(�ݦ��6�����dר8`>J{��ۻ�eZ�)_���F�U�V����j�~Y��j�ݽ���z�l�����.�|�Hb������Fm�o�H`�A�lPiM�C�/��6���Hփ�+��63.ES��lf(�C+3��2wN�Z� 5�n���Ӵ�8r�I��6��I�k��ˬ[��n��K�s���u��+"i���4x!�:�����j�2Bɼ�}L�"�
���s0�u������z�Ab�^.Һ����R
锷"viF[M����0NMX�V�����k:��)�g��1LCT�hE!�����I�7�c���J��b�=]�$�
�ʼ<N�Q>�=%�ߊ�qs�G���S|����Kp��3�o��Tו��Һ�+X�6��T���u�xW&x�t��c���*�꫼�=���9w*i��q��@u�V�R�g��{����=��۟k_��x�K,��g��@�A�J�$uׁ���qnO��a�l\�z�oKyG���*�qE���{7�T���~Ǟ�ջ}Wߺ���"ڥA$X4��A@VkE�BY��Ķc�#5�as,n�����Y;�T�J��\�r������
�!�1���i��9������Ul�������w��q��R�V��pw5t�ڿE����M�l�m<��.K����O�=�[��s�3�P�2
%M䇹��Dǽ+d�B���\�|���e�\�C����P����ޏV�U����a���uk
@Y�����p� .�ڵ��h���3����y�-H�����ۥ�c�AYte�r��� y��]��Ļ퟽��ﻑ�8��PP��22���Q �˭9^RE�j�RQ����2�ș����_��p��^���-�%�ryN~ή6;��*ϫ+bWL���끄oGM��Xf֒�(��޸'��NE%E��vܷ^m�(-@'*e�xm'wJ��v	��a���)�g���,tc(��^ם��ps��])���]�7�
� L�
+},�Y���/X�*#t4;��$o+2�Y�x�M�ﾯ���s��y����0����(���AG�&��cD��/?	s��uk��^k�H������=�zM���O̙���}�C���ܵ�㖁s;"4�)�7��r*��u�*��"ct�n%J���}D���g]�jh��6��D\��M�oYaI�-�{����LT֞y��%�}H�VS����+r�Ze�Gz6�,gG@k��Yc�2_jz��H���,�8[�d?;4D�Gu額}'
�^C.��ЌK��H�m�q� ��2B�v�r���F-m8���y��������!w��q7Os8rNr��d��J�h�k�I�������{�y��ܶ.��k���&	�F��!�2�,���� }��)�A�ǉ*k{֞P�ĳ�td7�	n��d!ٺ��ƨ���Eu�ԉ,��k�ݖR���Θ��=��^�s˵흑���=?t%EA.SoV�t���:�^q˺?�着�;'y鳏�;����$S�Sǥ�=u�a�&o���9�%�F��ξ⩚�9�ol'�u�&'
e>��Y(>D;>�D���"$�����3rɦ6@ci��&��\��q�ݮ��ݤ�������a�f���Ph�����^���51YVa��ꜳN`�cm�o�᫘��2�M�ں;T a+���l��)�=�Y<u����	9
EՕ��L��Ӡ�Y�`�!V�'��ѹf����Զ���%����Y���>Ngy?l���r�U�MH��<(�9;���P�]��C���aA�7�������[w��VW�G�MT��M��t�*w����*��G=j	��b���f�=GE�0^%�Q��C��-F�k��f��@�G+La^	S"w5+�[y�p"0���R`G�ӟ���e�[]<M���Kv�
�s:�\��ܤ��=T9o��ۭ=���ز���{|z:*�}a�� ��h��u!9�D҇K]�Z�n&�UE7ړ[&��V�y�9�P�&��������2 ���kj{��~�W\zNM�d����6�hq�&Ѱ�T�B|#
z�/��{:q$��㷽xELi�A��U�7G���d���2��(��%n�Z7Z�A�-	ds3��$
�V�Y �!L�"s ���f�v�X��'I���z5Y���w
�p��7j��W[F#c\�[�S(	'QFdx�ϋ̧����]�<NFr T��}��T4�\1vg��2����L��,%ɽ�:VK]�È7��UvF��W�GT
�ت���\��&�M4��$d�MFu��s��t����5`��L0g%���H�Rd�H���7U�,:78]���|�*�w���;O���NՎ����nQ�p�E�c���wv�ɕ�5����g#]K��VK:����9و��X{�Ӥ��ҙ�>����/htu���ڎ>�����Z�W��-�E��|v��y�9�%�Zy��I��2V*J�
bʹ��xrT�
��S[6Qiޠ��^��v��hgM�tv�'y��s��4���+�δ��6gKj�K�6�fN�,nkB7��B�S��Q�p�0����']f�X���G�N�a��������]�[1�4
S���d
�\/�>�{���s�;��_Y���3�nT��s��䝱�]��Բ��m�J��]M�Gf,��	��x�TW���`�X�]B�S����Ro+����lFx
e+������;�]����@d�qi�r�����Ti�����P)��E�[�(a1��'Ƹ.�����n���Bѝl�!���^�-���@��b8��\�<0��:��hu|{����t��'����[��|�5crn-�V!�qPa�)V���9y�ʗ�ii6��(��[	J�-O��f�������W��l�')\��(墭�i�a[��"�F����q^����:��J<�f��8x勖��
�\����:���-(c�Gz�LGbC��мTu��3%�w�Z,>�/'|��TF�qnAS�Uuw�fl�˧՗�Z⢀0��� ��U�(��q�اĮR��,@�[5L`�t9}�Nj��ea7Hc�m��w2�+q�͝2�I-158y��G��U�Єn�X*;��67��5�4I�����贞���yS!�;����9`E�S���qi^`s�[�����;�V�}YV���J_!�2�.�Gq�9#�����廣8AV�v��;��h�[�)�-��Vc����}Y��9.�w֓!�w�9���>��Qv$MdFىZ�:�ΧSP�V��S�3+�v`�������(�!hw���b˸p񸍀$�&1���/%��\���a(`��m��\���͒��`ސ�Y�-ᗄ��P��l�1T4�p��1�A���q�W��o�ޫ��GӡK�]I���7������}9w~��k�z�����H�,�m���|�_��_/��TE�V�9��X��a��qUPh4Nɠ(��-$M,DEU&1����A,EA�#s:j��$���֪����j�����������m�Q$TU]Ff �G
�DE4�T�I1IED�L�IpƠ� ��("kK���QIS2AA������f6q%U40SDRT�[)�Ә��"�q�s���&9j��.���H��"���:�jb�i�I)��h����M4�Q1Uh�AQT��U15Ai�M]y|�|	���L�i���G�]�ܩ�XRE�؍9��Y�7l �Q��_V�P��e��Hx8o�p#o&�O��P��ی�f���G�>�V,�KL�͖'E��sls��z���J��.��lNfi�|�{}�;Fo������2���(��<�դ}$���{���b��,��7$ϯ�F���5�{����N�M������ nв��S���J|��O�#66�ó�?u�X��*瀃1:u��q'lDT ��қΧc��W��o�>���C>fߔ��Y�q��'*���1���:tT&�])y�%'^���%��6YQ��E�U��v<ic�F��FM���YTR�����` ��Y��͝5,��Z6`k����l��e)��Bѫzb#5��զ��5��l����a;���՗7!'�zGp�c�Cs�2�i�\|�g�P	�"��i�I��õC�S>J2)���b#he��+�������"Q����"�/���fw'ڃ�JN�]e]�c�%Rk<�J�Q���[���e�S���T6�=���X'������� ��ÿv|i�L����Oʱ̴��z��=i�5*W�x��g��zѷ�nSMl����G:u��^��m�����ZsZK���/>ͬv�Ad�S8l���7����Զ����3[��xL�ӓf�A��v�N=���FF�Z��e���I0Jz����:XP*�Մw1�=��n���U^�n�b�֯���#���x�[�j�������g�Q�k��M�M��
MD�3NQ�c��>��ʃ+wNN��p��}����xN���=u?>�M�2o*;UF�k:�N�T�ֵ�Ljefs��O�[�
�3q�A[��ۗ�������¸�zie�u�[-/�-�T�`�`��c*H�O��Ջ;�҃����[�!�9]�eK���:�1��:��&,�)@��그�S�5!����e�wZe0l�]\;G|p�a����=�;&uM��ܾ����-s&��tv�L�}u�������2�/	A�8F���~�P��T��-�o6 x���0��X�|�kI��.��և�O�vw]����ր���)�Mfnc��	�=���"7d9�L�֊>Ɠ=�zf~��
�	�p��<����O,��t�|��e76K��F�c�q�� i�w�U�c5o�O:o��F�d�X5�Cľˬ(�Ƃ�rqD�el��P�D���_˫j~�»I���͞�y�{df�R�l���Z�B���§�9`-S1�jRcd�,L�� �4j��U�,�K�o�ܧv�H��̻��+���D�q�ݗ���5�p��@�q3z.��ZY3�4���Z�=��(R�4�dWqu��y��N���K�A���ɘ�`κ疦�V�RS�d�,�>�|��I��b.��U0`��ӽz�X�S�ܦ��n��`S���B��c�-Ǔz��J��rgh�Y
�ndN�/�h���19���x�-�-�����+��YT����|�O<�q�/��5��������D���\�p#4m�m�������&vo��c�qt�/vp��YB*��Wt���O�d�D�H������l�z� ^����\���5����j�F�L_:=WX�u��IӞ2�$��8�ew.Ϥ���|��u�G�OY���|�2��5J���W�f�ͪc�r�SmL����TdӅ�����1�=��ҪCt� �w�~�����ϚtH}�OZ�����&�3d5;2�Li��%w�UjkjYc1���ˡ��ú���O(m�GWf�m�l�"�z�ȓaS(=��(�a��|�f��հ<5y���b@oB��� �B�ݟ��܃�X��;�+����n�6��<�F�q9Q
em<��
�rgo�[�$�:��h�J��L�C�TxvZ�o�(R�u��qA�U��٤7�
1��]_�}� ���:B���U1����{�p��f�\�Ŭe�ϫ�	ձ52��9���&�R��QS��w�t�m�Ӛ�RLN�#Jl�F����E�⡖⼒P�薥��!��5w��FӚ��]}K�C��yU������x�$����w�3���f��n�֧���4L��(��]�r�՝V;r:y���^2�Sِ��,�Cao�=�>e��+Pܕ'	���6���6#3aѹt0���F?t;����fÑ��(oe�����I0q�`�[��ڝss�U5�k�Ig�����E��dUB}U��P�ӱxqKcQL���1ϲQy�Ț��L	�>�����0�f�!��h�	j�sZ$�U��. �.�t�4�a�q���0[5���T>(Ј4;� ��]�P������P�:��x���q1Rۨ�e�	��`8ocn0�v��ɡ��3�7D�4�C�'*afv�"�z�j�!�����X�a߶;�k��f�������� U���b�6xȔ�\�ڷ6����ǯ⍆�*�B7&�/�,�F0	�s���sZ�֞v�<�bV�Ѷ�>\�V����w�����!��]�����ٹ=]�y��[���l��)R�敹�8�&׺����j^�0ޢ��P���̻��z��
x��(K�>U�����I��e^h��O���	�]4C�v5�R��$�Ow6�A؊�\�8�&��B�T��e�F������]#�M���Ꞷ���@�s�t��8n���I[*7��z*����y\8��֬.��"LY�N�iЧ�dǝ�y�I9��e������Q������{L�	M[^S���m��Fݳ!wq�ȣO��q7�y-3J�ԘN���k�7a�q#o{�O���~ڛ��[��s�Y�U�PCzH<8���[��Z����@�n�s��P@q�-�'ZQ�5���k	m���B��h?�� UMQ;�[��ꁂ��U2���{��\^�����Z�5l]�_���ُ_�G�|�v�w�,�oˋ���z���'MB=��kpx��'z`�����hm�k�gP)����%麬�z]�FWa��S�7���qݒ��~��9I�i��������Ș�ڟo���=<y����A�U1���ij�A��[r
�7nKD<�t( �!�Z@/���"��4�֫��p�u;��hrX�xN?�p<�/�y&X�^�(�<�%	
"z��q��8�]��I��'���^���c�����^�����~���g��n�⅊0��2n�5�f�D^���M(^���OAP��z5Y�U#Jm�N�e����?\�p��]��A�qi��D�Q�. ��cF����6$�nS=�1�Z���8SZ�$љK�6�#N��W%����˰������v:v4#\2�WVw*�L[��t`&N]n�����x��&IBGdW�v��n��os��r�n��06�����t9<M�A�0"�XMbT�6�g:^�h�`�5蝪��d�sִ��n��58k�;�J�y�(���@�lNm �$={�לO�w�Ԥ-E�~�/ս�6����@�UD�I�����d��\�^��Um*(D�	Y�NuV�G&v�/�=���[�Z�u��q�n!�c5�~H�I����Ƣ����Z)(Te�Ғ�o
�N �E�DL��7�1�q��6/Y#�"�v�ُr�з�FP)ט�z�7i�5�'sNdO1ݦ��eDX5�3j��ԧ��˱���9w�kjOs�-ח�k�Se	޸����6���ɔ;� �+�n���:��"��Oި���GT,[�镛D�
�T([�X�ۡu�A���K $��Z�c�����|MkF�Ղ��XY�[�d���+ka���ƕ�Mo��b�SZ"fo� �����;����:����2���[8�e����Lcf��jԔ�Q�[��ֈ��{�17�
���ͦ�b��O����%���ζ8�kCs�=�GO��r��;���ܣ>��jp�vT�k1�e�ʠ�`�aS# �M6�Q�J�Rq�nْH��w�_W��m�M���t �I����5H|��emz�2���(���x��hj�҆����kX���L�k;������w�F��B���V^h�}׈/�׼���>R��L_�ǣGj�v��2��٨c��>3<Y�1���D�<�U�t��^�I���z�u����&BNV�sY��O�<��W��Ö�,=-��L���F����}�k�͎D���r#Lk7¶T>\>�Q���O*m�{��W��G}�^��r��fRux�+K3�lZ�fi��z^Δz�v�H��\�U��w���Rp�(~B�Qef;�%����4w3"�b�����K��I6�rE9���Ec�l��+��"N�i6ӳ)ӛ��7TZ�*D	%�r�$Q|W�s&�-��#g�2�*'w_	U[��Д�;��"��=�9Sة�G�}:C��l���&Z��\���|��HJ��ۓ�������Z��"��:�"T.ט<��6��<4C-���W�����#�!n��kVt��-��\�y>��ͱ���*�t~�v�}�y�q�m��Խ�y{Q��7��]��wsѵFcKt9$�Z�����>Jz�06۝�М���m��^=���敘��M�y�J�՗G/<Jx�̈́���[�x�4@clj��I�~�͉��Ci��CLgJ�G��P/�\�0h�o63x<�9�>>Ȫ��\��.���ͮ��8��|��� V�c��	�����I'ot���Nv�j�L�����A>70ĥ�!�w�� \�ܚ�bG�G�n�kQ÷%s�3�+4�s���u�K�8%��k�^����Ջ1�ǐ�j����%��gQ*#�E�-.����Gh���"������˹Q��c	�f�[Vv��0d����5��ˢ�3jwww%V$;O�]9��͘ʕե怾�S[��&c�+�>�V.a����Q�/�OjP���䮩���i����-j^����d��\w�{X
J������e�`
�4�jdE4�x)d���'��2���A�S])�ز>�:��0���d	��͡���\�z�Q��󱍝<�C�r��>mb�oGf�nD�$7�O:��CR��@鹈�ae���v�������F���}ZhMn�;Gm�/L�ud�-�Ӈ "b�Zk�S��֍:P�5�YW�2Ѿ��|sV����5&��m2���|	֍��{:�.���za��{V����V~�ה����ݾ�n��ᷜ��/;�e�X�ܹ�g��3:����\���m���R���wmX<xZ���`�em���ԭ;�=9mp�{J���aYn[9���]M7q�N�M҄��z�Gf��;{�)"ɣui
(�0��Ωb��R�j-���=2�=%�ӽ��K��X�G�/��/�D��4y*�U%�e1�U�vQ�sOR*�� %��P\�[�J���)d*W�Ks�Q�[��]"��=H]�|��[�KHJ��w�f2(>�kpse#;�3�wp�|���3S�)&�ג�c^���V\�2���N�_�JmN��[C�ǬǗ���0�-`ټ�X\[��	�g�ѣ��N;�>�ġ��r�L�XT���.U����-\��[0;oW$�n84�3���*���%������v���Nq�b2檷�� ��s���߾1h_]�t6KX�.����uF�$�h��Jtt�7�QUD�KRm��*�&h����lMELm���U7[1�TTDDMDGQ�
�h��*���ULQDDӶ�*h(��&�����U%TT�1��i#F��Z"#c�T�uTQDAQ��u�KSG]c�T�E1D�2TA��TI�EP�QQQ7$�\�4�MUSUM���cULPUS�3!�H��b"&"����)���"�j�"����1?C+fK���1gY�/7x��ij�%�Ǫe�݂�W��1t7~�dF����x{���T����}�l~���$�{��T6�ɠ�9W�>\�W=�A}����e،��%� �B7RjB4��Sk�>�O��na�y�9>�}<���e����b6PFz�1���8�g�Ճ��[�e���l�N^`�����n�V�>��2�i1ph�Z3bt��*i�O��N�髍�b�i/�xNj��}=\7T�Tv��&��km+��l��n���MIթ��{.�n�ʧ��s�u�Ec�����<��X[��+@�:F�dV�TVjQ��-�Y険z��ƺw���LEc�"�f�U�ʓPX$�e�y۸�eIv�׺��;e�Ƭp����O�e%~�@�i�̔����p�c6�����u����Լt��uFI�a��ܦG3�@�
V��x���)�qy��m��s���U#P���wi[�s�V����Zc�C�/�����vt\�D���=� �ݼ1@�=��~�f(h����0���t�t�}[EI��t.,��� }����k� ��ɖ��E��ѯE%s�'|\䶂g�߹�}��35�T���"������w���Od4A��]1j"�6���������1���3���!�hRwUp����e�����ܽM�c�}���t�ۆ �[�2+y�Hގ�U��J$S	J���v�E>sI�%98�UC(V�g1n�E��+�b��P��N(��gpQ�Y3�E�{t��z�T���聙|���SI���P�F�ګ���6���N�*�G�%M�U��9�-�"o;IZ��Ճp>Q^�����dղ�*���:崩�`�G���8�9E�/|7��qM��_��}�+��1+�6��yﷰg+�?Z=&���9Dh��N�p�L*9�!U��pU���d�C��h���&�v��}��_k��`�K��]�r�;�K8k	S������#�ƛ7��:�d:*��������8������iy��W���61Q$��A�/����n~P�R��Vvn|��Ӛ�-xi5ݼw��C�Y����r����7�b�<�ϛzM_8����N鉂�y�)c��7tϭ�U�=O�0���`�|j�t�@�:�g�¯��^�D*z�(��y��g�.C:8�*�C��7	63=�M-�5�[��`���R����ٕ�m*��)�c��H�[a������[.e���5�U��,�lSV��y�屚^on<zs����<S(�FYws��2w�`�0�&zX����kx]�����A�Oo �|�B,�J��Tr����c_k����TJ��Pގ�i�6��5�u��H���e��Ami>���=��j�=���,��#�/���)Ѹ�Z�����$������'>Qt�D�°�7_�U��}Y;zzw�cq6�m���q��²�3E���Eaݶ�:|�_�r�N7���XoJ<p//86�jtX6�u�~���Y��b�tO�Ly[c6��"�7L�;�.V�g��Q�&��O���H�9,���ܝ릌<-ݛZ�������e��.�YG��[�ႮueǍ�[r�����2&�ȍʃRc�Xy�w"x��h}=k��ﮇm��',�9@��D�hæ�@�h[=��۔�G���T	Ӫ(\d�k*��RF�p���\=��$�>n��/��t�eIx�%]׼Q����i���������;LXZ�)K.hs���w6�
�=���aLt@���zN�n�ɀEdy�`2��Ff%�5�$:���*��ڿ��Z�J���]mN�+��9����#�n��:�ho��%��%Q���l��C�5�_T=�j*�a*�Rp�����=Dg�	Y��\&2�5엂�K]�_�.LΏ��;v7�c��Ɍ����q���hCܴ���.�����<<=�ŴJT�2��{b�c�m����\ǅ:���a�V�c��Ҽ��ߥ6]<��&[�}�:�lL�Z��;�8�5�7q�D�����{�oG�{��W.��GNn�w�Zݵ�\*��K�l��8&�+���z:n$m�4��V�{%
� ����⃽Kh>��"��=E?,ϼ.����
*Q�$i��^���5F�x�;Y���x�`�۬)(h4���1�Sg��f*Ŷ�|��mҫ��И=u-bNk��p���b�^�Q/ڭ�nz�0����I�93Tm��
��7�5h��L�ͽ���X�E[*�.1�+��]Io�Y=�uu��+�cr�^�[��0e�LL��=��2z���u�ڔ����{^1��-F���1������d~�	��M��b���Z�WkЩ�iHp�����<v�D��<��%�}_W�:��B��'>�EkU��m�pV���wT�G��Ig�˟'&�1!p��iBŜ��or�,1:z˷B�R<lG���:L��"�&֊��IR�G��x�_��c��4~���;�e�5uA���5oJS`:MZ��&�H8;w��7GN
�����cǶ���=�WA�Ɖ&F'����g�qa��o7��*4�2P��Ն�<�]�xL��Ǩ�7�4m0�{�������j��8�y�G:�wU�'=���O4���N޺��l+D��;I�l�n�s �B�P}p���L-�[�x�<���h�":{r[L!�kK��90�Q�&�O�(���\C秜c��{<>�G<��%R�kF�;#�v_���0�ǌs����؅���,8d.̖�ˮ��A��۫���$�����h�<���B=+K�ΐ��X�V�"<d�+c��~{:����%�ɕb\�N�	�e���jAG%u��e����U�����j�����6<WX����T�1;���EX������I$�(���񆭷5لgSB�>O`�� ��xM��1���S��[�M�}��+0k��VQX��E�	э��I����.Yu��ݵf�9�_��������%�Q��|r����J�re�:&��7�dg��{.35�T�e�;�����B�|6�P���p'UQ�n񑚮G:E[r�X��NwF����u�&��{��o.�}3��"��r����ĻT��������؀�(��tL[�2I'}�=�_v�ݜ�N�㛽K �]A񷶄S�[<ْ7��i$d5zE@i��V�q˺�T-�c�@1(����^���U9�ګ2��%�:-.~�JC�>�G%S���~��(���-���{5��W4���Q/B��-s�!�H^x_,vM+�V��m{$!f�I��b�z��P�)a_;�s��}�U}BVU��Eÿ? ��t�9���M+��]��+�Qz34�m�;��1��Ȳ%��M�"�;���ܣ�uP�uJ�D͝�Z�R-ȏ[�L�c,�w��.k(�e/��1��2�u;5��u�f9�y��NHx拍鎃{��3�,<�
�cX]�j��4Z���>A����vBp��[���5(����{�W���0��.��z[��Kµ�<e!}�Ȣ�ο�I�wsU�{L�Zi��Nd�\=j���枌0[:_3Ul��S`1�{-�{��٫�c����I��	͕D��1̤'�R�+.�96#n���zZ��7wv�q+��b=B�f���
��r�uŚ�����s02aD�8��*KV�)���w@%1уrd�6; ��'�7���gq,;w0����7t_s����R�:L �cx��c���A��Z뻛1���g��A����ed���=��Y�������O��m��9jb��}Z�T�׊�Կ)�S{1[����
�S��q�y���?!O�i�����Kn��z���'.-o�i�	���sT{���IB=$pէ����ȼX�.䬉��"�Ԗ������*���EMk�˒ic��S��^S�^�C-�3������W�o����5{�[^�=�@ǟ�sF˾ �s���J|ӱ}û��b���J��{�|�7���Ԉ��Tc��y�b�NQٹ�UM��E���m���f*���	&�iS�5�FT����,Ǜ�Qurt�!dT#űKXܡ�7�j����uf��=��\����I潌�ǧ���
_�T dԭ���/D�s׿i��^��\�Wv�R�k�nC����'��u�j; 9���J�5(�z~��GX�T�5KY���5N�Rjv*�m*�͌����|�OzJ�#nk�Uؑ=W�5�[[;�F�Q-��!�����Ҩ�O/�Z��GXn��q����=� ���ө�7���AD���)�9�Xr޷����dF�f�Z�|y�U�7{zsU���f��.-^��|��9�⥗S�Vk��zח�X�t����Q���6�dhʱ�{h�˸ug�֑,�z�����-+Ւ�4T��=g 
|��*�D���iʦ���B��u��ͯW��Q�Taj������s�D�{]�Uf�N=�7�)�~RZ��1��O���q�I�S���ۊ�2�����gj���nf�Y����]h�դ]E�4E���^����*�C�X���۪�0�g�.�c$m�~�/��(n��ON��P���jK8�t�hU`���3���x�-��O8�#���Z��J��mUe�F��Y�iP��ʣ�B��d�[;����uD!���?��ݼea�ܼ���m!��(�A+H��
8���{�y�$�Cm�6�3�(�a�E��2��� �\��^ ���vv��1�c;���Z�+`��ͧ��U�B_Kc�ͺ6����x��K���t�������Թ�д�+i�l��c���u�ڧOW1�K/�R�_N�Su��U�Cz�����Z�ռ�.�5r�gegdH�Y�k ��u�(�Ŷ^[����T��[vFv��ëSݻ3&+�.��O��tx��K��w�ΥY�����^�(d,��O�[��7����O]��5G�N01bR��*�kB�wN�Y���j�e�z�a�����k��"���¢ʽV����&�H
t��%���}W�\z�4S���e��C�-��]ЍSu��"�v����4��8���3U Ȟ
����9q�SprF��{��{䐩�R��n���خu��M�K�6��*�[�OEJܢy_h�he�P��Cu��4����}i_[ F���b�9Qg;/u˶�=���qY�f���/9p����Q0h�.�5I��^W~ �DJ"�*�4��	(��Py,�I6�F�Ą9�m+�V{�M�D*x��a�v]vY_p��GRQ 5�W\�xZ{4ݪo�ꕐE�;����փ�0r�i�YR1��P�!�2���i=��N�����`Ay.k0��� �35b4�`����R�l�&Eb=���1����
�ni��CO��Y	ʕF�8�FHxCS�KH/�~�����U(!C;�1Г;L<�����2�9���x"V�^�*���	�ۦ����d1�GW�@��@8�ؠ݄'+���)�9dǑ%Ѩ�Ҧ��-���D�/ZB���q�ˤ�uڃ�]��m���.HD�h�[�&JT�7�i�o!��y/p]���4P�@���L�v1�7�]:����dJb�Z���0�v :
�ח~9\�%��"��fRG^�$���`�+mҥ!d�r�v�>��5�;$��!U�%�Tu7�{��J�h�S����p�_�a3�PSebv�����{���>N5&S³��}`#�8��!tYSnJ�	drEZ������Q�\��.W���u�¥q�p�v�Dmj�w9wt����&YL�������j��S���(��������`�SD��AMUQr14�CT�1MDS�E4��11���PMY�)�*��5ELsj��("4:*������@QIJQLG!��\�EBh�UCIZ�h��m�m�!��-��JG:��R��j�(�Z�a��EPE�G!8m��(���(ZJhb)4�)(����������*��hZ_~/�v�]����vۮum��:�fAt���=�w�NH�2���Z�s�˽�����XŐs��y0"���=� `b�i�v(�.~	ߟgt.���9��v�wS;&�o�̺j����C�`�N;q�W��˪CV?^L��z��'Nd���/]�Py��:�t���SAmX&���c7XJbl�)�f3sj��T����F��S/��lۨC͊���9������[AKY�`N���Ms�6:{��m��:������㶨ה\VVȧ��W*��R&�a2�r����g,gŘ�Ws�q\*��w�B�x��/N���ǿ�׆�5;�=�;�	ʯ+T����a�8#,e�e�^��vxk�oe0X��r6�6��U^�������!l�u{G����W5�&�^|+_�Z�����(���uC��r���h�	�|�`W�k8��
�����#sP,��PU��X��ɸ[K���y��&�&����q�=�rayg��� ^b�ef�ɕ�"ƪW&4d�wxXԭ<�LC|��ur�g����3�*C�@m��D|r�꺥�]�
fU���'��_�̔r����ۜ�Vy�h�}��z���o�̝�3{����vYj��r�$c�5k�%{)��^��1q�Z�~B���p�t�蕕�21�d��OE���d6nvW ����Η�AKP�Zq���v�t�Ǩ�1+������bs�2�I��Em9hOW�ۯ]�i�ή����{�Uf�P��lF�|S�J���S���`8d�T4���m�Y~�]7�V4�K�%��$�õ�ks��v<��+�ĵ"�ɪ�`��N����bM�������|�f4�yN@զ�l�Uv�|~�����2��rp�����]��{��ɑ4NV�Ʒ�r�dٻyۛ���>��'�B�C2s9����x������{����'a@e�\:������wD��]��`z�,,5�_USY��a>����ּ��g�:b�t�H�95���ڞ6q��6�b5�2�˿�9_O�z?�M���*.+I�ó"E�U�nv�L�inW�؉�דJf@��[�'}�ׯ:fF�uV��L{�t�J!3��OU��(�J]9R����b�pL���)�)'ȕ��3vx	k9)5o�^�k�²�#�AКO�mS�э�4߲�"S��/ V�����&�⋎c�b-�,�r7�6j�߉��˾�q�z8ǭ+���B��f�ڻL�gލ�Y+��60��m'�!b�B�FYwf>��tC=�s�Q�M1�AE<����3A��/�T<���6fEPylk[d�ņ{�G7Y)����8����˯����D֯��������\�u���j�s��i����љsl7���c�>=�eȜ�B�Mn�-��Fd�rA$<z_<3N��[1閶6����c��&>�l��b� �͏����4���ƽ`9�Z>��ێ���n�j�O=q�6F4���\ݝ᳋.��SQ��A���.I�G�C|�}���~�{���m[-q���؟4>��
^2`i�$c����]3��۔c:����nM����/�蝻W�E�+m��%JzFYG����z����+u'ٚ�8U�T��� ��C����<��[
Dn��{2��+u��f��[�3��R)�K��}q���dҭ����g�.�d�ܞw����J�kv��b �P%i�7�q�22!��K`���cc]G\Y�Q��'Tx��(�ڢ��Ln��nMw���X������OA��-:�1T�O��&r�ؔ�u$m�t)d	�5^Tg�`�iWz{����I�40�'�Xe�߮>v�X�;B&4w6�L�4$j��p�!�"��*j5���uf*�4EX���4c�쫦�{��n9N(�}3�˙ƕ]�bn���:�W����v_E��������G����T�u�Z����z�-��Z~�U%���*��
�E��'c#Yd�RG�f���p���YGK�@]l6�B�%C*M�j�nl~���T�T��{\65�9�A�c�5�f3P�&JYD�^�r����r��<a�
�G4�-@	A�s�3M�a����oA��g�B��I�N�'+-ް��l)��j�ʓѩ<���W`Ʃ�eP�)L�ℶRz��Zl�+|Ǆ�q���\��c��y�w3񗪈K���D�ɻ[o�¶C�|�:���9"�cN�Pz�u&~���:��vfN�f��H��5jIvͲd�j���F�\���cQ�zbS�۞����x�2n�'��N1���q��z�YJ��]���P�3aȇ���v$���닮�ڂd�~#1����<�m�&9�&���|�Ե3Q�R�;�,�sŻ%���bA8$F���p����{�Uv�ܻ8I6,٧2Lצm�L�1�OFL�����$s����������Ue�z��2�2y3;`�Pl�m��lS.��'p�	&�⍷4Nq���l�V����HJ�чf�T���f��OU�ݸT�
��r�&n����/E)�c"��h�ܑW��4k04F���^��Ҧ�|�^�g~תw���u�\_uU�~aw����t~�5lzc�'�>��Z�U�U�;!lXb���!��fji^�q0֚��t�\�e��am2ծ:�j���D@�uuW�������[�2�>rCJC�A��y�e�v��g��٬�����$JAH��=�̇�d����82�[I���W	e�X;�CZ\�Z퇿_��޵�6A����MŮSnlk�t�7]:�M�#yb���}PFM�qE0��=��/'����S�r�wQ%A� ���VE5�7xKS�C�4`o��Lep�Y���Q�f��͇�?< �T�������k���OEH�1Ztr�z8׹rҋ�P`�����f!���m��U��g(���.x8n�t�P�Wh#ntH��P�``<q�Z�<��xY�y�M�;�X�ڤ��#��YU1��0�xF_n�ħ��Ca����4�rk3m�Z^ӥ���u�WX{�'��[[x�Vk�@�X�F�1�K�*��ug� �j�ⶱ��n(�ՙ�"����2�Z'��ОE�Ec�8H�����BWך���*�&�B5���r�Q�2'y�N_Hy��lx����Ϋ��3{ԇ��a�n�Bo�1�׽>~�{�_!�r��s-�-�IE�M@��2iUxYb�y�=N�idvX�����hu�F��i�z�e�Sʌ�)��Ʀ5�Z������˧�*w�?T�5�m6��I^}����1����9m�0�θ5s�݋
o1��|�GP�����ˑ�����p�s7J�ǽ��!�X�Py�m'Ng�O�S ���)�1���u��K��܏<3��ɐ�&K]l1�.E��:�j��*��p�v�f#�[��y�cK���P�	�����hokZ��1[�à�l9���h�U�޹�=3w>�3�j�� �r���*7�vf�ҭMV����_|h|~�i_{����&�M�.󏵋ej��ަr�!9�b�d5�[����*�wg�D�VhSv��^�hN�n�4�� �*�3�[����?�ڪ)kf�[ u��b/E�3F�EQ'�6v�BZh�V=i*�7
�^5U7�r�z�S:%U{Y��Grܴ(�-w�;�qw[�Ǹ8Ǐ����(�o�����;�H�*��b,;2J���aP�;�<bt��fo|��t�|�rr��np�V��`W
�c�C��׭�:�h�M�L���zV��9*��2���u
��!��9>���ed޵Y��� _Q%�Y��i�}�W=53�>�Z[��8���W��]����+3:�l��뽽�!�LS��ĉ+#5m�N���ɯɿ�ʑ�kU)�S�m���[��H����w��mP�n��G-�aا�8����1Y&���u�>ۮF1�K�Ẕ�xNVi'Cs��h�o)�ސjmewAL\��[r���1n���v��'om�.0o���H��ao�!�$5�N�����튉m{�Ob���ye�gX�,��b�v�q����]tә�B���3b�V� ��X�ѫ{b%exb�g|���{ٗL�7xU62ᶡ����C��?M٨벸�w2��;fR�ʌ���ٻ2��;'z�S(NnC�#8%K��1���Um%��띖*�>٫��5 q��Q�eG�f�u����YB;���Wp�\��������8�6q��č�\omn�v�N

[�Nuom*gM=J�޶���q7U��?x-ԭQH�އ���٪��3Q�lr�y؅u�H�ύl5�[ʻJ��T���bkۀ~�u�v�'�xOM�}��F�ݺaV)��d�W�x�=�Q��N��Ւ�o0-��L��j3Eq:q+�Ջ�!����Qie��;�i�l����j�#V���
.ؙxv�m�H=p6�mPƟ?V�v�wϱwC^wY��҄���~+X�KnΜk����Z�F1�bƃN[�6�60>/F!��l
�S읁��t�Q��D��ssE��<v1,�5���E�Ps\�+y�S��!�C�Ǳ]m�܈�S39w�(htr�%\�1���]������W�'�����Ū�w��T��hǥ�g�[r�G��ڊqfZ�� �4l�;���F���X�k�}��|��i1�y���M�k�&�^��V��w����.3tY�
&)�.�����{�����t��Ox��C�z��ec��C�.�.�	M䯺���3;M �>Ә1�jk�&gJ�>ciT!�܀�{`;t�]nup� 3X<����R�"�5Շ:��������.ż<��ٻ��[�b���*��c���_lAF�K����ob][H�)�B�{�3$�3:���QhQ��w֧n�<�7��k92�\��8���__+@��]v.��(���4��3u.ĺOv��X�x�na}i�4�4��趁��Eշ�4VM���T��K'�n����b �A�r9��V3��p�H��ze�M�;���.zc|z�uӛ��G���x8�1�#�šɍ�z��e�70K�z�q��%��4wq#��	��7MQ���/x}�r��Z|������v�z1��֖����Ή8��j�4+3�L��r�.3�Ԕ2��=�$�+�A�֥hb�q�N��V���^������:��޲�K
��s3F5�b��%v�\�L��uI�ZwT��W
��|��,e��hR̙�Ѹpe�+��g������w��+ePT\�W]t#@����N��ai�K[6�Wy��9aJ�Ֆ��^TKT��=iX�sf�.�p1��M���1u�U��[6���_]�º��NM8�0LX��|+�-`Ң5K��y��gbnᙉ:��j�=GW�/>l=WPf}�h��Q���H�X�ֻp�	7GJ�Y�N��N�q=�;�!)�\;�$F�,΢6���rico��4�caE�J`�j��2�T�c2����R�a�f�,����YqIa���i�u֔RW��M�'U��吔w�t;\W��8��2�.�с\�`;�B�j�$-gu�f+��5u��Z2 �� ��%̰JL�VE;�t�R;,
t�����3��GىՀ[S����Rv�*=}t��&-<6��s�wyg�&�Z2x���נ�]��u]�~�Z�t=��PE�i/XME i�i�S�RR�Ji4iĥP�P�!�[���j")j*Z�������B��)6�T�@Q��p��&�V�H�(���h��u��
(h
i(�Z((��]34�SM�hӣ��6��M4�	E%!G ��LCA�Z�KIRi!MQ�N�5@P��-	��J���R�6iM@8��AKO$��%+A\��N�,�����Ϲ7BK^lNYau�k2�L�xz�u�s����3����T�V�q���.��������v��d�@�ޭ"�"$��J�Z���������h�O�q"0�D� ��Gt^hZ�:��C�C��'E렣-n��&��sm����+�1��,a!�_���D���"b���d&����v�z*����^<�ڭqwYYqM1A�'JJ��ŠS�l��[9=�Q���u�'�ձ4:��������.օ`����p+�}�����F]����o�]�D���Z��t�HA��n3��9s��pY���)�Γ�U�2eP�k����T�F�@�U�����)�:��Zt��
�^W��ܙ�Qt�:�Q-"2V
~r��y����r��R��7!�+G])gH%\�}ޗ7�]
��o�}�:��r�&���Ջ�T7=-�n��o�&�*0��m5�ܮ�ƴ�� ��Y{���Ӽ�G��n� �vr�njx���V��T{S>��͹��g��s�X�,��e�_5�aG��G�eo��XMs�幽^tA���J�ǝ�*�wUP��g�!6�!�^6�@�rHU8DtT�S"6gm�n]�P�*��],�
�;)��g;y����LV��S��Z�4�E�]l�;aq��v��JJ�T��r�_b��/�3;TPlcb} ݓ��C�gm�+~P��V+����Ja��Cu2�������t٬���,�[�i�/Q�CF�|Є�I�n;�VN���&4�
�l�p�",�*��&����V��D����v6���E[F>��;8�0)�'%=�!ζpW���ΘL4 �~���Ԁ�qWR��6G6�c�XkHNk�<� h�Q��q<kk>�uc�S�V�+Gxi�V2}x���.��O�ч�����M�k3�����/�<U7�J�v͗ڀ�!�Ǿɭ����{��"￾,���$�c�s�7�6g0W	4�z�֌��N
T6�]�=�X�%5ڻ���#��[��$B멵zb�^��7��Z�NP��͝��>)@���-��P��p3u<?�5��ɴP^����s��H��>]n�jZ*#��D��b}�\
��u^���kJn*�Z�6�UJ�ԝ:զ�$ړ�t�0f);�>��i�>�ƃ������챉�܏�	]#���<?c�[<��>��W˺�*X�)�˗�o~�ho�(9ʧ����J��g����5>�'�좛�6}ܹd�c�s��Ѥ�G���_ȿ���h��������r�Ӻ���wOyW�ܨA� 텶�u9�9}p�8DԄ�E�V.-���`�cNI�kђ�ٗ�
�[?2�7L�=��W����q�A�C�^�m��y��1�h��{Q����+]�r�Ϊ�!���h��Qs#�z�mf��]pk��f-m��EZ�gӲ-X�(E�ƪɚ�:
�(���Ø�ź21�C��PR�V�z��χ�q�����gV<��nu[��v��L`${])d"t���;z�ZH*���MZ��K���:a�z���Qܧ�ٗ���9��+��Uf�Uq`�j���$X�p)l��:�3D��[���zA=l��ΝGٝ[��p�jUV�Y��0�:�J�oZ�hD���U^���������\ X%�g�Wm	޸Z��/U�·+��T�n��},��]PSX�檵��cD����A�?jN�vv	e�����o�ە\��ga�݈t�AY}�����{j�L���/�/�׈/�ȡ'�2� *;vOّ�Γ;���i
ȸPN��z/hJ����V�� �m�QS�.Z�BOʆ�z߈li۷��d�ne�aK]K3��[��u�U6u�lN8�C|�,ҔL?Df9�s�T�N/#}8���k-�H�����5~�yL��������ذ��̨ܻ�1���SfW��Z��\}�zs�e�j)>��z86lme����꼽��44���,�:[�`N@�.NNI:�v�R�|$^ �p6�����Fh�Mː�i�:��/�ŋ5$wv�*���ȶa�^�ü6�!0(��s��o^i��[��P��*��%�xo�ElƆX�������^:�mU��Xd[�Y��w����W��x���@�a�ݓ�V������W��-P+�������:]��G0놔є�ܳZFfnf����� � �
�0�^5�=Y�X2�ȹ��J��&d*C�Q'p�E�Z�+�"{��s�}g{���v�u�;���ɔNŒq/6���=��EH�z��Nw+��̃c�vs�h*�ն���G�'1��ֹ���?ޛ�YIC*w�7�aS�9!��|��d>ٗ-c�==�u��&W��}���jz�y��fzrS'#7Y�Պm�%�R���Vh�%��� ����f�S�}:v��W,���.�K�+}=;y^Q{6�3��W#5�_L�թ�����Y���6/t���V���Qi��8��Z_��:����J>-�S��5c���:z��U�YFu�������x�;�g���ȿw������g+Т+�v���PU���mTM�;xD���ON/����F���E�K�����?v��������;�!��{�Pؔ��\b�����%�3�	�����!�R;.o�-^��g:��Vj���7��;���^ktR�ޘ���+nݷb1�
��xt��V���D&$ݣW���hDwe��q"�Ig�
�A3]%�o9 a!�b�*�3��(��7�������M�6����^�"�=u�l[�`Lŧ�kڛ�ú3�c7�c?,��͇�Q��o��1{���2�'��E�cu�E�=�C8qǹ�k�3����g؃S�����F��8��AX�J|����-f02=&*aL��˃���n�-�k�e둊��S��[f�* f�Qm�������i�����
��B|Q����z�|f�3p�^��(N��l֙�ځ6�{A�E����B��Os�jXP�;ȕ��sZ�0U+�4����h��� �JuUxڥ������VQ;8|�����Nb]f�(�"n��Ð���Ԁ��ɳ)�,��T��=Os�[KV�T��릭�>�T9�3T�y��y�wm2t���e���I�)S�}�Z�*<ˠ}�8wNW�\�v,W9$ҨP���̫h�B�J����Kyn�EO.��������S���i�װ���P�.��-K�{z��{����T��d	��nyng�>�8o���yάz�o��tw�s�|���F*�sR��&GޝFh���ʩl5
��X����<�U�!��f�2z.#����qeݶ5�ˑ4a��f��1Fc׹κ�p��J�n�rVUr)�_
C���__%�,�[���&NJq���.�!�W�&�6H�3Pn�x����GkN���~^�?#�C|qR@�����_S�ۦ��g�����%��k�w;[���뫇���h�G��ܨ�(�#kf���f���h\[��I:æ��B�7s�P���,1��0�!cQh.��n�l_�,����Y�Y����~n�f��Ԏ�/Йۨ�Hf��.�u���K�.ߗ|����I_8+\�a8�����Mcb�S�w3��.�3!���=l��/����A����1�|���\(�����󐙚<�dNtZv�sO.)�<#���y~	��4tS&֝�q�c>�`U��rʙߞ�n�N�QgN�Hc�씆�_[[��%�^ܺm�rVVv�%$�
O�g[�Kx%ҹ
�������yK��;���]n�靈�3NfH�X��`������`Vޢ�nf�y/Z�������Dxt�jj�m�f]�Lk`�:ފkz7kz�絪�H�����6;���y*�S� �\���#��_L�3��w�HJ��&t���t��.�lG?W���M/C���0S�xjR��[g��=�����ZO����`@�Q�/n�ǎ�I�۪m��Z`�'�Ʊ�j���s��t��5m�� g�[#�}��?-�������9g�|f�\�F�@���wc�P�f�!�|e�x:���Q�s�'
֘��и��\U��j�M�rK˕!��U�Nh�j�np�����*]���Hw�x���:�Р(-{J�s��[{}��{ mia!1�M����Ġ8�S���A��7S)�ߊ��ˏ>ϾN������t0h���b=�h�����TEU��fkq��4N�_Jj�v�zV1�ױ��`Zr��3����s�4�~#����t�l�ﱜ^��HW��!�E�g-�;�X9S<^�fT��XgK�F���]�g���Y��M,�
3v�kG�}o��'���7�̇��X���Gy��R:�Mwi�j�'��H:	�A������R�x�
����tV�l�������ȏ�}�����1�S���T�5��d@M	����;��;N3"��o��}����&A����xgJ��}Z+�@.��E@\��M�{�%�C1��.eߨ�R�f<2s�_��>���n����T?���[>7z�Ṫ�$}������˞D(�'$e�S3sW>q��+�agz2�:�zEM������(�}s�65o�����э����;�ut5�C�(ϔ��������5Oe̻�pä��jO�3��/�٭h#�vT����>Fm���υA�B.��n��Qĵ?JV>����s	�����3L���cf���&���Lö��q�Dg��g�Ni������5�I��:����o=�r�w�ŻJ��M�VnoH�~d��E�i��4��`�F��z���-�b}oy�FD�ʺ~;}�#���Pf�>��\>;�7�=��LӍ�/�7K\�C�c�:�u��	F�#�F܄V+,rQ�)��VY��\UJ��v4FNSM��mu�Q��*��/K$7��_�s(!����Ht[Aή��ݳs�I�*�ʊ�E�P���#���zo#M�NHIB3oF���eɽ0��t
r���d5��ժI�:�Դ1�#׫����]���"�"�m��P���`R���Z�3c6E����	��	���.���G��p�͓q4u�Z�$��B�%�D��hnq���uew<ɡ5�݃K�-��^e��W��$�ſr6N�]��.e���w�h �`� ���Y�.����X��մ΢d�qcrv��=��q��
Y�S|�9Q R$^�Q���WF�o��l�>�Rd��ػ�wpSu�7k�t:5]��-֖��çt�F265��dV8�C��`�C>��Bd���k샍�w]r�(�����37��y�3�C,��e�m`E
�h�|���ҥ�����RJ�PJ�,�E0썮`��Rɠ�ֽ_�fv�d�K��Q�+qd>TD2�>֗Y�N�q��*u[S��u0�H���u�B�_m$�-}���f����겝F#�t��Pn��Y��8���;�ե��
W�JE��7��;Z,Y�ZlluTؙM%`),#]3-[� ��L�9X�yգT����wCy�E�)�����,�L���l��5��o�ֽج{��Y� .LL���*M�0�f��I�T��Wl�`�(>e�蔃>�S��k�m��fv��-m���9OL�G8
�,��M�:�}��,��h�u��>�j�����W�"�v��Q�}7����.R2����� j�.7j��-��b������m���"����Vb��m7���ʻK*�L��QB��v8�xf��n��5�'*Q��'>x���Q��h*���f��!]��
�����a��kk�Ֆ�NN*�PMɽ�[V�����
��u�.P�R��p<s%�K��7C:K��
W�a�;�m�{�X�5�C�X�[1�IľtZ���:�r�;�Z:�S�WԎA�ODP����eq��(�k�A�I"�
�F�]49�L��k;y�P�t�1K$���m����Z�m�Lƕ[:��{��i��R1���|۽�3�]����;y�:G�0i��|���AJy�9wwĶU�D%jj>������߾�����Gw�(��z�F�
SJ֚i��V���EFƊi��l4�J�I�QA������*��ur�m�G"$t<����\C�
B\Ƅ墊B�(Ҏ���)��"
���4��(�@F��T��)^�H�A����H<��ry�+��eb�Ru�)��h�E(�z�ՎKr^��^��'�LF�4(rCAE���Ju��EFaM�m&�	����䮬99s5����u��9w������y�;2�/���S�������ʄ�7T�
��$S�~j�S�L��w:��K�)2�ehn�Ԯ���~����T�}>
�V�juIh��9�qW]�	�xv�j������	�-Usk_\K`wE�;�{`�嘺e�`-��>׹�>��p��*5��|H��4��F�9�]?2k�,d��R1����\ �U�:|� ���c�|@�jT��l)q>�4�]݉���,���fXO� �1����/��_Y#�<	IP{Z�t�ty����D�Z���5�Gw�尽x2q��%�	�.�ݭ�;��ؗ�~.��6���a��y�W{��[�H���Z2�(S�9����9�q��L���F�Q����̩��?}#.�~����?��n>�?�]}k�L���H��W&�舣=�ݭx�[�n�M+�#_��aR�s�6;E'ֲ���?U�a��Z�r���Ekk0�"&�;
������|��u)�u�@�]8�flџr}�ެ�+������8& {X��&T�vi��R0�a�w^ms���������]jbsݙ�C`����|4�:U�hܼ��՜N����
@h)Y}���s����<o�jl�� '����E0�~���S쯔����0�e¹����A�c�5qyq��){l�բ�u�ۅ��O B�ȗւ��}�l��,��FO��n��=�&�1�L��Ν���M/%���}U�-�s!��Q-/)��k��X̅u[������ϼ���������6PȖW�����Zr>�}͍��Z���l�.ӌq3Z<n�S�;5��)�ä�)�fŇ5x\����E��,�Ϸ��d'u9B��������wJ��\������ .��燏ضmR��9]�ws'�0�}_{�^��m��u�Ld_]SP�^��Nܤ$�a�[��W�-��dWJjw��9�:h��%�ݙ��Xd��b�wOUq�#������T�v�������)��i|d�_�S��f��Փ��.�w(~,��*3��k�H�/Xn(mQB:83�QQ����~�_�l��l���E�h%-dI丐@��B�����CB�r��VOA�"W�=1?o����X L�O�+���)����ќzs�cy�oO4���?
���Y��R�{�^���坫�鞟[����GgCs�"`K��5@fl�U�rik5�_sT�b�4��©L��:�%��U�X?r��E^_/$��<~'���vW���wv��t47��6�'�ދ����W�Ox�x+��8(w�Ǵ��g�{ڟ݄a�p�^��Œ�˄��haFu;K��iؤ���uS�=�I�7�y�C70��`2%��lQz��Θ�i}Η��6=��ڮl��I�������I1��L3wd1y,���yݬ�0����[�E�7��e~͆K�!�V�A⪣�w�9j����1�~�/�Z駞��&�Q�7�|��oj�/XjP�����s����I�m�Uc4�q�
�)��{`$�5E4�I�>�e�x,C4�W}Ƴ���t9��Ͷ�#h��vq=�n�<�+
ۯ6�6�� �Ou�j+Z�ķ1�#&uV{�O�ˀ8��ċ�(:�~%�[�mW��jy��i��r�K����12˦�1��rRV�s;��A�V
�UnF��]���ҟ�0<����ި����
ĪwK-q��%F�aiM�5,��q���%kgVn3*	2n��<<6�L@���k�t���;)��O��=���yR���^$;��k�Ǒ0̦�OSܱsh-�:��:|h��)�t��)��0�TF�:�p����F�K�s@���ݝ�f�F^lj�/�皭ݵ�2n�^w���^�f��"�4�Q`�}��3�����.e��4-�fd��Gj�ƶd����Ǣ�?3.��-����;,�hn�7�����v6C���iս�k�pC�N���]GE�_����\�~�~?�ȯ&�;j�|�1W}pde�Y*:ˋ�FLh��y3b�kByQ�s��h-�1�t\��Z�:�C���q������:�l��}�� ��?%�^	����ӯhV��WrY��s���G&��ֶ�sf1�� �����\�'I�X�ؚcWi4����˜�E�^�:zwv�`E��|���ֲ��L�S�=���1����a#fF��Tn��bǁm0��P/�
��U��0�9Ζ�KGao{F���@7wœ�I�^��F�;��&Pv�[��J��{BG2�&��/�w�v��`�9�7�X�ˬ�[��0s1��{���E�e"��T�a�ҐS�:����H��-N��~���v��zQ��9��5�Je��f�1��cZ���?�G�qc��i��NnJ��2|;�[���+(���aN���)�'�񮚽� ۦ���r	�2��3��=F.�p�΍��é�?�$UұM��.أq�6��l���+�c��w��}�ŹI�H����ţ^�yX��/a��]����*�-g%�ߺNLp(��m��}�����y�|�>���LO��8�i��p�|;��Wc��'�o%������<:�n�d�[�Q=��k��H��w����S�	�W��7��#�yP���|����1Q�x��R�Ly��B0��1��l���'p����T���\�)���X������<2k&�GC�c�r�A�Y43����Tv�-�ׯ��0̷s�w�y�?4s�f�;��������Ȧ^��`���^:��.���5�,w�D�X@�5�^E	���ў�h�-�t9r6w:��D�[�U�|h�r�yv4 ԽM�N5�r��i������!/y<k�]8٤5MYک�}2���F��S�c?���zll�����w�b9���iТTƈ�r��R荾��c�9����
)�Y驦�kE��S�ͮ�6(���}���!����|�x��]a�p��ǟl\�z=�f���6U{%˳��qCz癴M�5Х�{xe���{ۊ�`R�mi��0_m��S-�٫�d�l��S5���a⧯�<�%���;�)�/m��(��Y"��L;\�!H���~���ŵ:�i3�x��ӗ��)�Y@�:%5�ʋi׶]�m�q����jm�f��qᡅ�6��챞]P�7676%��S,�%�5ð�ګu��Ӫ��0��ӻ���#e���Sn��[�Lu�p1���s���~���lo㢶d\*�p���H�o���n\��5�G.����_���=ۊ Z|�.��y��t�[�MK���\)���3b�C�e��:��]'��[�`y�Ǯi�j|m ��7޽�Ԟ�A�x��F���(�*�j�)�Қ(5 ��/#���Ob�u���W�&�\¤Y;�����F��y�&#G[U�l	,D�C��`�]dYV�ѩ@�����H�����i�h�tksH��@���n�r���d^�K4Ve�Q&Z+�"�O?+��D~̓���GF��n�29���v�5;��9��3c9kvwg/mj54Z_®(���x!�k�cny�ጧwm��eR�G��zcz}.���t9���"�%[]u�ʌs7F�hi=�74�p��:a}���9�;1���;��4N���6�N�i��C�MץU���4�q�)���\��X�ȑ�� �7w'�w��b��	��������V���U���
�j�wY{� �o�rY���1Q��o�֫}�z-��NV�����<P�<4eyG[شW&��8 �e����_��V?Wߧ+�[Gˁ��8J����D����8��㮇��+6�)�57���u��,R̚yκm�MN
U�W�Y54����)�j��UU�s��crn��L
��۪�S�7��~$./Ous��ip��>�W�|��0��v;o-fe����j�&����HC;���Y�Ыf�U�u��o�֦Wdc��Y]ρ�9���2�V=��A�v����Y�%����[9���j��x{֑�J͌��=y��u�6��zK�we�����[�h�76�ri����6�X<c��gM'����?�l5>;�j���Q�Y�y	<�QM%�R��uq�y��{΄-=��/�U�:�ͷ��,4��f�1���rǞ��2��;MGћ9Yy�O3s�=�W�x��s�;y3<�7H��/\��߉�ն���'�����}Y�\
��/�5���PYP �U�Kן5>�T�gU[��e=݋��Ys:lc7�N7`Ȁ�t���<��MN��{�O'�DfK��5��ݚ� q��+L
J��| ��o�<>+�.��4����h+���[�5����fT37�'�۟��i�(�m:̯/��
j 8/�����P�V��r��5��q-�vg��s��}�T��g�ڋ�z-�^؆^�E�M>��ʳ�H����۴s��3Gt&w�t�l��jm��;} ����4�R���Z�z�m�MKUukEЖ��'DX#CI���&Tfܴ)EbKQ�pA+�����
u� �/�N�����H$U�yz���:���jo�v�#v�&�#���uLegu&;��v(:s��2�v휗S�n��Ur�u1�QC�1���k[���s�?<��e��==���]�H|�k/L��k!���?rj�������Pu*�k:fm�~xd���[��0�h�a؅�k����x�5��5��_�����P�L�T�y���@��0lznl��Şc��������;M�����+�K�Q�l��'e34x��t��5p�4�»����CCv��z�b���He��P�*#>2΍ᭋ��~u���~�iZ�T�V�T���ϗѥ�'��l�k������t-�и�ǝn��H]�B�#�;:�Ǝ��`�76�~`$�ُBÝ����~����}Iw�&�T�p�S�~?����̣��V�=�,���*���_p�s�(tʕ<\]�ojd��T�߂��/������rF����ό <��l=�$2ɟ���aWۦr:�CQ�v:c�.aK�)g��g�X�K�����]���q�8��<p�0$���b�yWl��6�ж�W�r:'�[�5���)�[��p��_t�أ�}`,t�'5�}[`��鎜�GK}��s��k�1R�*&�L��}�%����?���B��>{��W���ba�>������P���D�7T�6ut��U�A/ŧY�\b��9�\OPj������
�,�8�����ee�k<ҫ�&�Sv(-=Z;3k�|~S(_?��p��|�� b����V�̶�]ã\p�4��ֺ���������?|Z>��%OΡ���S`���6��=�C��T�ݕ��W�C��#�v�y���g�t>�6�"]٫��֋�~����--=����p�2G1ʠ�����%�Ѿ��u}���aӥ�ߋ��;��:{�Ճd�yj��_NIf�Ι��U3_?.�7w����j��П-�Ŵ��/.�4�F�J!��5r�H��n�Y
Jfˇ�s��ǅ��r9�:!�J-�K��ĩ��SJp�b/��8]�O]�)4��U�H�L]�M#���.�����{e>Fm��D+�lS�m~��[3����0ƕ���Բ%��4V��K��<F�ڲ2�`�A��&vVl���Re��z�����ei��c;C<�D,'Ǒk��qL\I}r��Tlc�wkFMZR���"y��2��ˈ��ek(��4��L�-؛R�KB�.k0��P��ɧ۵���+;��n3�E�ÅɁg�|�e��0��Ѫ�ŕ�uN���"��wǣs�"��Q��3vI��\��[�����%Kw}��N�u��<˵��퐕pK���v�U����	ޗl��й��>ִm��e%(j�9�^�U�*o�^�o'����7ǝ�s2xv
���PX���'7q	�ᐾ1+8}��vVV���Mo<ǙG�Q�P��y��Hy{+3;I1x����YY/F�i:�;�n�9pf@��E��n�,�4(�/V*�8�0wBa:�P��]u��Y8#�7B��eҭ)��
���b䉻���Ki⣋�K*���M���]�gXH6fʐW��dOl*ጜ��Vʔ(��r.֛�t.�ϸ�|�YS��|�9�d��E�N��$b)ӵ��]��8-ɠ%:5��j�1n��r�u��Th�V�D�i�X� �=��U��,��qe�x,+�H�����Ы�ZՊ�Z�o7s]_JZ�a�ɉ2ʁͮ(�疦4oIG{��ɇ�˪k��e�����U�@7Q��
�4u[*�N֊�[;M/���<+`�B�832��+�t�1k�B%ۧ@M�Ee�r� d�{����nӍ�xE���$�p�7xrh�4�l��(k��0�)S`t�����Ԑ��B��f�+��_P��qp/�m�]یUL���D�hL�.��-�_Ⱥi�tVl7.��`>��%���8���֞0i0+x{Kh��{#����8�x��`{��\���!6.t]S"S.
��J�9N�e���xӒhN�ي���l�T^�[Bf��J�%i;wpw5�m��m��A���Dĵ��,H-�B��_tT�օq�]��)�b]Ú�U�MD�6��S�ի��ϻ�������B����� ��hv��Þ��*R�V�)�М��4 z����#���:T�6다���䩥y�Q��I�T�BHR��h�Jit%)GP�AJd���A�4<�SHrz���ii��J\���@�N���(4:/n�NA�l�P�� rS��t�������hBp����CT��u� 4!��AI�ꐪZ��˥W�7x���N���4F�淋�^iq��܋Z����,�;F�Z��:M���j��o�q:B ��;b������YNS�ST�i�ۛ}t<Fv{V��8ȶ��\�5
ޙ�&܈8�����M��)ݯ�uƐ���!��9��S')&��ئZC�,� ȩu$7���a�<��b�L��D�����Oa�.��dcLgH�g�ؠ�ӡ��->�r$Q���x��t�Ǚ6X�B�D�NVf��c[[o
��ʯ�.]#�"5�=ö�E�TKe�����<U`G��f����s�E����	�)Jf�����5�}l�FK����Oufq�k�c��Z_���*2䴀�S�iC6Otҧ���D�q�B�B��K��k탶�O��ߪ 
��w�*����]�0�v��7s�V���hG(�8||�1#��V6�z^Y�{g���;0�b�Gs�<�^vƝ����{�p����j<l�v��R웵�Dt��m���cL[D�PY4����������I{v��ojk��t�>hk�4�_rwy��+,�Wp���[ٰ��s� ���2�Fd���{֦6���@YR�W�����[��(�ژ�#0n�L �u�_X����.�Aw]�^u������[E��3e�'Ox�'���o��V�����oGF�7
Vi35'd��ιӺ/-@ �Զ }d����:�=��3^P;��!��&/���~S�'/��*����=)����%��[�ZX37��v����{5��w��5Hl�����Ӯyƕ�eSɪ�<�oc5b�qԭ�Ө�Y�����g�>��R�_a���,�(L�(<\Uj�kP���'Ҳ�{[L=�N3S�~jw)ȸ�!�@�	<6���'o&*������ד���ª��X�Vx���nu_:�V�ѥ�������~g�5ޕ���^7��pX�}��r��g������k�j%���ts�9{�r��u6$;�q�;^j�D���!LIN,��ot�W�<2�Q�윧̩.�+���[W��F�!�R��p�<=u��L��_)p�Oi��. �埃���ҥ��c��z<+Z��x��h����h�W��$��]�ޖv
X��'�j覻N�-"p�C���茊�L#���hNM�v��ن`��R�h���_�[���m��z ֭W:GZ�y���e�i#���}��O�����o�O.���:/#����:r\PO��@퐲�#��4��+ⓖ��'�|�����)  T�'9��V���~[�a1�6T\�A�DJKc�8�w�g�������Mq�O��M�4w��Ha���z6;��r�i��iM5.�T�;"����o����J������s�A�to�8�dN�Y�@�s���ιٹ��2@����|d#C���z柗g,Ѳ��l<���n
L��O���=Z��������	�Aw����]�6�}.���ys�dc]���鄱�6�΍d͠'�T��c��5(�~���t��-6����ߋ �SH��>Q�>ض-\��s���Mu��~����� ���cG��Y[ݰhoCO��gAykZg_�T��|.%���G�����gڃO�	��b�O�4ӯi꼎ֱ\���렯^9��T�N��܆��d��+�2n⭗�L��s��=�;�Ƹj�P����&��Ƅ��[2�)�a5��ߟW\ S�ױ�}S�h�s���t�{X���#���*����N9վ��?~&^>9y�\���v��Z��}C i1��o-�4�(�Wni�;�;��Щ�[�rzɁ���-l�X���}e����pW�M{�ŉޓ>�b��=<�J���@;�P�߰	�lR���i���P.��ʞkE���R--���ހm�H6�[B������݊���jO3*���f۹����Bv����`���n}#"�HQ=������-�F�a���I�G��Q��"��75��(\�.P����cd��kwM(C&�	}`�:�X��]�p�I��dƵ���0��Q��g����}as��9�p�5���0nm��v#^�E�4���D2Nͩ�J�i����݃�2ǜ�������z={$���K���
�3m��-6�����+��~n�����P�6����gn����0ۻ��ލ��E�0�=8�n&��հ�"S��B�C{��	�l �S�f���{X@#4h!ԗ��.�>�9���F
�����~���䧕e�ޮ#ή��xs�5�\k:ޅ�ms��?��MA�^�Nj�&�v�Um3�e�Ƴ�;��(L����:�b_��Λ=��;,	�j)�j�g�pY���89z�.3u�U�Z���d>w�Z��*�;յfW�Q�=�/���x����A9ۍ��t�,͔�ُ;އ��?gg����|�:�D�}��[x����:3[78on�~�c�>-9Z�����_�Zo����ᕪ�U�pF:-��>�>��Ș��'[1</�\��s�m�S��a��>��-��"ة��y���=[xT_K&��΢)��Q��O��ߋ�$:�L�kRy¢ω�)f�a��qK���W�/�_�¾��^e��r� Ș?��lwacX��]�����$�;�l
����	[�ΝU�{�|z��klA��4��Dl�T����c-�ﰐ��	�I�B3�\,M�*^�U�]�w����4�t2�_fH+��Y}끭j:����L�S2�;�}�\����y�=�+�Ah���t�n��d�t˩7N�ʼ/���q�����"J�:^{��T�vAwX�ι�6��H�V0Mk�n����jhYI\��{�=�W�N���ʧ^NmJҝ�7B
e��}܇����*��9y�IL����$:�����7���NU����='�5c�C�O�����5G5�<����N�j���6_v�i��dnL��n"Ź�z�5٤��/:�l�c����nZ��
��R���Ķ�F�11�C�2��S;JP���]@���`dWH���u�;��tJ��Oד������4��;�>6;�wd_��G��]��w+�6?��e-;zr~�*��m�q�qӼ}Ѯ�[3iixM{��c���Ī��]�\�4xڧ�U���x��
�'�����ك|O�vc�=�a72���f5���'b���=��ż�,�p�醪�Ɩ�05;Z��͓�C\�<��������y�ݛ��(+)�i���.���Um�x03�m�{�e�fa�,�M����n&��:��΃�m�U5`���c$����|����u����Ң/�i��Ѫ�Ez��n�3�zhg
�Ȯ��ō��=Kj���Z�K��Հ2:�����J�̕�qݰ�o�(�����a�A�V�V%��qG����k�,�Z���;"P4��!͆��F�+���@~�v�Ow�{����ϥ�\n�����Tiy��g�(}��ﳗv�������'�}9 �r�a�tG�VI�|{�ض�k���^�'�rxP�o?�qWasʖyX�|k&�}壼Pꄍ�5�)N�O}L�ޝ�`ﱝ썋����Y��*���`�,���1�����;����~�p}Z�b֎Ī���A?*������K��q�a'c�Br����~|.�t�)x]��r��?�a V������B-7�!4v��˥Z���~ٍ��nf�����������v�<�z�Ѽ�a�o�2�:�m��X����m�q������=!���K�5��eK8��5s'x;��Iz7�,ZF�P~c{Ӫf9������sE�I��$tskWo���'\�9�����ij���xm�S�:�mM&�����������X����n�A���[R�!=�@/���ၬ.���;�b`��x���v6�嫶���js�X�k!R6(HJ����J����[�y�1�F���ܱ��	���<pa0���2W[yl�ij����~�(����5~8U����+���m��A2��1����*W��p��%X�0AE4k�=��i/l[(��*a��\�͂�Αü�k��Y��5�[Z��Y�r1M��"��Db�ѐD�iw�z�f5=��E[N�gj	4�����q��n���Y5�����ڐ��t�՛U;#"l-��tE7k�D&��%�P|4����&�mŴ��r:-��܈�eW��j�o[wU��V�ÕБNQ�l����06}{%���-�=s�,v�6���p�L̙��X�e�1c�K;sږm1�\��?7qx*�V)��*�O��@�ܯ�ѵ��"ڝ퓜�k��Ĕ��AUT�_�3Me�7���?f}y�ϫ�6�6�E8������^{���YBQ=��ñjRƮ��G�7KKoK�)F2���TO�5P�ιCc�9��A�֟!\��Z����;毩@�;+��[��{�V;z���&��V�
�Mm�o!�D_T��]*ĕ�K�$��:��1�!�qq-���c��ni�]x/w��r޼�ɝ\����J��;���c�.�6ഇ1��^S3l�ȏus�3M��Pn�lov(3=��W��>�H�O�lOİ��j�6���K����tw=ᱭ�~�1�S�ro�S��N6_��,����ٌkO��2u ��G4���=�s���2�73-�?r:]�X먬Vz����ʾ{)5{a�FXh������V�c�0ز/�V�����k;_a�a�69�_X����Bi���Q��pY�	MC'���u�U��ܖj0��8f��̵��x�Ž�����1��&�"_��V�>��y����γ4����z.�����M�2./�a5Pܑv�˻_c$T��ڻCo���t4�����K�<A�Z��i~��n1���ک!S��8�ݙ�,��fq�@�t��Mڄc9|��n���At�n$��֥��v_7�g���I��c�P��˪��<%��?^�勇��P}t�|>�ς���A��a�U�$�1���z<���V�˽7�Eh�P�AyN�7�=�b��ܩ�����9o��8Ҏ�t7��FXn���r�Yf��vj�6��5o^!ZӇ/��/Ô��|fZ_vY�q�V� �0|��,����ξ?T�3��m��\8d�ֻq%@��T蘠����Ԑ`�DT�������ST��x�~|�h�ۋ�KkKo(	!,�F�`ؿuD���SuQܗ^i������5끩�U�3�m�Br�ڽ����s���w�u��:�A�{=�O�F���F�����Z����ݧL5�g(C�y�{�d�c��o��n�=>��3�Q�7���đ ϝ�DJ�v��v��VI�`�n����ٲc<�@���Ls;j{����a��3� �.�+�%���]46dw�ÿt�Ѽ����]�@�ya��F��[K�j�ez�k�wxu����q���oө�[����[���׽�E.���eQ�t������Ǵ�k@�O5h�� �3��R�+�΃�-�[���p�Mh�K,Ev&ԍ$Q�嬲��;�XF�R��ۗ��<��2e�;���>�����]+�{JvEMv���Yۭ�8�
�rO(��.=��S��;��U��U��Ԉ����%����"�̱��es!�J1C���o�e,[l#P
�ѥ��|b���Uڛ�C]��,�Ʈ�ӧ�=í�)D��Ӟ���v�=yJfd����t�t��Ms*ֺu;b(������ӟu� I�i�H}<c��w_�-�����v�{���m�)��t�s�Q���h�`�!t&��.1;��f8gc幷�P�8:r��p>ݳF���.���.D�),����r�8���[�Jj�آҀ�{�mq㌥�K����^�0H����2�lk&j\�9i&�Շ���D��xѸ�h���k��B�N�)�8��K4�tg[�3b):��T�p�dj���&Nڶ7��ԶK�*��r����"��E	+����J}[���9mM-V��|�[F��&0-e�Dh�٫���Z\�4��VMsܷ�E4,�Z}�#�s�����7��ڳ�c�r��]ދ
V��Gz��m�����(��X�XY���PϮ��tN$˻�ڿ�����S������v�Ԟ8��(
D�I��m��a�F�	W8!xV�MdL�$^,D����"���O7�_��+.��찳T�O��կ)E�w%8vN8�o`�|4e�I�_p��������q�-�W���z�T���x�a���w�L�R�wHManƬկ���|�����/N�A(�"(G���$�\9�,ܭ�n�.�ŝ"ǒ��S�f��_<9��A�t�*aN�RcזΞe!�&����/fBd��ޮ�R�ګ�N����J��n��=LJ]��{7`�`��QW�v���P�jX����I��EX�P�aݳZ:����ϧ2񧱇O�a@�V��L�N� �n_lo(�ݮ�[x���@s���ed�G8�+t�c-8�aB�k�]>�/�a�8��&6�����uѾ��U����3�ݩm�%K%��8�"\�2e\l+.����4U�%L���o,�|;�0c{�OT�6�j���fow]���*����{oV�VQ��UAU�UR�s��@�]i9-(s�4��-!��˕�u*h�.�+H��h���B���t<��4 rI��yu)I�4Ѷ
�4����Z4�z��S�y=su'#Gns��=�)h4%PU̚�&��N�����QBrIʵF�ORi
9lC�佧Aԝ�B���kM�l�Q�҅=l��G]F�����	\#m�4b�y&�F��=��(�y�x�9��I�)%yD3��d�tʆ���4���������ㄺX��v:���N��OQ1���Z��Κq�}��W�wH�
ܲj��tPͼ_�_k��JF�?��U+T�Ϟ�����g}�� �_���D�6-�ϕO��g�-U�J�J��$:��.6����'x�����5�8�8��?8��'�ŧ�u����CvV�0��tx3������Nl�ǌcj�Q�3�X�LZ���X�E��.tb>���}��kV����Ys�9�Oa�s}ja�7�.��)�v�I��������Y���z���}}��/�#X�d�ٷ٘w��tcZ�6��ܔ����Y��gV.m�L'*ߵ�5,��}��@�	;Ӎ�ٮ�����s�&�Ͱ�*5�xcS0d���-�����k���;_luL�����c&\}�B��y�n�_�a�4��~BZ��yK���.��х���T�k�@���7Z�S���~>Zh����� �
��>7`W����qF(������4�7v<C3e���gE���<��;��y��'o�U:�����MhU׳�	μW.�P�SKy5]{��\�WD��������8-�c�HNjG�����sNv��q�� k��q-�/!�v��G�u5��ث�#d�N$X4�*)�zC=V].lg;��P왳;��%wPgs��!]�f���/�8vGO��v�3C���S:֎mOo�������л��ۛpC�jf�6��v��������@�� ��P���>��f�N��q���4tl?3��"���GR�JC^�LF��視�{d�&*��u��f�.�瞈,bw2:���ni���[��lq4l�Q���ޣC�栃��0��Ҟ���B!���R�c9-������^[��<I�U�y6Eg /���nN��Q>�:J�O۝쳟��ٮ? ��Be�l���b�:���fH���4�w��q����Iݩ��3� �0IP49ח������0��|���P�]��ݦ�}ϧ>�3^�;�x-"�i{�=x��+V��K�{clUM3��K����
g�nwYt��Q���K"���s��`l��->�MM%�<�}j��sp����R��z)' 2A?Y�俫ՠR�c	MH��c�ѹ��ymdG������ ��Ք��R��ye|1P�*�,� ����f�Pw���tU��n�T�o���'�l-�i�>�=�ܮ�v<�9�x�x4B #A��]݋���՗�i�����w���:��1�6�˔�4ư���V٢kdwWb���|����e�'�����䃴�u7��K\5�E��0	9>k��M������6[�9��Et���ԅl���F2ϛ@�L��D�zN��X#��N����7���XP/e)�:�X����È����+�����)��nW� ���)���>'�`׸�<2yx�_s�ރ�W=y��h�fw�spEi����
����]��a�-���;�>���{����hOC���t�=���RDv`�۝�9��ё[Z�ЩM� Ls<(�o��cs�;�s9��h����������b *��ց��KIx7��'pVi��O//μ��&���2i�*���5p�n�h�W�<x�{(�۪�J��/��!�]�[ru;��n,�7&h�&�q���]���k�h[Ҷ^C��SV��TC����c�� �91���T�[ h^��Y}jI��#6���T�եF{�%�t[.��&�P}��#������i�+�[�O���J{Q.�rK��K�i����f�*]��t�9eo����yH��"�o��um=b���F��&�*	}�SOP�w�5�3y|-r���ڬ{�za�s�Wy���|�N��n=@M���22on�U�b�Bߊ�ge�s��	�ɥ���h`����^�/�������B�1�GL�4�����`ð�.�]�>����&��v��ywd��X���ieoݐ#�k®}͆w_�.X�`&>%ϗ��=ΠT��?rk���n�`0���c�-�m�-�0֠��whm�r��q{���1��Mfc�"� 6$�n�H�1m�񥵥�8EAT��0���E����0�&��ly��]P���1�#�[*0Y4��J����k�B)A�޵�T�K>�n�\(j����4P�h	�����|���oc�߷����``K�Q����ż�S�W3��D��ʭx�{M�D����ʼ�����!A�u�1)f}u.�aj��!q���a��E{82xƺX�_�*��&���DҺ�֋�pew\d��j��C�N����k�Z���\���p��� ��r�\��%���e\�B�j|OV-��@�TP���w���۽��������A����;1���B��c��S� 3������UC����'w��fX_hP�n�~n���t;_?k�B�U�`dV�Xzu�wT_nD�!�Z�[lD�lC��~w�b��8k�ݝFHV�R}��WT��5+�Y�:S(�(�.�qL�
뫚��'���-����M!�؝z�(�舊��*��웅�H�9#i�=��_E{)٫z+���T%�����}r�:�v��A;����X�^H�Ϋ*/��W؆|�W׃U��W;��pŭ+�]�r�ߍt�k�8�������i�M�`�ujH�n�Y�l�T���L�溷�vְ�ؼw������<!<��v{���h�U�y�94����TSm�nW�C�Ka���y.0����Թ�g>,�k�
��f�%^��&-C&����-Dd3Sg�#[q�g;���@Cm�{�	EZ����Av ]��ɲZYՒ7Z���kn�9�1iI�"�/��m)�z�՚	��l�ݺ:��w�4��<͂����6�+j���=��G�����}�r����&3������3��D�;�:Q\]��=uţ�\�"�O�s����P�4}-`_�U�����p�}%��qM�XsL�L=æ�\�߆�`��-�|������?��Yzt]��:��>E���o@Y�v�~O/��D3 �1�'&���W51��v�ʊ�y|�Cg�i��,
�LӃ��i�2����Z6Y�M�S%��z���s�+����}G�ϓ����;����]��Y�ٲ�����쑘�tL��#a���\���v�t�7�&�a\�|_� >'�����غ5z�4yO��o�s�'�X8:IxI�#60r:����%}+
���~��#ҭ���C�ɏ���������.�W)�aM8�s��vh|5�d����y��,�S�����ݑ��!�<f�O��g^�t�K������/9W�z���0~�UA�3�Ϧ����҃�o�ਿQ�6�5%�mu���3um�w���H����y˪�0��#�%��K���e_9���;x9�ېe1�@ƺ.2�Н���]�W�w>�*��h�e�
m�ޝ)ee���_W;��s_=���b�HTf�i�e"�59a5�9�����S�l�`�b4�1�)��6�D'M�03I�/)���SAQm��zmYQF(�sm�8��A7AU�����0��W�����Շت�f4�<�S��}xLkb[x;b��GuF3O��
dTm�2][r,ٔ���ɗ<y��ݷ���+�A>��[���=��r+=Fm�EG�,��,ћ�@����o�,�����4�k��Sk[���,ٖE��7�ĊFy��p[l��q�]������'Y55��}/"�~U��M�+�8e�#"���ξ�YP0Y�Z�P�����"��s>t�b�q���Q��'����>˲���h�'/)N�,��t�@��Ju�����N��e���d&zt��=��(`��l���25$�VU�Ή���k��+�]���;G�׍��F�_7A��@o�����c��hg��j����뾈V�v�ʗ�};E�P)e��7"�11#����n��Rc���r]����.3|`��[u�/�����7�O�5�>��ʾ�,�Ļ���H�������h���x�z�߽��R�@{�����I'��Pq�\;gʘ��l	m��)�yg3G��9��x�cr��i�<��,'�69�s�_+u�u�S� �Ķ}�[_a^�ޣ���Ql��K�7�$�C�	f�e642�{t�&=��&�Kl�.︢��]孇�,':�_��� �~S���~�(^0!L����zg/�vl ��;�?p�P{9ei���ľ�@e�?��i�Uڵ��9����)N���̨\H�ڐ�i����QZ��h7L����5�5�f�}zY}O,20�a~���0*o�Z{dٲ(4\�� �ei�_|Gb^��W]x��,�#�����w��n`���^(_LS5=��
�H�/r���� .;� �n���U搎=��ƒ��(�5W�
3�@���"�C�F)�06V��Sg��QL& ���U����a��oY�=��XE:ͮ��sEB�*��]���c-�tUΠ�Ӈ��0��N��(�MY�T�F���<IꎵI3wY�y�J�������`��q�p�ĥ.m��}[�`MZW�uҫͧ ��¬�cM7��x^F�ӎ� �'����O�M9�D�T�Ss'6Wr�]}l�^nv��Sp��\2暨����X�@�07(J��ce `�j�Lf�z��5�r��w�ͩ�p|k��&�kl o���gE��Ȑ}Ы�z�{g��jѿYl�4v��|��}m j�����ӌ��@=S]�Kge�3{��Z�����P��f�Tw?;ؕ�=̅eW����#��L�6�b���N�["���w;oF�.��2x�]V���x�T�b�jj<�������f�z��8;����7�Hَi}h~t��#���������&�R\����5ӏ��+� �4=<ձ	�Ls?<�x]�޸A�⏙������A���2.F����*����؞K�@-s��2(�WU���'3���H�}ijX�m.��>ضc��Y[�g�i��|�N���hN|�#I)���㟹����3�Mk��'4����ܬ�usR�Z]Dw�l+�UI+W�k�t�_m?íz��3�נ��A�9��\��>����r����.
�;��:��t����� ��h��G��p|k���	�j%g�=m��w{-����L�5���X��y\S��l���9_��3���u�G)��nQ��y!�j�i �q�Se�_�#0�O1��N�!��sM=�X�\��aٸ	�E��o=��H%��-lZe�9�2JWfcg�v_]��#����@�U<ϝ�On�}�9��h���[�vZ�����rΖ6���S��o��_.��4�>Pl>=g����i�V�q�<6u!�Ӄ~p��-�}��v��b7�Z��	��X剑p$�55y�kS]L�o4���WݙH�:��u�:���M�)HX7��ݬZ��9h-�� ����.�^��R��$���tk]Z��>�M��&l��^���
q��d���m���5��O�Çv��Z]Y�@�Fqy�c���uO�> @��������p�8@�k����ٙ�UWP����r����t�=���q����;V�ECө���N�	�]�6(FsqP�yl��Wy�c�W8(ޓX%vM�5gJ6�XJ˖r���p*�d��廬;���nM����u�u�`�*l�Tu��^�Kw��ɣ�:`.d�����S�T�wvNר˝i�5�¹#a��J:5]է��QKݙ�K#�Y�4�d�}wt���u3�]�+g;̦��T���]J��1ف�n��	�!��Z6��$�t~��*��	4UǕ���0W�|��&�U�{��,�!	�(P��:Rnw;���ޛx1����L�v}��9\��m��WX��k����4��}��Ӑ�T��[H��ٱ`�x����*+?U}Y��%1P�9s��P�Gn��cQ�x�� ��ih���>�l:��09���g�-�|8R�,���d(�2�j����vs�]�ĺ�@>�f�O�S8�s��P��T3eb��6�����s����ԥ]�q[7��ٽ��u��V����4�ϰCټ�| Xue��&��`N�
�=C(�
����q���Ẕ:i�C�"�ݺ1��� ��[����8`���.��F�[�5v0����˹�1}Ǫ=W�Wn�����(�TsP�5�g*��0��d���j��}J�w�e�&N���WaŃ��Nݙ�k�|�Aٲ))�"��Y�:\�vw��6vN#�Y�$�L�I�[n�g7dv�7h��(=$s�E�u0��E�t����s�T�RεR�pݑ�/�5�:���r[@1�z��;^��;�b�\E��S�XQ� ;hwT�٤n�V�m�+O������	u�QFcx�w+�uzv�uFqvo6����:i�-D���Ȭ4$b�����W$���Z�i�:L�ڬ3�䦁R��Q��c�2�\�(�ӊ_Y�T��j ��C8������@��u��$^M�++m�	�5��\^��Xᗶ��E*������՘{c��hd��,�.j�gon`gU��hm1�u.?�tyj�}o�g���|�@�Ï�Ρ�@�NH]!&��ٛ.��,ť�a��ϫu���g*s���.��8��F���{u�{J�'w�ؓ�#��/8w��ۮ��FtyZB����!�#��(+�1/&�rG��J ��� �e|�AK˨;G �ĚR��k�(NN��`9�]��'EݲQ͍ 4�CE�A�bF���i4�@i4��#�9��T�%������ri9PP����-�P�(.�r@t6΀z��\��4��hM�:Q�4��P�i��
)y':��H�cB������i�4�E �����_\���x6�����gKZ�q��E2���O�������k��'�^�s�7�S7�7��Zw~���;j��fO�L�7�\��������+���Y����}�q&���ݍUM��tp$�4!*�z]Y��]Y��|��W��;e�ۭ}Wz�ל��F��薔�#�Z5�:�Mw�`LW=��]E�f��6�S�;��H�C�ͨAt�z�A��§�{�ӄ���������V��;��<�#9�%@�P��Q�M���>�/A��Fm�zd�ɤ=��]����qg(m�kw%��a����&��v9���c!\�iOmT�u���Jtro����d{"}��WAU�&�TG6��r͹�%��zV���I���YAb���s�����<���|wcF�u��Lm<xeϐ�r�K[&�ѝTKoN��t9�k��R�,,��_� ��n�|�}�����,|ҧ�r"���-��0�2)��_��f�o68O֖�{�<�������*[��LI�B~�R~�[ 7S'uЗV~Z���>G�P�{˞|%]^���CR\�-��V��]�L�ܚe9:+\����V�ͼL����%S���V���֢B��;���Eg�@��S��$ϸw�U˗���;\=�����^��?8=����v�~��n��K���f���o��ccL\�Ql��[>�A4�j�̹Cy��zv�Aʮ�Y���p��Ơ�CL��.�6S��0���fl�;�t�q��*i�>ޚ�`|���~��$��!a��Sl���jlԊz�����QA,�g�5W��>2��}�R=��o��W����Q�[[V��S_�F㈋]}\Yc��1����T>@}��"�}��1$ğ�A�+�b��	����|�폳y:xp���ތ����s�%�8k�ϭ�;(v\�����MRm�-W����7�
%8ΨL�c��G@fu���6a�� RhD;Z�׈��҄`~�t4fZJ�k�^)���o��5�~�(^�Q��r����-�����,�3�'$K,�f�P��~���y|�SNn�"�J�Q�Ξ�����t.�׎*p�ۗ�"�NH�.XF�D��-�X���amza����F��ӡ��k�^g}�*@�� ���=s����_*�t�!r�Ă9pծ�˫y�y�Rĳ��v3��R� 2NI�B"�2��Ia}l��v�[H�ml��F^ԃN��6ߊ���F�U3��wr몝V���=+5&�_[��-��ֺ&1���|��Y����:.��#��ט���g��s$�!�p��-$�4��}�NXWlCvY�#f��=sL��&��E��qs�����DZRsZZӇ4���?��.����Nq˨A�"�>�;��7I����Ծ��\��Su�.��ܰ:��M�	w�]a@�F<�Wow��h����Su_�b�H�G��x'i����Z�u�~�F�.;���Ƽ-�O�<~��Ǟѕ��JCӕ�*F+5�E_���K��/>$}�@f�����]��@�增��ROG��	k��J����������Y�w;3�F3;�IHR���j[rQ��ɱ�}�:���T3��.vލ�&�3w(v�g�wsc|-���;��Itm	�+�FAn� ��ZqCPk.}2pվ~���p<[ew����b��̢9�[=�:�m�>�㣶��b�˂�i�Ӝ�s�9��Q/[Ӎ�Ꮪ�i�;����R �[D�sst:kb���~F!�s���r�O�&Ӻ���Yպ��r+�md���i�K�+#��G�ny�lB`��<C���R�sS����K��M����>4ytl;�u�Y�#M\�<ێ��t
)�w��ۡ�
�iV�SKH��4 �ZZ{u�z�u~���-y�	�W�c:�v.MQ��d(�g���]ہzN��*����E��	�KC��w?�RW��Ѫ]Q���a0ð[�Aen%(�M�vSR{.���a��zQ�����Z�u������||X�puE����C���@�������¾�t�� ��׾g���s՟a��h�9�2�.	�Wp��u�\�I����M�'�LZ�ɞY�r�p���-�)��D�c=�E\�w.c�`F(��O��h��G�=/q{Sv�v� 7`��ޚcWۯO�S�L@�K�Ç�G�Z��\:����'���> ~vXZp[ρ����& yf~�z�O�Oޜ�8��Z�x-�Dn�3��PQS����R��j?++E�LUõh���p��R�A�Fb�� �`�4]Xiss�?��S��|]F�:䷏��%������~��5�fTM�V�k�7�tS�[�)8�����RB�34q�!ۙ��ݘH�ܸ~���v�=g�Z�r�#�sd����j��:f���.�b��#��ik����;�k�
�ý�_�4U�ki ��;���vm�x�!���d�4빠
Hܻ�t�~^���+D����"/L�>k��$p��@|�}�y�����޻�~�~�ʗ�������%�%5��Vtr;�r��Ϯ�M�EK����'{g���Y��3sZ薔�!&�^�.S]�b���_��=�&�]�<��6�5��l�#s�N���������[��(����ɥNvi�"�u�1k*vi�~�[�_ ;~��ps����ب�yx�\���z�����Y�%M�3��A����8�� }d��έ5_Juϟ�x�|*D��[S�c�껂2:�E\����<�Yˇ�\�8v>������T��Z�3�%D����)\^q�s�(��{!.���3n�d�]n�u�����@y[�,�H����C97ٵr<�t�jɸ���g������s���:-�O��t:(\Jkw����Z�X&�xڍb�g����lƫ$�,i�gHMm�0+r:^وn���)����7[��c0���b�RS�e�qa,|�Z۵���	����>���s��/q�X���r�P�׆�ݥ��+a0���������8���K�@}�~I�H�!l5n�f���o��E��	�j@�Mm�d(�r�4��QT�ƴ��k,鮘��aNwQ+296�ED��[U���ͼ�Ş�rzd��[L�&�uI���7�M
k�o�]���ٝX���͍��S�=�e�i
K�Ʉ��,fM��zo�1dZ]�O
�,����6Q�g����|lBX����	�V�����w�~���K1n��ԡ�Xy�k��Ls=H3l�m����ኳtum�B�iq����\4&��Ý�����<�����9�b��?M%�N�4>S~�����cj���fI���M�K�v%]w�g[�D�΍]ǣw
���j���8�D���'�3�������]P�pөۗʩ�Zl=f��8�模�]��ɉ��:._q��Ұ�1谋G�d���O�9��9��?�L�5������̍=]�$�$h�W��j���nF��Bf��$_\�e�ʹ޹�5�du�-�f|��h���r}~~�PJ�U��sa�ߐ�����{�x���#=ӌ�.F�:�g�++oxt2o��Ƚwjj�rD�gFk�ɱߚ� 7y|���zfn}����o~ԑ��.z��0Om�,���fkU�1%��/9�t^c�O5ʕQV�+t�n��~O�~f����d�����u(;�,�;L��Q̻Mʭ���������(x���*�|*_��7k\������㜎j��fnF�z�'U�LZF�]4Ȳ�H��)�a
D�rL�mi���.��Y4����{CO{&e�D���n:��g�X3�������vw�3u����!��	Ey�[Ԙ��a�=��׆8�Z����!�}��G�D�%��c�:��zR�����Y���h��/L��'���.��z�_�]�����W6O�z�=��O�6�)W;�ˬqT����}�N�L3���ԝ�#�٩���MlR���w:i����ӑ��s�>|h)���TKm3�K3l���br���)vuu�y�7���3D�M"�4�s"��y�}0�	��j�j�o���t��~ɬ��}���0��Ι���4��e*;���YF���W{!MV����U�=�����j1�>ם��C�����By�z8�]!�{�ڹ�_^v#�򅞊�<Vc��a��/�T[D�ܖ澘��.��߱D7'nq�CG=[t4������a�Koz��_Y��J�P`� 7�O���s�.{նþ�R�Q��	����E
����m="�2FҊk.�V:C5q���a���a;Zf��k|lnSޑ`X�\ ��
���!���1슷W��3�O7vY��ɬ\HP��.CGl�;�4��U��[�<ju�<|��P�s�}��#fF����{�>s����3-�g�L������p*J�a��LYwHj����(�fX��Y��i�S��L��;�sdO���\��,e髉jY�8�o%�:�%M֗u�@�k:lZF���#��kf��[�$��r�Oi�wJ��Յ��"ڏ�L����}��@-��oX����Y�-&�k$Dk�;����$n6��j9�v�uF��k���e'YA�S�oV���j���c%��kL����o�]����ӄ�H�o v��S�o��v;1dֳ^vPi�8�N7o�@���:o*��A���w�	�n=	�<1W�_|�S�uL�+��jnb�Ol�b���D9x�8Ĉ���a\ Ͱƶ-���\������=Af�|`p���k�xe��>���w������$9�O^.ȥAu�s3�r��X�y����4��{oz_���Z^��&���we�23d�wW�һ�6l�f�h�¥��R�L��v��m�SJG�tKw;6����ha�ǫ6{�[����x����aȩ���B߿R������)��?;e�ܜ���t��P���kn�GV���x/s�><"K�f~L_�c!���uf�fR�됃�5��]71�c���.3�Y�u����ۍ���-���4�R �pc����uLdw׼K�����r��v��\�6��E�+�EZ�\3-�Ǝ$o����<7��&��z!2�{	�O�����i�YAS%�V����nv��?>\�cGk��F<��%�lsW��߽��~H��i�1�[p�Ƕߓ[r1-<���C���,�=S��k1И怌[	�6ӆ�aк�v���ˣ$5�C��z/���g"���F�`���9�?o�@���":'.�r�셥ٷ_�E�W�>�n��y�d�؟����xT2�\��sZ[��ݻ�tct�r7v/ƣ^�pr���lc:~h���(~��ڸGc.�,F=y�<MIx.?�/�@njT�eA�C���'���S�:��U���2�o|a4bV)��ذ��5�����-�!�@f���V��:j#���V����kGds�
5��֜S��O�:���k7����7���6�ݠ�3^�Ʀ�x�.�����'3����H�i��UUR�/�M�QK���������T@S�:��Ew���gy��y �{^7�>����۸u� *��C�R8�#���B$�".���d@y(�x��@xBiQ JQĪ��"���o�S�|	�c��u�M���
  rD?1|o���7����Go�����~����{��*"�����&(�����"���b�)�*���� ��b ���(������(��*�h�I�("��*�*"����")�H����"���*"�i�(�)�&**�����j�b����$�����j����j��*�����f*""��	*h������"*���&j��)��"���**���(� ��*������**""�����"������(�����������)�* �˪��O�Dp�`�Vnf���]�jBv�
��;R{���K�����{�IA$AETEME2$IA"TR�A�2BKE-S$QJA-!Ĕ�%E4A4KEE�D�0DT%UI0��CSC5$�4UD��3I�S0T@�ԑIUQASEHL�P�EE5D�CQSK��ERAKM15�$10UEL�T�y���c���*�
�~�}��G_���%�ؠ(
��wUU?�2�&^k��˯�?<0�?˸?b�]�@_��?������'�=��X���330��}/���%����<��^ߘ8@w~���z:�>�.�@_K��v�	���I����A�wS���:�,�v�(�A��B���jAT@R�����\��n_��r:4 �~�@�ʀ����AE)@�]U z�8c���$7���/����w��ϣ����� �x��7��P��Ҋ�
���3�����:M����q�=��~��a��Ӗt.��E�Fz�~���ύ[��{>?�' 
����훂}A���;����<<�������G��a���x�N�3_g��rF�t��3��s�S���������>���O�U��Ay��O�B �g����v'
?�8=���O��|@UN�p>�T@S����n=o��FS��zhc���!��vL+�;�����N��>\bI��</�X�'�>5� ��xpP8��w�@�3����w��s���i��/ =��`P�w�c�H9����y8�x�; 
��Axo�}���	�!����G�}�0�#�~�O���?��g�9z�}��:��ft̆fyx�p��{P���0��<3˒X|0�>`�|�{3l/��*�
}g�~]���|�
����>����/ր��H�!@��
 �@*
Х
R R4�@
�P�%*��@#B�@� �P �J�R !B
4�
 P ���B��R�R�*AB ����
R
4��H@@(��"�(��"#H�H"�B�!B"P�J��% �R���(	Ъ4 � �P�PR4 � _˸x�B���S��@_A�������^��/�������P��c_6FL����@i���o���A��?������xװt��k�(���� *x�?����l(�RT��An�:;��>���A��ϐ{1c6������>s4<yf}0���)��~'��|¿;��_��>O����P?@3�Ғw
v����54Ũ<Ł���a�&��v�D��?�`O������|?�rE8P��TS