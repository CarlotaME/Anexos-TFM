BZh91AY&SYL�ۉ߀`pc���"� ����b>            `                                >� T�'  �  y�D�� �   @��(� 4  `�    0@ �    Z     �*�(I$D�UB$B��T
%J�PD�T��P�Q���)!A@ ��QѢ��_oERJP�EEHu�;�kH��+�:��<����K�;���q wn�Z�N��*xz��8�V��     u�^t�u(>C��C�CsҪ�xj���uR�p�6����1�` 9�h�\�c]����������Э�=��  �} ����
�p*�
�"(P���}�
w}����޷�^�\��� �;��C�����;�����>Cý/��ҍy;�}�MiCg�o�оJ7gG����8 P�.�*EJ������������}�����R��}�A�W{��t��Ͼ�@}T����(�} ݎ_@�W�q���s�X>�   �	�EU*�n�)*���$;j����M}h�;�� �C�K� i۞��<͞lֆ�i� �h��t�Ǡ��R�� {��8 ( {�T�V۽ �9Jt��T�� �����CO3�C�:�!�g=R��Gv�U4�jWZ���{  
  ��w �y�I*$�T�!I"�| o�>��4��n�� �zz��s ��V`�c�C��{z
O<�W�c���
  _|
K�}�н�@y���.�s�H�8�z���g@z�<��{�h�#�T=`  ݐy��@�!UB�"�B�eE�v5��������G�yE -���W`�������u�RW�N�(���
( ��>�p}��g ��%D�G��9���r��w�"< � �z��&#A� �       �� R�@�&i` L�T�&�IR�      Lʕ(�T�      O"��H      �$ꨚ�1M�=@ ѠU4I�I*�@4    ~?���_����_�����7�����<ǿ|z=����҂���o�R�W�H�?P�������_������
�?���m���U��	���	)^����1���~&?3?#_���oFq�5Ƹ��1ƸӍ���W�8���3�q��q��k��q�2�8�s�.1Ưc.5Ɯk�q�1Ɠ���4��A�e_&K���0�ej�4�2�2�4h8�q��P�J�*�R��U�C�WW�1\i\j�0��8Ƚ2�5.1\`q�q�q���+�+�WW��h8�8�8�^�W�2�4�2��Gj�0=����W2�2��2�1\i^�+�W��C�Qƕƫ���U��*�ƃ�K�)�C�3�Ըʼ5WG�2d8Ը�|ƥƕ�Ԝj�08�q��ʸԸ�q�q�ᣌ�WWW4O�D�Aƪ�J�J�J�)�jq��!�ҸԸ�\i\h8�q�q��j\i�1\`q�q��T�Uq�q�11��ʸ�q��(�Iq�q��UƫWWW�4i\h�Ҹ�q����q���+����W.2X��8�\b��q���q��UƉƪxn08�\b�Ҹ�q�|��2e\j�5.2�5Wj\b�R�Aƕ�+�K�U�+���1\b��q�q�sJ�J�P�Q{5.2�5W������#�Kсƕƪ�!�+�IƇ���J�J�h8Ҹ�q�q�q�q��+��q���q�����%ƃ�'��ƕ�U��8��A�U�U�U�U�+��ȼ4e\d\j�4\`q�q���q�8��J�R�ƪ�ơƤ�K�#�K�+�K�Wj��	��a{q����"�D{�4�5Wz5h8�q�q�q�|�d��\oc���U��s*�R�!ƪ�P�3�GW�5W��q��Tq��.0d�2.2���ƣ.5N2�aq�q��I�K�N5.5N1{�j\h�Ը�{��Ɓ����\e\e\j����)�N08Ҹ�q���q���q�8�q�q�q��N5ƾMƼ3�q�5Ƹ��/�N3�\k��\g�N3�<1���q�5Ƹ�5�q�3�q�q��&�1�k�q�q�4���q�����.5�=��.0�/cS�N4�\g�\k�q�lg�g�\iƜc�q�5Ƹ��k��\g��\k�q��_&�k�q�1�8��8�k�iƜg�\g��8��k��k�q��c�q�3�q�3�q�3�q�k��7ƽ�8�Ƹ�Ƹ��8�5Ƹ���2��5Ƹ�Ƹ��q��k�q�3�8��3����8��8�5Ƽ7�\eƸ�1�g�q�5�q�c��\g�z1Ǝ5q�k��7�\k�q�q��|��G�N4�xg�8��\i�k��g��.5Ɯc�|�gѮ3�q�5ƾq�5Ƹ�c�������� M�� �>��d�(��lσ�$��e8����l���6]��,ԦNls;ǻ8�09���Z�J3o`ܷ[̅`k�N�ݛ��L�-�i����r<Z�㒷(���0���z�v٤<�Z=\�`ٹ��\���0f��laGJ�YO��Cz��-���7x�9�Ӷ�'�^Mܸf*�ݬ��r$A���w(�5�mJ�:&3׎G���so=��7�����x�b��]�i5;�ɻ6��mZ�;�f�F���aT�G`���KSmg:��+Ǜ��l��S�V��oe���9�ŷ_f]�zL�gqHc�ГU8�f�y�Iv�xfb8�M,�Xs��hzH�f
Vrג`��w#4��
���8%�F�h�.H'l��gT�{1-�r ��"��i8�qŚ�=fI���:��o4�k��5��	/	ŉH��w9��?�Jn��2֚���?X���B�P�/Pĵ�9�ιi�	����u�vv�$�n��K[pU�L�/t�j@���d4�V��0�[;V�MU���{�y<����0vD��Vƅˍ��5���ꋹD�;Mp8����;�^L�Ȳ[�����5�߻M���zR���4<'l�q��g.�&��X�L�1�8��}0�"#��7�v����y���;��Z��'^tRrՌ�F�]�؏��i���&:U�Z{�t�d�ُ��.e�O[�l���ǌM�/�r
��`;�V}����%��w��Av��Q�����ʎ�J��@�`4�Vwm��0�*�z�%E�kw����<�Be��<��f��W�ҵ��5�z�P0��\�b�֥�;�]��Rә������Ym�~�J���^�?d�3&�39��tP�3L�����q'7�ҲG;:u���D�܊j���)���R{MK���Bm[ynu��9�;`}�z���t���D�h�p%�����z���<ص�� ��Gmܛ�a�A|�o4����Z���V�Q�sW������v�ˣz�a0��jQJ%\������]�3X�nhZLd�:3/i�[���q��<,�ÌiAm(R��ѢzZme}wk��Rm��{g]۶n}��#��m|���m���z�#�%	s����!�v	��CF<�}y�aM]�w��wNq�XFmx��a��Yd�vh����.r������{.��|#�e5a�+��'#~Q5%ᚕ�d�4�f���푓�eP�p��y��m�.g#�e7���~��P��">�.�5��D��un �� �/�&�ŷ�ع��74���w����I�DΊK�M e8�7��Xa)�>y����یgi��$�iew
h�{���+�k6r��0��Pt��.�����Y��oZj�S��\�"9�H/p���`d�c��;���@�g#�L�ݸ�ϴ�1���Gn�bN��N��3f�˼�-ܹ�N��-ݢ�Q�{�<��eq,J��L�u\��n؞g	�!۴4�2M�cՆV�����V��q����u-�37r�r�ݣ���Ur:�	�'P��
d��p�1q,��95��D���3��r�"dHv'�\����#��:ŴSz"����:
̰yc%�L01��a�raz����9����v������Բ�,�-�)�Yg��f���󷸮r�Z���8����qF�:�.�,h���s좥��wGrݎ�	�^��gO�f]�f{Ga������Lw�v-��������=����I;y�HA!�`#��3�8�r��3�L��s�X�w����ʲ�kZVn#�q��I�����V�uMG��tЦ%�OY�'�n>�`������t�r�yv1�7ps��iӱ��yK�%�֣��m�3�cK�t)�9���.n��=C��ⳳn���5�]�*�$uiVw�n �DapG�;c\��w�QXsTSQQ����C�]ň�&Y�)/D8Z3\�������q��9���",h�U��Y�',�[`�5}��c��:Nm�����ipS�*���v��i�i�(��n/oN�]��F��띺7BFq�E�F�'fv���:����#�;���͘{O�ڢS&}S�w��5����H����q���ҩ;�M�:�&'�o�y�Ծ�E��fb[��Rqs�sw�`�'�o\P�W����Αm-�[ ��%`�5�è����'��`ee̓C�'�ւ95C�3�ӌl���9��n�����gϓ�b�á�Q�V��Ͱ��9��ky��צ����\7��W�s�W�`��){�Om]Ե�4�wb��K��мV�a��Y��z�����D���E��Cw��%�e�9��qvD�\��M
�[�Y�s�pƺM�޶tԡ�%P���X$��ތ�Z��w����<��u\;�7r�[�Ė�������C��f�����f�*X:=z�H�'Ϡ{7d�ۅL}F�-�r������c����\wb]j�0^;D�7�Y�L�&��:N٤Ÿtt%�/.:�ĒہՎ[/ܛ[sY:�����EL̓����{�I~ѡ�x�L��^nW��P�|����-��(�#(�����{F����a��s�A2�ϟ';S��BK'&�FX�&Nds��wQ��2<}Uߙ�[�=��s��W$��w3�B�ٚե�zr���ܲ����P�=���Fq�z�F[�އ���.��i��n��x#��xBfa�ݺ�ÙB�7O^���Mִ�V��"�9�&TsFb�����Z�Ψ3��rW5��vB��t#����屎��2�NG9n���wZz�\�Ҩ��������U�7k�"r�΢v�u��ks����{w^8c��:+�k��0,Or�8�.L�˭kY.�\�[5��fAt�Ù����k�ޕ$Jט'	�E�똆.!{�۟`$\�ʋ��ak�m�ڻ!���1��uj\U7j���}J�am�]^U�NBokx�s^GFi�ū�F�ȯ<]�0�����yi��'1r�]�w�]�x y!v_5�sIr!m�;4�F�,���PTk���'ud�Ϧϣ�4�x�kM�������n��#�c,)J�n�\����i�S}ِo��ޙZ}�jq��Ϲ���_qV"Ҹ�˫J𻙁��켖�s%�5^����g�X#�c��vt�4Ê��z�[	���� !w�.;ydyݐY�j���t}���v�yg��N�:�Nd��6G���$��9�{7s�qY�	}{3NM���[+/l�7ׇ�u�����g�.������w\aC��ȱ��9-�������8��I��B���;5��!w�\��ĭ�>y�󃓳DpntdV����}�&­竚xM-��ZŸd�Ni��F�mӋ�q�i������m<VL����[�Gx�&��H7z<�v��^6%>j��Cå0Y+h�$�-W�wT��you[�NԜ���%�a�&s\���sQ��$uvE�c�s������Ӟג���s�P�TD���u�Kt֬��p�i����ًA�m��3�{��zÛ1n.e��sy��Ϥs���6�n\�p���;���9�w�6\]u� ��c߲�'�f�;���"Z�&�`Ņ�\	gn�P̝�[�o[66ʪ�|Y|�7�B^�p5,�6��c�=�껷nS���s{�R�u^e�Jc�=���d����=Fٜ�p&�/}t�wy�n
Z�n&WL4W��hV�;ٰe˙�n&Z]���iӪ�'2��S�;��ĥ�<��^vv"�[x'p���0�ךG8�@�&c��ĴcڇU��+8�o�Ly�Hc�-,���MK:p��4vŊ'Z�v�'?�%r��c�pN\C���C���>��G.��.�.�V���6r5����2��Κ��nv���,��<L����"�.�Ac�&mލ���d�a�k�R����吃�v��7_�7��}��2n�m�.Ѥ�x��u41q��f�y���U�(���E��I�r@��H*7��I�c��]5��7�θ�G�[�bڶc��}X���Vv��P��̳�ݑ'w4s�THQ\��Ǣ�����V���L����X�+Ւ���0vb�C��0'1�m˸xdâ\�ۓ�̐<gQ-�0�V�puKti���[��*��;ft�$��a��7`k,t�qy�c�7ob�4�������cRy��6W�N���to��8\��D��(�^�G<0{��]p��K��3)�Ed�j0��2aA�Q����[��=v�C�3V���wv�\���v9W]�yL?9����u�΄��u͛y�`6R@p�Bg]��[4�X����9�c"�*p�=ٻ4kRf�I�+7��u�=õ
Ukm:�ud�0Eq�zw#�g)�U[���b˖飃�p�#��Y�9�L�>����(���㋗jD��z�� �����-L#����m6���M�=w,�3Q|�<3fI�9^�3�R,�vX*f@��:�F����J�Y9Q�;�8^����[�#��)�ԼM]����r���#Ns9bJ;�PLY8]���Pr�N;��i�ؗwq��;w�	�'N��|�lѼ��'��O����6�>��)���Z��>f�#5v�z�ft'jvW�Of�٭b�ذ��wS;_[�:vݻ#ܸ��>B d��`�㣖�s
|/%������^|�9�MCP�/s���.���Kp��ed��,nf�ЁJ�7,:4�[�3pu�Nk[�1U6v}��X�;�nWyә��]�d䠽�r���_ݑ�[�9=[Cґ��s}nn���H�q�ϳk��Ƭ�stp��O�ϒ�ȊN�Y��'3	���U�q�s(���������e�(n�
��L]�63�iU����Î��ڏ.S
{��f�V�����e�NIZ&�ᛰ��c#U�TFw%�Z�֮)I=���iř��RZ���U���d�g_���wtfL�
䔣�M��h�,�vHt���$t.:��bܻ� ��vK��[���M�c_zP���T�
�[ّ��>�c�N�W_Y��9r-��]7���0s)
4\�f��M�84�\H�ή�t��^���rk�Fe9�u݆���om7�14���5�2�������6�pᐾ�:�W���e}��ʲ�R�k��ɖ8�%���s���k�'0�^fuը�ݲw�̘��ò�3�0ާ��,��.��R1S�6Uk��"ySSW�6q�l>����k7e�j�tǸ���uv�j������H��s>z^�+�<Ɣ¤�'J�wf�!\�'��U�W�z�E��n��sSڢ�0��?��5�Cy���Yg߱���#1:�#v���6N�:�3��#��������E��GOt}�/T�Nᓯf����Wt�%��$ٹή�îr�%��e�bO>Է��#�HJ��n��LrwW��#7�P�0�d��	���-�Y�t%�.2օ��9ʗgQFv�eL����TRߢ�ؑ�k�};�4�ˑ�Ai�K9��Kr	{a�3]�Y�b��T���+��8^{�۹c�ѳ�J�â���`�l�ׁhY�q��Ͼz7h�t+F�\8PV�pEF48���D�H-�i�@�H��fPMA������Cd-?2�*���Ț~81 ���?+���G�HrЕ@a��>�,�&5 �(���6��(%�����hǒٸ�8�����xק�>�����a�����#�H8��/~��Z_�P�B�����TA��}�t�@فb�+��b0V�hdAR2�@�B\c�Ϩ�@��&"�"!����,�K�ɁR2`Ԃ�D�}���E�� ���ab/�[($�r�(�	��F�<x,b�TJD�0Q7tL@����#����g��c kA,LϤ���R���T�@�𨎄d#�E�7�88Dy�n�!�O�t&��
�H�W������!�_��;�l#����!O�D~�6!��:2hk�LA��=�?�*�oұ�=�"e��T3O̎vϯ�0eC0l�h���t�IP��lu�<)x+>XcM��	����C�
!hŃ,��v��v����C��u���-���5�=���fPՀ�����|U��Gd�-�*1`küGc|7 ���b{�چR1���%����!��/�����K��,����8w�ăP!"��6!�Ԥ<�}�W�lJ��8|[Q���4xH�z�
Q��2 d@9���e����&=�-�J�0$�b�#��z��`𩈨� �b1�c��#*E�����/Z󵈰n!Ɔ��BPx��W�'��7<c���b�a)�5�"J-�sBO��e�s��C׆����~p�P�F!�"$��hɃт�A�~8��<`�ǌ	��_`�����<���z3�΢���8<0{�}���3�~T�Lub�b�>~��FH!`�:��GM���j����U���T@KDt!xǤȢ��хPx��C�y�b@�#�l�nA��������ω��
����v�(�~LL�wE8,�*����6�z `��!'�_�Pvh6
P�|~�1�`E�H��M�+#bP�����{�a�L>���e!S�ņ��`����7P��D�S�ϛAG�bV$�B*�؂����a���7��J!ˆL����h8�Lac�T�^RCތG�>kv6mЦ��DSb++�% &������{��/��c��_ƻ���|O�M���V�&ʪ�6���[+aF�&�6*�6[H�T�[R�ж�m@ڥ��h��l��6�������T�R�Rl����6@�T��!�["�m����V�6�l�[mB���I����h[P�[(6�
؛E[%�����Ҧ�ldڣiʣ`ٲ!��)�-��V�ک�KbVГiM����dSeU6��A��J��[�<Dm�=Dm�-1Ѷ0�m#i�|�Ǌ�<lF�i�[Kh�[lm��D>x٤x��x�kF��i�c�4�YlCKDil-i�!��F4�"1hű�F��������-���CB��1h�h�Db�i��FDx�1�ZxcKi�-���#ű��h�cH�YkY���"�h�����H�K[H�H�ih�H�i��4�b4��la��[m4�զ��4�Z4���F1��ű�"1���1�����m#M"1h�"ȍ"ֲ4hƖam-lZ1d"1Ɩb�������M��cE��Ŵ�D[�#1�,�1�Z-m0�І"0�H��Ki��CH��DcL4���Y�cO\x���m-���4��K[�cHa�[Kh�1m"ж�g�[Ƌx�ilGZxh�[�R���kh�š1��h`<G-��2�>�I",�PY��S�n��.f� ��a��{^�ƻ�����F���B�D&��60��K���Ko��R�	�,Ĭ��Tce���(Ͳ�XY�̰5R����m [��ur$�0B�nn�6�`�W7#M�f�4]nB+̩	�[�v��	�����H]���ȝf�$o��B�ҡ�t4	�M��v���e�'��&����ċq�כ�� ��r��3j�e뇍��E�!o���~Ͽ�^z�=��^MUI���""}~�_}��=���ߨ  ��>����*?LjI�����N�	h1��F9�e�)�(�Tֵܾ? ��q��^�|�^@��՘��=�&n��Γ�S�9����3���h�uS�=ի�����*���A�x�p�����پɿ'0A����Ł�Q��(Զ%u�ey�P�f�deI��ǫ����l���Y��^`�W�"�ڷ��������usiY'�������2ƄCJgi!kAh;�qʷ[��Q��KFg�skk��̚�|yu�W��zp�sΚ7_�Q�rx�e�n,��݇��I��t�7�N��݄6=��4j�_��VއJla�z/�����n��^}�r��nڮbA�>�>L���S��ʋ��uܹ��v�v�'��s�=��F�f�'���(�>�~�_t��xc>�x�h�)�)'�o���>��e�se��;k�f�sr�ɱ�:�5r�p��1�o?$����IjA�!����e]K�L�DT!�-0��bUYyXC{O������fk�˹�.ޯ�>�����-D��a���u����>��K�ΞB9x�����T.6�N�ny.uaܣx���]����zx�9Q�^��N����f��
$��}es2,2�;��ԏ�Z���y�瞽�Ӈ��YgHt��ӧN�=:t�N�:t�ӧ�N��ӧN�:t���ӧN�:t�ӣ�N�:t鳧N�t�ӧN�6t���:t飧N��w�m�T�}��^����S~������N��#Tx��v�(�D��y�N��*�(~�e���u/�q�9���3�=��gl9��y��*��3{����vE��tU��3�s��x���?@�����B\���(�����0����R�w�P��v�=.fo��窭5�ק����b>+�㖨�3/g�FWi>��i�R�}=��i�6^��_!�1��h應^㝇:�g��yΘ�/{�Ƶe�|د7~R�q�'˘9��>0����c=�1=�~E��w���Y|���Y�{���z��4{o{th��[&�����o�}�S�e�s������<;����݇��{isE*�t��(??M���8q��I3���C(������e��wS"�y>C��y�%c��z��!�����f���}|M�ى8�_mNb^v�nqw	�������+G)���^پ�P_N�b�u�^b��v�ۏ�fu�ܓ.��Оc{�I�I�q���{%���x�>g���p�<)�.��N.{����ef'�~`�J��.�A��K��UE{�.���ޙ�g}�W|Ç,�͝:aӧN�:l�ӥ�:t�ӧN:t��N�:t�çHt�ӧN�:ztt�ӧN�:p��Ν:t�ӧN:YӧN�:xt鳙ɬj��Ζ�W���\�������{��%O-�j��7R�%��ZV�xTv�~�9΁&r����|s���O�_�	��
8�\d�ߧ�����F�s�8�Op�{��c��)������c���y�O�H���<c��\�������ǳ�}�p�2!�"~Y�B;'
3;nOIv�n��t��E#��k�������!���8�1e=� y���)l��y=kP7��\%���}���#�x��+������c�.��e�������]>�>��{0� �Jב�}�����a��C���
��}���`:������t�8����T��9��0̀���c��_Ah'�s�|3-�L}�TFyy�u([л(�=+��޹y���i�{�ѐL&(���`HfDK^Q������|Ys�� �z��kF����mcL �����OI�x��P��#��kA�ۃy�C�����	�?a�f��:u��tp�>n9�p�0>9As��|��~��ejؒD��q�}��&Y� �a��Z��]k�0N#<���uB0� >a���ؗ�9���z-:�f���`��?/��S#�Y:r�>m�nr��.���o��
V�$�^���L��qrÝ�;���n����OW�?g��n�o����u9m����X�_)W���0?��!�Ai K~s�s�ن��Yg�N�:t�ӧ�N�:aӧN�:l�ӧL:t�ӧM�:t��N�:t�çHt�ӧN�:ztt�ӧN�:t��ӧN�:t���+9w׺�;����?t�};X[��7���ڸ���A�Z�^�J���5x=�����DG��	�x�z���ဌ�1�ӣ�ܼ��L\z���];��<�A�|X0��>�ǽ%nN�\ቁ�k3F���Gy�v��w�f{�!��J�ɄWQ��S=�d���/=���d�� b}���mp�{�{�wuT�z5eM���/�Pr�|����[z>����_P��V�/�)OE�Ңc-�aŞ����C¨�L�x��_���g���Z��u�e�������i�$�ΐŗ۱n��R�c6�O���W�JՔx����#�����W^�{wv�����϶�9���s�$��l<�S��<Qx�C��rb�%k�z2�Y�Y=�p��zn�r�9�zsp^��7m������NS�>�a����f?\���QJ�_����=��[�=v{2g��	d��5)��8.��o�a���rqۮ���m �S�3��#���|"���S��#��D������w<>��9� �N��e��RfN��,#y�Н	i����ۼ=���^��{Yjh�pK0{�c-x��stg�5�w}�
a�ݾ��!� '�y�$��V�Ӿ �F}�GEp��w��1gX1��D݋��1��w�����\���d;�������< ���ӧO�:t�ӧN�4t�ӧO�:t飧N�:xt�Ӧ:t�ӦΝ:tçN�:t��ӧN�:t�ӧGN�:t�ӧn\�V�(���{�7�K�9�Wb�o^�����nfx��zt]���C��KE�
�]�}� _K���Ǯ�B��)���mS�Ҽp;؝�7��t��q�����c�=<P87��.�R���+�΋�x}��4},���S[�e������a���wT��h�5���}j�ֻû�����)���'�N��}�{^sl���*fY�8ٟS���ܩ��������{���]��(Gޞj ��&���-�^�55Eঋ�ӻ�zN�/M������׬����?wȼ�B��zq��`ޏ��X�^W"3��sW�2�8Ggu>�o-���j	y�X�}��ζ,�������W���f	iC�~߽����8�z��ᨥ{+K��w�o��mt`���ø���ˎO4<�6@_m,d�oz��sȍ��ï��G�M+ݛ��2u�Q�d\��+�ќ��δc���z�,7�V83k#pga��.���\�8{U_���,Ćq4���d@��.ν��U~�����'r�tp+��ׄ=9�ۅ蠋�=}��k�g�#;���/ذM��7ẍ|���=���#� ��+�x^YuQ��3ݸ���~�q��z}��?z;���˞�������ѳ��,���ӧM�:tçN�:t鳧N�t�ӧN�:t飧N�:h�ӧN�:t�N�:t鳣�N�:t�ӧN�!ӧN�:t�Jݰv�y�����{��Z�|���`O�{�&}*��<���<�҃�#����K�U�X^�=�g�C�:L�<�]��V���ׁz�=�����$�����n�i��N��[Kp��S��=�u�Y�7�^���jNA��6��p̾���m��w��{n���_C[FyǊoA>�o*��+��W{���a^{�{5=������&c{�{�������d�QH�`'�(wr���Z�]��a���|&�.��s�n�p�fկ�����K݇�D�C"Ӱ��R��3�8��CǱ��e�z�]��I�i��1Ȳ���&�j't����j��*���۔;0�j��N��@�{4�3������Z[Ҧ�&�p{ϣ�r�pB�Y܆a��<r{�gO���P�yk����^٧��c�{}L��y]�6q<��7��r�m���qN?3(�\�:�H̊��^��2���j�.�5��/:.��z|�>�y=皝F_E��K�A�x��"𖷆����aV��0�-JS��Ͼ�o!����>H���-*Tb��63���ەH��{���}��5�3�Y�x��� ��,��ӧN�8t�gN�:t�ӧ�,�ӧN�:l�Ӧ:t��GN�:t��ӧN�:t�ӧ�N��ӧN�:t��ӥ�:t����I��hꞘ7�Ԡ;���cϲg�m�:��l���]�=�9w�^��ͽ��<|��fy#|{|5y>oΆ��pe���4(���/\���D&,�xRN��[B�&tw�
��秔�j�o�f��؈����|gsti!��yg��`V"K�L�Y���4<�<�I1���gK�O×���7�nd7�P�<B`ﳻ�d�����%�=�p鹃˶����Mw�fx&N5v���q���xh�F�<��J��7���G����ew�X��&3F����ݘf8W��éE;�\�P��T�7��%�}�-Z���*{�^X�%���9�:��_�4��܌��0�#2��g�l�4��}���m����<��^{��U7Y��_9=���7�}�X=�?c���^$�������5��������K�'$�WX.���v��|T���S@=/�'��������k"�n�W����oy��{qt�l7�OR����g��O�C����b���r�{�ێ�ך!�~�
+�>�2��iQw{������r�؇�&�A�����v3�o�[������N�YfΝ:t�ӧ�Ht�ӧN�:t���:t�ӧN:YӧN�:t�ӧL:t�ӧO�:t�ӧN�t�ӧN�:t�gN�:t�|߸�c^K[Zכ�_A��C�|�g���e�`CWl���f���g}9���N�U�d��XF�����~Ë!۰��a;l����;bcD�|�#��ˍl.��&���'�ޤէ6x�N�� %<��zb�>"?wC��J���|�+��6������E,�R����.����\��[oZ1{��l��JOW��<�G�{fa9����oq}٧mk������s`���ܖx�A�a���},t5��4�ooq~����ÊX��c-&�Uyº�0}�a�Oa���2V̝5�}/��o�#�}��bO���.�7�?I�7l���w^��f�����X
�Rn�^�0t��Lv���{�{�9�=���g��s.����_vd�Ύ���w�|>嘆�$]���p����,��I���|��*��}�<���gnH4��{{��|A��>xM9��;������ѹ��=_Iw�����.;���|���j;7�/��\c#0G}�Y��<�3�E� �a�<1�'Fi5�?[�ďC�s�8��1^�c�!���4��	�D�k=W��\�(;0_�1���x�#��������M�*�G��s8���R�cV�>�|��ɻ�����<4Ce��çN�:t�ӣ�N�:t�ӧN��:t�ӧN�::t�ӧN�:zt�N�:t��gN�0�ӧN�:t�ӧ�N�:aӧN�r����NwZ�ɯ=��|������5��m��$�o������%=�eT`C=��q����Ta�ȸ�LA<*2�k>�+�罠�}Ї��/{ϛ���;/�k�����pKq�c7C�2�|�Uw�?F�����3խn9-�9��.��}�8t#�̭k+�\w7f>/����6�ܘ=;`k�Fk�fgD����B�k=��>>[2ʘ��OC7w٨�7�E�;����s,Y���M����]�ϴ:����ɚϳ�|�0F�n�voq��dɄ��RڳN[��E{�s|4_C����%���f���k���r���w��vv�>�c���TfУ���p�����������'}�{��f_ykSyn*�i��P��Q�t���o�n������=Sř�4���;}��w]��}w�ܽ���-[w�$Z;a��P��ѭ!{W�S~�7/�,�wg��]���n���&罓���V��l�F,i�.>�ɩI�r(�����T�|�y0���;���y���t"��ڭ���>M{4g]w}{
ϼ�9=����.��K����9!�Ww����p�e{�]�3t{���竴\�\Oﾇ�\k����D�,����\�5�Y�^罾����;�3�k�!L2O�^�r���n���#��[�=Þ�N��㗁7�����b��=�	�x��6z�_y�t�̋�K5=ŧ�f3���qv�4��H���Lz�Q+������R:�ө����+m���4�������~�0��B����}ͨv�۞�1�w���g.�n&�)��4�;�_P����y"��a�͍�mS�&��=>G���i�����>�{����|�h��)�(�A��=�|�	��t��N�?�m�'�;n�����J��T���s��>���5��z�(W���9�--���7��G	�l\���벴�E��䞎��k��O���M٘'G���7�=�K�vRT�
\��
iHz�݉-Пl%�r���>1������ޛ�['c�N�R�V����s ×V��;�F*M�ֲ�!3���FVF!^4�q�%_L�3u1��Y��S�ul�d i⽄m����A>o^-G=���&w�a��gs,zW?r�A����8l=���޹ڸ�	k>^����O7��c&���𹫅��̍��}�u�OfX=7d�s�gC�#a��i�j��䷵x�ۻ��N�;�ף�2�4��fs8�/Mw��~����������L�����2~�I�gN���OϽ?>�o�n�b�m\���d J���a)T���)���b�S>�i7�O3�?�}/��Tİ��������� UUUmJ̮ʪ����EX���M�n�Q�t�V�Ύe��R�׉�-\X8M�n�[����n�a�˃Q�))�s�ƴ��fīfD��f6���īCYl�0�db�jj�m;��k��KffC��Y���vkFl��/kb�tM�mu�+�3%k,H��bέ�T��FԠ7i0�5N���F������1�P��e��kN,���Wk�X��V�"�m�.ؖ�n�GX%��sn%�0[a�Z����Q���kbM�	@#��=��:�J3n��ilL4�Վ1[2�ʹ��v�	Bՙ)���^��n��\�H����� lSKF�:���@n�gmɹ�.�"1!�)�lF63K�P��Vm��:U�`�ԍ3s� .!6��*0�+tF���D��)Bڒ6�	�`X�l�K��-*�n�j9�Ȕ5�:�fPeڄB�ԡR�{;\6�4�v��Sa��Z�Q��Rۃ^m�g=��l%,�SR]
���lօ���1�5l�s�P�G8��4��s%&F�R3-�r��Wb�K�ޡ6�4��/,(+f/R�{`��%T�,�.���3	��*le��[[�[SD\K,yu���x �M��x���]5��r��#J�Yek66\M�w1��д�aq-�e6�xt��P��nW1�@�a�E��5V�]�4������gMG���^��ҁ�5���F�-�b�kc�pvR=���
LK/�h<d�D�n���.��'[+(͋�%��4���T��4tvk�X����mkC;`cq0IJیh�-��b(�qB�f�	f��44�B�4ۣڅ�s�sp�9���ٰ�G@;lH�z���B����	����a��#�Gkɿ��<`¥tw[le��Ъ+Rk��T����m�F򘼧[�a6t���IfPb�vF�j66�.�1!v�5��A��2ޭ���&E�g56�2��-bi��a������"0�"Jg�S��aM�]�h"���J�3�*f����Sk�
C�����{���ں�U5�:�X�n�̳F��0e`�4ͽQ\FV�IA-ICB���	^�dٰhj����B�\��# �1�glmb9�c)j���i������v��DKI�t�t�K��Y�BW��K��. 歰�[�d�s�]����rKV�l���i�R��)� $��&��ـ"c��+�ѹ�gF�VZl�Kfs��R�MvqIT����06�hR�lt����R]q�<Oz��S�p;u���/S\ؙl�(;m�n]1�3��gV�2�`Љ7V�����."6Z�˝s\�a�F�p�֖.��������Q&���Y�ˬ�5�w��<v#�L��A%U�n�	z[�2��ܵʡn��V3[��#����,ye���Җ�n�DQi=��9n\֪��p3ce��!�a��T�s�:-5�(��؈[��Li��Y��K��u%�b�a�Y`�Ů�ų67P]Q�d�4�IeC\����AB2��R��m`�6�c�1.[lw,�t�eγS[��.��A�,Z,�M��j\K�0V�k��`�nҲ�"�c-�YS"mt�C�6�;�3c���B�ڨA"RjYvs�R�q�0�قU��]��
f�IN
�]v��r<k�M�h<�A��p�V0�,�R�-�h:�.�H�hkU��r�ضa��,�c�3�����-,�1�����08@�S;K�h�D\h�y.X,L.��J�r���c�@�lq�)�a�J�a���լuN1�\B��b��0�Ί�bM@��l��2�5� Њ���5�]k�#H��[--ɭ4��d!eu�h��!�P�����J/֜��R�v���K�2�.r��:�.��n�4��T�
\�f�cd	P�*���ێu����8[�k�4�`�`�ۚV��hY�eY�40CB��Rk3-m��ȼՂ�Tu�f!6�� ��Zeᙢ%w6�Է���j`�W��RiA
�n5Zp�ca��l����l�t[��d�#qk���`؈����v56`K] mBB��5Ix���-�K
H&�w�Yx���Z�!�gU)]k6�D1���5M���YuM+hh͖ٞ��J��2!���!�H:k��Э��p��`�n�$	Ku�t�����Jb�3t��XJ�8 S2�u��Yf0c��к2��a)\jR��,�%���XL���H1թ��]Z8�t������ZCQpi�t֙�*)Ƭ˳��ʹ��p�Se�A�ru�,+
�V2��j�7Y��m61,�3���f&�kI<�!ub�:��s��4cf��Lh�%a��Q�4�a�V��k���-ym4��
+wVX��3�v9�n�2�˗7JDa�qCfR��6a�%iYhBR�:�*�1(��tU4�����G4jBÜ�d��Ōh����`a2uf�s�ͥ�Z�-ݮ%��V�`�],�̷��6#j�\D{A�@54R���4VYW�i��n(�ƶŰ��K���2V�X��f���Wx����mI�p:��Ĭ1��ʰ�cB�=�.�%ޡڭث���h�]4Zd���i�3� �klb&S�JK-�lk���Ba:�d0�#�Z(��a�r�:с���P�R:�8�	)�ՙ���C��1bT,�KraV1�,�Z����/`�!��]q���QN�'v��]H����ur^p%[siv�@lc-X�K�-i�5΂�;.vՆs`�v��Ěm.���g��Q�L��u�n���M�P��QxH%Jp��f񝥅�A#�v�&F�b��t4����V�[������u��Q��Q�\�S&E�酰.�݁�=E�]�f��C��f\�:<��[�v��5�5�飮�uF�@��ˌD3�:�A��!0(f8���x�Ň{��m6+�4�R"$���H��a��ݴ���Wh]kD�hj˔щt����1ɩ��Ơ�t��,`X���j�Z��VԦr�P�<)��l�:Ɨf1��^�
%ҽ���[u8�G*�M�!��Cf�Wu�
�̺��]\��v���K �K,��E�\�Rh$:�vm�b�[�J�t1E6b%A�5��*]l���Hƚ��O�\C9֚�
�˝2��-B�z�ir�5����j֌���ң	qx4�Be�f�cu��`X��;��1���놡6c\�a�%�m�"Qj���p�ѥ5���i4֠CF"�l� �[�#B�X��+L�����¼"�i��m`���+�n�6��f�hʘl�\�؎�m.�%ׁvA���s̰�[�j��3J��Z��l�f�L����s�	��²�ԉS�J��B7Z�zⴤB����4(��]���t��n;g80Mu�cA��:u�{uF9�1��-�63q�SkA���]v!sH�&��f��%��@դٕ�,H�
VZ�U.��!x,�(�V�bi�и��a-"�J�&#���-n5���6�h�ZU�Y��Ӵq�U�M ���u��FkR�.��S5vuZ���mue��=k[ LZpj2�(.��"��v�RR�,��qy�b��i�
FRMpZ͍L�h�X�2
2�n9�܅�3�x���-
�5-aT�6��&��GJ�KfQv�R�X�vR�f̶�R-���5�XX�PU�c��q^j�2j�0oU���ʥ�1N/�Uqy�kcÈ�cĬ�ݪ4��q�雗!t&��I��F$�R��bJ6�\��XE%�,��&�J핔�Ʉ�iepL;F�1��n����f��u!@�<6a��4��L$)`�⪛��sk�jK*���j�H�`SF�%������M@���B�V�8[�P�ۊr���܋4ѕ�-����!v�$�8���q�0t��Y�5���%����-s˸�V ti�j]m��2�Q�+��-g���ј�5KKlf�I���WB��&�7
b�M.ս]��L̅stcͥ�M[��a.���b�4��Q�Ԏ�		�wl%yF�v�.�3��X���K3&ë���V*���Ċ��Wf:�͊���Yr���e��3*������"(��u��ۖݑL�������������������K,c%�2�K%����,�cLE����hƑ�[M1�Di��0�#H��1��iѦ��Di�F��#Li���E�k?>cm��4�n�=���Ye�e�[��3!^�7cCZ9Yr��!�m�g��kg�2����u� �;m���ymllٲm6���YR\Z$��%H��|Y���gOO(ܤ�	+wj��l\*OZy�2�Wֶً<i枱�ՓV�!���>>>:���\]Ԝ�\!��J��Z.�TE�j��K���ª!�M�<[�ff3*l[5�����M��R�(ff+2�f�k6^��=�'�1���ca�x�1y��̫fd�+2X́��Mxt��Ӫ�DV���ZR$
�.Ժ���'1�̉��g0�I��2�v�-U"�[qWՖ�]ȒȂ-kT$DEE"%]��:h�çN�:�%��ϳ������L٬�٩��D��Q)�ir�qvܼ*"TD$J�Z�����i!kZ*\Y���><4x||z|y|g�ɚƼ�Y鞱�i�6�msW)R�����%���nxlчM�:zxy7.�O%�L��u*�%$��*�I���1)p�]:t�8t鿧)R<]�UT�!hHmmKƼ���ix�Dj�eze��F||p����{��T�+k�^m���fl��m[����U\H�V����y)%RI#�D�`C��N	8888'Y��˪�"K��R*�ԥq��%|�<~���8���dq��"�!V����LTY��&ߏ�>m�e�Y��\U�ҫ@5ͨ"\����]fu,�b�2��츄s,��m/#���8Ԣ�;&ip�b�/�m���m(&�j[SY179ڃ��T�,:�m�v.VJ�΃�W\�M3�	,n�L9(U%Chf�)Y�k(1.�0��m���|d�.�3ԱjTaz�1�v�`eb�6T���Pԕc���G��`#I�Q��2�e��2L��6�C�����eQf�^V���h�&VR-N]�MV�mh�0�.f��9l� ���A�Z�m�v2��F�C��Ml�1r�LS&��*1aM��6!�6�����,Y�!�*�[�R���qv#ЕsP+���i��@պ��Ua�ؔf�2�AͭX�Sd^�4ƙ�� 5\*�fi���m)P��9m���q-Pe�mk��f,�	����-�,,�u�ж��*CL!+f�%&�Z;&�%�
�\a�$cv��K�[�u��K i��v ;.�� B-5�)�[H1��ۨ6�Aٚ�fة9@I��6ƚِ�Dʦ5�ƶ��٪�u�*�kv*KV�(� �ۢK�SB�͛a�
�WclF�����ͰB)��`v���K.�=��hMk���9����fͬk�ݮƖ�R�ț
�xF!i��;7s�vK4�ѧ�Vk7U�ȉ�汴���*�`R׭�.W`��]v��e�X֬��
���i��v k�:����5��7lRT�,T,х����Y�A!��T� �����;���[f6�5b�R���E�ª���Ǎ4�oY�"�F*�=�Ɨ�� ���.�I=:t����-Ւ���6��F��K"=m�l[K-cͽF4��1J�j[KhZD�,V�jVV��4h:6ж�,���[���H�T�G���"��T��Ky��`@�m��U��i�,�=F[e-X�� ����
*+Km{���������k��`@�`����_Db.D�P9���7[�j^�.^f�)����a�[E*E���=��˪tSzey��_\-
�1V!8��m�^A�zX���8h��J��bUئ�YP��U�����q��H��u��lj�ft����@Be	��T�`���dc�e�`r�_r�6���%�y�z`�J��pV��I�,_Z@V����ұ/[Tobվ�ו�;�@A^�����M���s�x�1`�$l����c�R�m��z�T-��ie�"B�,�� �_��g���^��lj�f{u�9�٭(�h=�@������,���j;�Z�/��8���bd�[��Y!w�{�c���!�*�V���v�k
L4F��P� H8\mh�l�݋�����|��^��ڙ�gh��r��9�	�UT .���ɐw_(;�_��gWH3Ѝ݃8��EC ��3T</U!�A�3/�z��.��fd��V:96w*'_廾���@�UI��wix+�J|1	�<��zeD�=�Q��!4����Mn��=��:��U��g���nw�`����o��¸c6I��^�<��j��X�8�c��$��,=3��$��Qz7v�U�؅o1�}1M�zڢv��ʰ*�²�ӫL�'"2|J�cif�ι��g}�6U9v�����D^���%*q��r�|-}��ϿW�����ix	��v�ƨ�d�۾�H�˯^��_g�?W�����dkI�=�÷��1������y��qR�<�|<EFG����������!t��v�}q`�g�ck!nE@��c]	�=2����׫�5�
�4 �̜l��Q�8� �0lN+P�j���������{��N��������T�̙��j������c��� c��Z�[-��w��tf��:�������p����ڗ�	�׻���w��oY��*t�hL�f����b���׏���.\<���ϫ)���}���~�x�!\F��4�v�bW��-0�ٻ>��?�U��|�9��y�:�ȭ��3ـ�/�EU/	������T�l��:�&Sf��N�^�]�fCl�{�k87�ٔ�6��sn��{���l�w�^/7�=�G/qF{{M�o�
cqy*MV+�*�����^E�F�z��97�">��t��s�p���^��\Y���8^+� �k�f�k���O�
�4= &��T�m�����RY�J���bgf�E�**�x�K
7��2��h�Q�g�<I��'�@e���������ͤ�2�|�Μ/��kO�պz� �F <MU���zi8��}����,d��׼�͙�{U�y����&M�l��'td2$'�P�����v�#6��;�;�l���M�
�7��P	K�*Y�AP���;sj"�r�� D�2d3����>d����:$ +���Wt�i�moE,�r&�i�ҙ��wMQ��:7*��-N���C@#qT�R��W�a���En�q~�Ĥ��� ���B �+�r��e��֟��5��Z9��Z�w���u�i'O��d�6A ��<m�|�M�kM��k1��m�,�i�/�̶Xm���;W��i�*�;r#4(��X`6�dÛ��ˁ�F�����G�`T͚iL՚����f���C��Yu�x��-h�b��5��[y�#4���	e�M@�͗gi������֖� h��Z���6$�h���* �۔ͻ6I�Ѝ.�h7bYMA���i���ڍl8�amö�e��]�������+U�֐,� 봺7$Hذ�b?@g��
I�~>���_u� -_0�U������Q�NrIZ�ᙲ�5�?�ʘb^K@��K���M:k6�TVg}@]T����;G/)�t0����e�v������Z*ezf7-(��:���)nT��[N���S.�VA1l'lư,u�N����E�����[.�)��dIL4�c�Z�����35�F�}��'���#h��3V�� 5%2�>�`��}-�#łB(ԯ����O���p: \�dV5e��Y��,sh���n�]2ND��ʵ@M�8�^�ݬ{͆م�ym[�pײ�) ���B�zg�hS���d^��Y1A�TE��E�<�
�Un�\d�ֽU�{m��¸Z��rL�lE|�-�盺�Ol+ާs�]�G� yx�+}�w�ޣgom���N�`���gS��x�k�����S8=/��O[UM�!M��苹Y���� ���R��$M�=*PV[8�"&^����k�l6�,�˧�[��OiY׼�{)k��L�J��BdFUA	�.��Yfؽ����mOu�Uh�/?�D>�V�	O���݉_ �!�aH-}x�>��,e�Lb��u���2����%� V8�C9dd!+@��/��Z����sަo�JgA���%Fj�h�B-zg��Tz��f�/g1�䬉�.��ͭz͍�Qyw�N��	�ױ.�qnϚ�j������������O�u���k�}���=&L<5'N���)��p%�2b.Ue��6*Mx���>�݌��
z����}WK�T-�"j��S��HL�&T��;��G���������� �n�������� � ���u@Iy�ʙQ�_N�m"v�M����}��q-�@x�TN<�cSct��!x�������l����P,���,���cpL�ǰ�Te���.�w`3�t��^ɸ���4��p���3����`0��\YW�Ԁ�?u1�B�[zb!z�4��T�Z��uR��^������Q~�d�w��>�&^������ʙ^����PK$��w'"��DDee�\h��q2�2���	��"�6��W�� D�����є��s;P�cRuV��u.��q'��z��̖(��FQz|�86���;�=��3?_O{<���x$���"�k���#�r}��<��,�q�f�A;��n�4���Ӣ��i�}�o���o�{ ����-���o�_V��2ȭY�����&�J�mv
gh����]����ጔ�y����_b��W�n��T��E��蘌����Hӓs#��g���j���������7��H�܊ѯT�o:�T*�l�m��A���A|ɗ*ey62���7�d�1��rrvYLnb�^�BeXQ�am�g-�1M��/�^�蘌��o}p�]�ٌHM�]��M�%�b�g."�\d�V����x�M�����T�&T�k�epX"g7.Rp(;�E����-.�m�����`;l)n�ߑ�G��d�p���<��U�}�0�<��!Fb/�H#X8$+A��і]U�Jڭ���p���q���ZG\���c�&��Z[U�����4X�.M�R���dICGX2ѱm!u�[	����@a,s1��%s!E��Kcj�GZ�#,�b���b͸��iB���B�1^Ġ)���o��pL�[e�](�X��G
���*��r�qn���R�8�e,���	t��G��a���@�]�Ř*�B���=�X��O��q4�vj��E�sf�F��Z�5���4f������[2�eX��-m�I��e1�@vl��&�Z����z�[�"p������H�������n�	������ux��@h�jbv��-�� ��5>�-ʀ�Z��U��T+���5�cq�.� y�)��f� 1�C�V7
}{��{���A��Ѭ^t^�W9�)�&`����A�4a�j z	�T��e��������e��27jV��S���6��2����҅eFxTee�c�l�Y�-f�m���ϟs什|S+�%���>���ȳ���l�+ �� 5b�������C������5�iY��f�3������9ޝ��<��ۻ���Ѥ��{�>��4��=�����9��.�z�+��%�f��z{���y`7�8.�ڰ=`�+΋˙����`�Q�~=��ՠSlһx�����Sn��z��}���ʠB�R),������A�����8�1��"޴E�{C�<�����j�-�4�4n& y%�f���R�<m ��*����僻v�B@�q��şȈ#&)�XB��5 K�Z��PT��qG ��L�LP,��ھ޶L�
Gv�5��N4�]�����M�vo_	 0��q����%V��ةa��m�ލ}�{����-�@ji�a2�̶y�ߛ���{��o��[{�VU*���::𸨆�t�<2*���g�˹j�eZ}�vz7��2g��<�w1z4�Qs}u決�=�>�1�ly�w���^v��C%u�=�K��U����2,~dBG��/G-���[�{�}�fye�_u�=���=K��T��_9/{�1���{s�"����������QO-�f�y{]�:!8]w���#sVg�x{v��������PS�}6�+:�����]3(�ק�Y��{�p�'�Ǥ�ܮ���_{�{�Ҧ�bo�Js$�[Z��+�U��t��<�ӽ�1�U�=JS'�����o�oy���=�a��ћ��E��i����<�n���W�=�s��pt��OA�P�nݽ���;#Ϗ�܏oh�-��M٤c��k�X�t;ψtNA��8����v܃o���j�tE�ힴo��Ǉ�ۚ�9$WN�܄{�����7�ݛ��<z��S�{��W >ѣ�ƽ�)��sB�ox��^�ܳ�^�y������;$�f975k���q�Y���U��TlVJ[o��/#�K9G��}��N���օ΍vVbp�~\�ݜ{3Nc��v�Zw���z̍׆kx�v�ݯyc�W�g5g��<�a=�O�ќ;�k�����G�3�7�N�(�'js3z{��*~�6�ބ����0��b��A\��q����>��ff/w/7>�W�z��*Ҥ���$�J��$���d�"���%q{�ˤ�U�U$IN�4h���㧕M�(�)"�R�H�T��Z��B��t�F͝:t��Sr�5�H��L�hܴII2���Z*TDD�J�0醏�=:yM�wRH�R�erII*��J��R"I.%I"JaӦ�:t��n�I!%J�����O��SR�⤐$Hԥ�JI>>>0������{����$��\H�D"BrRJ\RD��EJA!$�RW��ƍ6|||xܑ7��! �H�DT������R"��\�*���0����ӧ��P�.�I�$8� �$����1	�za����ӧ���*"�f6��6fl���ko4��@�� �rwv�������B�=" �BR H�#f�m�mmf��E5�F>���Fd�U���p��>#����/W��\�f ���G���=u�2_'x����;�jS����+*?���58H��l����}��k�l����\G��R��vK�s|o�A��O��V� �	���
 �T�� AU7�􃏙��cv7o���77�>����"����G����8��=@8Cʗ����[Tki � '��AG���b��Pn�8�l౩��( ɕІY�RX6S��I�G��U�O�]=#���ۧ��K������v��h���hG֧�A�C�Z��ܲ?yo"���b�J�Rb�&�1���Q����ܽ��s{��׿��]���{��R���K0V�ޟõz�n�Ks,Z�D=��尃T���.���R)�9���vqu�7�z��8�`C��E��]���Wk�:C�]�/���|�^`n�5Kͳ���x{�
~"Wx�����4�,[���#���&
m3���9b���F@���{�ܲ$��3K���l�gs��'�u3�}/6�̽�t��Ǵ�v������HIe5 \�p]� �����=��4d��I�}�����g;mw43\��- �%x�2�	�ƌG�6�ܾ4[�s��``�d��gϟJ��k�l�)e�GbY�5���<����n��?	B�Wk�! ��A�<Ʃ��
l��u�9�\�=���;J���9y�!<5oc*k�X��y*���u80C�>����P6~�6���p�\C ��A�5M�M!������^"6�Ņ'	�@]� ��h�.שN�� 4:g��n�l���]� ��L~��gu0Au:��yzl���l]?۴�Gsz�{m�!�R�����pۜǽHq�A���m�V,C!@f�q���UI� �/5ST�vLm�&Ƃ�<u1�ȧ�wDR�x� ���p�BH�Cw�� �ˣ3��&�7����{�|�z�b�+���3�d�Y��>׮4���X�q8qjn��O3�=���yx��R󳿧�A��F I��P>χ�n b
6h������4űli[J�[)t���Z1~�t,��}=���f\K�SW ���2R�]U��`rBl�k���ie�.ָY�c��(�K�6-��Ұ���telj�X��5�L��+�3+JD]bƘ&�=� Ҧ�iV����Yq�b�K0]��G��pƙF:��5��[mePkM��9-S�R�2��u&�D��4UY	%�SqI{�}QfM[Wk�2��ɚٛ�U��Ѭ	�-]�CCƢݷ��S����=|D�E*����+�w%�����w��>���>�y�{�zMb`}4�������x�{�O_�؃�_!����拯�ês�S�E���VÀp�����5�s3���x��{t�-~��9~>3K@�OMU��:���6l�<4E/�*p�q���^�o"h�4��J�`����w0�[���w��1y��V0oT/6�.���-�W���J���~`쨑��	����^A�0PA�R^��U0`jz3�8(��p�`����Z8tVcފ~`L��`���oTެn3C]�(����!�x��_�����E?_�V�k�͹v�ljA-�$��U	��c'%ܗb���G��p>�M� �[�nА�S�۶��ё�p�"נ@�K���HB>9�3|� �7Xdn������;a��<>l���iPy�4J-���0�_gq�c�/�۫(\��:�������o7�櫓�T�LS�r����܎i��`���o�ߙ�=�,��/��Ou*l���\A�0 ���T�E�g�g/9Us�-^{z����eD��`��z��cD�lȿ�*�`��Y�Ϝ��~�����{�2��s�+̩R���%���}�����ܬ�!QC��A��Aݦ���vn�}G������� ��Q�ɘ+�{����4����j�T����v/Z
S
�CzԪ����ie]�� J��o7�R`A5J��q�j=�fP ���F�=Ͼ��?}ٮ�4\;��
Q���Mi�kYA5��fɍk5ws)���Ĺ�m�KYc%=���3����x��Ki���[:�@N��5��������xH ���h�W�)A�
+�ջ�u�}�V�
�	�A��
�i �=�w�|�b�AՊ ���h3�@�`�U3x���.��+IГxx�jw���݁j��z�vI�s�Ԯ��g�����q�r���mѩ	���>�3|���8�~�닩�~(�?���쯩��?|MN]��/�'-1U��||a��x��i��L��7C���ۜ)	���AM��rxwɼy�O�0&�6���[�m{�X���t������+����`Am��v�v�p�Tɉ�
]8���t��y�p���q���b����9[Nlcx0`�M�����hKn�d�LH���`�mv��66�2���Y�o=��5Dz������liG��wq5�w]���x�+C�+ ���x�T��K�R`A}*�פC�Тl8;h1u�xb��;7�:P�oP��@�f@2��5wGf��	���"T���;�L���'��T�������P��u1���%h{\A7h7����"�#�Hsx�� �P`�:֚!<��^0o������J���1�Nbb*�m5�vc��6t3��cO�P��k}����:�zz�׹�n^~����?{<���CL�X��f���i��Fy���擧��!*�$%B.�.y�W����Z����q1� �
�� �7hk��}�&�Ek/�t|'t��C����� aX�� �/8�o6����� - ��2ȟ�C����l��gCe��l�/#L]�֯-�5�Kl)0�p/��|�cT��j�vMU����O�%p�\D �ۓ����А���7h7��A���7�p��Uw��(����#��y<�x3x�˹�ĸNb`A�RX�gm!���n&�� �"���	�"�wk�r��螊7cD��X�&���c@U/5/T��&�#_M����å`#����0���<j�x����5�W�4�<(m�n�`Cm�{"��@�ZB�A��l<�UH�sI��2���	����ʲ�o�. �yns��`A3\.�f--�<Y�3��4:����yN�-'����xl��DB�|vיZ�U,�!l9����a�בfX,�}L�5w+�.��<n'�Fi�x�4���1�DcF-�42QS���t����$;�R�	P�y�"y�d���ėR���KM�K-�����;ZŖ�
����ƪ�e�@&����%:�7U�Zٓ4�a`fh�Z�^R�t��G!����X����Sp�f��Ԕb�b��+1`J�ɭ���tf�B险Fu����u5��6�\�j;ij3$3���픎�J��,~}3&ϰ�Ia,����O߿��e��,���YfmG�˷54�����M�����H�_���6��R��1y�c�sI��:"8�A{6�Ե	�*������� ݩv����Wm��V�e�/i����0퉬�*�x�᰻�Ո1�y��B:G6km��|汳�ӻϋZ����m����������4����d��f�j|���K� � ��o05	���6ސB�T� �����0�\�o��b�oo *��^on�p�:.�`N�A=��ɝŃ�( �~of/5��לݐ��1���EM�Ź��\(g��&1݁�zEl_1��^�kb�� ��6*?r�A�� C��O~��<�^M�!�,̳��W!\J˜�-�@�B2��aO|i������� *������	���J{"���.^�S��G/T���鼀o-������ń���}R�h6ޝ��ٖ�8̨l�!�^HzO=4����{�
�^����=�]LJ2ד�fRMCIe�dRl��Ԟ�W�._�Z\�u~�����*���xyX��xhcS^�a�Z�G���5}6ǰ��w��D����[��*+�^��߼�S�>���L}:�©�Ʃ1�!�)Jr��%�/s����HȻ�3�i6�x�/ުB�"B��`����BH�A���`���^k'��}�qަ\^�x~��_|ϵ<�O�G� ��A3HLƩjs�ʃ����Y�ճ{,�A�}�F��4A����h ����R��%�j��'���y�E�������iK���i�:P�u89���1b�Ĥ�$йp �:��W7����	S&���x�Զ.��p�\D`��4"�P�k��`� �퀻�Ѣ�u�iu�<�e� j�5�[Fn�;U�
��Ľ�7��#�U)a���!�9/=-�yi=�׾c�ɑQ�d �6����K%�Zg&�;�G'Z0�{��� �������ܽ��7��aiIk��=��R��3i���������{�����)���Z�BJ!(L���y�ڝ�����Ϛ���F�U�iQ5����v�����r�>��8<��!��^cv���9�b�jo��5���Љv(��w�QӇ��B0�d0��9�W�$T��{ڐhsMSZ�ڭ�Vm����7�'5{�K����r�L��t>�0S^ҹ?�dM� HG��t\�WJ!.lx�i�ql� ��Sx��~�>�e!>��$4"�y��05�[Oc�u��a��aU�Hf��{�,���>�؏~�rٵ��^x��5#����zyz<|&�cfVmj���v���<�/`ER�ل��|4'��=��G�}u����u��fD\��Z۹��ꛅf�]������ �T��9�;������d�;�pC 7h_��^����v��tM!�"�1͢�mz2�Y��?b�c�<����x��w�uS���\�^��ݛf�C\af���O����:���l^����f1%*�ĪBU�!��j���^M����O�x��0���v��hA�J\N�e�a�� H3��5n���Ӊ�u��� j�8!v��vë�^"�/1�Fn:���������C�E��]y�]t�0��r�" YdD�N�l*/�F��?��^l�ES7�5H0�76��;mR�9֗�b�89=�� ���S	�L���T�OTx6Q7�Ha�M��0����MFI�}gD����u��U]�h���dxo��r�KbNA��ޤ�T�� ݢ�r-St�z�#'bw�=�.�`8%�1�

�1I���
@`��]V2��������!�|n�oL��T/]D��9֗V!�y��7\D�����3+�joU7�R��`*���6�P��w6h��)�YM�m�H�LA����Ȼf�	�����8��d�ĕ��?[�Rr*m�)�š.8]�Te'��/ U��n9ݦ>�����f�<흭a�S�2�jd����3�ԓ�-+s<��y�z�q��8gu{F��ؑ:p�>����b�aŞ+Od�w�9�OzY��o#8U{�F��g2`[�n�zVj���<C���EѤf���2S���Vp��[�y�J/b������a4�}�f�"Mw�O�ۑ�0U�<_�����D�5���+��5Lm{�s�ϱ�gp�$�o[>a����gb�v����mB	��=r��:���Ľe�ٳ���}
�0���-\4����,��P����ۜ&��/����̓����{��{�s�����Ӑ�ʍc��M���js�����ťбטow��w�A����K��D%޷�WWbN�ԙ#n�0�a�u8󞌥I[�nכ�E�b�e�O�!�эvh��D��\���؟��P�v%�������Y�N���|z�YSȰ���vf>'�C���x�k�
��s�g==d�����kݦC�P�P���Ңt�p���+���~��u�W��W6꽋÷�����D�>K�j��m���̾�{�S��oeuڢ����s�XO��ۍE�HUv�}�1踾��>���vSJ8�pB ��h�s���}�M5���>�y>�6�Kr�#�P�,E�EI1�>"}�\�hl@؄Ҥg~aM"cO4�N"U�YՍx���3W0����#���4���~o�:1�C�1'���� ��/�H)���os������Ƒ4ŋch�F��Z1dZ�if��0���#L1�cOQ�#Ki-Y��#[�ֈ���1Z#F-�<i�-lx��4$��Y�l5��
��F��4%��খ�M�&&k&v�"Ȁ3A<�<E<y"f9��R~�� ���� �ԁ�8! !��B�8 HG��0��Çǚ��D�J���cF�֙�e�l��ͳl��z8�>8��:�5�8"0�0 �^N!'Ӥa*H�I�Θxl�ӧ�#<��H��H�p@�FH���D�"��i*I>,����g�ǜ�*n.�w*T�I%IU"[f�[[M�ͭ�Ƴm�k�'�=0������ڔ�TEn[3[Vֲ�|��Ͷٍ���UV0��!�8t���IP��"���H��H��"I%$��B$I$�*"zC�OON>�NMK��RW-i�k�$�ٶl��o5�f�66�6�Ą�'Ht�gM�:y\����� t;�|!{�@�cm��ٖ���ٛY�ͷw� B�+�B! 	� >� 8$N��=5�j��z�+e��Kn8a8�h:����mZ;M�ʘr(��6��U��G3��	�����-�l+�2�qx�T昗d��&����&�$,�C�gL@�Z:«�sZR�Ɠ\�-�B���5�u��e�D����&WM&������b�X◂�JXg$,Щ�s0�{�ݴ�	LT�h�2�hW:Sk�6��U�A�0iIfV�fA�[qSXKI���k�!����Fzb�Y-�`��������X��&�ݵ�{,���X�l`P��e��3����Ah��d�\X�GJ�cd4L�ZE��,e��R�F���]fqJ2 @��;��ųM�i�Z��rʄ���XbaB�ۍ)�)�(\�R�Y�.�B�	��a0�8e���Z�:mlԄ
��
�c�&�!����O�n�"2��\��j7J<�٠�U5�@p� �3t����.Z\��E#.�	�;Si�4Иf���6Ck���9�uХ!��ܬ+Pn[f֚��lR�fb�1�s��ƴ Z�jD�6.����*�mR��,�C%�Ri����Lvm��,�)���r7vִ�ʡp�c�͑mն�vכA�4�
':U����"m3��]\�4��`�å�ؕU�2�A47%�6�Ss(��"Z���k�ɒ:im���Ikt;6���-y��B�`h��6�R1�n�g-*R�x"䘷Y�M1k)XЊ�L�nte�.�:h�]L&�2Ц���6�Z(
��B�;mb��6����k��+Arb��7�o[���6�2h8M[ND���t0�Z���©�͆"�u�ɊC�����6��cXU�s��L��+�-X�p���UUUWK	�FXBXBXB�a&�3\ˍ�W�fd?�HH�"$����\��$�Qr�ˢ�!d�T�Qs�&VYt�%�$��yk�`;����v^M�m���oK[]4V㉳� 8s�^j:�j�qv,e#�s4cZ"0,��&�9-�Q���,�li� ��������T��L�[���c�V�ED�3qc��b�idLc醲�m���12��ƥ�d�F�V������&��#Q�c��ks2�6�k�^�1��	�I'����i���.*h��6�Jf��D-Ka0�Se)S<�����|��Ob���R����������f��M�a�>j�gϲ��c#��D�1��%U0$za1���rS���F����#.h5�(�':��	�^`{W��gU���@�Zi{�� �0`ER`5L'0֧�@W����=���������@�d�x��P�U&����AE��=B���x@� ��& ��T�[��G6�W\'��M�@�z��h�����0��Y���p]��=��	�ڱ�OI/�����+���6���X���gh��x�D�!�5I��R�y*���#�0ZFh�BO=YO�������e�]�db��n�b�����X� �6�� �D��y�F��'1<fcF����ڑV:&s�M�����x��5�z /�i��K�@#I�������n�3ҞbU�jS���3,8��Ys�`���+��.�����	�}5��c��hw�3��3��վ��m�x�^��,h��̯V2�}��G�cI���  �<���M�����6_9�>��Y�mq��^�q�
f!7�k�H�`�+�lBH1LƩ���l�*���뽻�q1�i{�Z�v�����5���ڢ6h^�:+�r2� ��wPb��յ�>�Vth�X�ᔃ3wd���i��A[�����A��� ���ug1m��7�Լ)Ds��m��3�8N&Z�a��pn�on��MA�r�|��;M	f��F����ߘ���3��l6��L�ࣲ��4�`�2�K�[n��[���X��k!T��4D�{�t���af�\%�N�3���G~��n������ޢ� A�@�Z��:�#�״ɢ����eH������Y�Ah���1G�Nn�]��h�+VC �PD�߷��]{~�'��DO}�u�s�0�ԯ��d`� ō���J���&yXL/NY��y����
~#b���7y�q����ʷ�ԣ��V�U���^&1=i<4�iLAHJ�.R�J��;Ϸ�_߿���=�,��C�A_ �q����Z���Q�	K����W�y6A�a�8C-�x�Ր¤?b�w��Iw�j�;��1�%�|'�x� �A5j�"��^�`0�oQ�\nl�T<6X7��H�¸u��X�x6X���*��R�	�Aܴ2͛�k
xQ �H�E��'�D��)>M�y�@���af,����i�J�q'e�O�3W�|��X ���l]���q3S�.W�'D�;fMDv���_�?}��-�'9�#��T�,�=��A��f�K[�!��c:�;Ԗ�^�(=Y����m\��[w"�x8��V�1�A�ER|*�b�`Ɍz��G�6���84_\����� ���	�o@�O��fB����x���`C j��l��n�狪���n�A�A�Q5����5gf���iF�!X���U�Fhb�*�"҇'��#,���9O]�����ý�ʟcEcU1��	�X�X�XҬiO���eU�o���+�m^,�9�$���G9��[a���i�ֆ��VCT���_$�֖v%����3�Ɂd���8l���wV����� bCnc>�^���4�{L�7j]�s7Z:c����ډm �r�x�ڽ��lѢ��T��k&E�}�&�N��S��xE�i�{��A�sy��k7��y{l���k��o��Tᷞ��5�� �ի���y������11Ƶ �)� d���ܗ1�{�4���!x���!��1+�(! *���m[��H���6��! X�C�y0
e9��dX�f�ׯz��@ ��1�S��8���{%p���n �p�D=��5�����Gj����{�eF�������� 	�����\����/0�s�s���踛ɾx��A�*����Y��ʺc�HF��Y�a�;�H9E�.휣%�oq�"Jgxsu�#/�O�p����n�	a���av}�8ot�|�6cH�a�Fpn
4��q}�m4ţm"0�EF#KB�5�$��%��ӧ}䲘���cDc*���JVT�B������O{f���rbRVX���a�JMe�Y�&��Z�Yj�	���J�.%b\j�!�6P�
P7Z%f��PѴ��-l#�%K�RR�
i[R-3�MPK�43�V��SpA,�J<�<i0Lm��8bHT��o\,6
2�ͩMo�2�-[�j�:f��u5�]�;2�3t�B,�y����������6��\���[5���͑�fk4p�RY�)3�ř��H� !��1+�+�q[��d��k4v�bA�ΰ��iJ�A���pA�P_��5��4#�>W�$����C������V�c����n�Y-�/�d/x���L�U��H����/��r�����L&eH9b��9Ӓ=�1�9�a�s&�Y��Ϭ���dܫM�ޞH�.��<�֘�D�`�#�L�W��n�`M�����H0�bbt�k�n�L=�� j���u1P>�A��A��1h���^n`�{���^��b�ڎ�Y-�-p��H6X�t� ��}��"ƹ�gK@�D�@p��)��m�!��4ÐXa�X^��3mY��`֘5�Ԛ�[8��<������c:����p`�2����#K�VVE��E�x,�ِ����C�T0�
��G�]9�c�jT���Oe�F��/I�Y�J�4��1��b��(D�2��ESއ�ox���y���{��[k�;f��X�Kj�6!���Q�`�K�����h�5�cP�������XԏX<1%�·�\���א���l����v$=�;���
�:99����L3H>,ʕ��D��qi�R��/I�����>��=��~�L��\��x�oYt��	fo@L� ��cjC޿y�7�|��LA�M��w�ܹVVE���`	V��^�����x�:��`}x��ES>4B �
�`&_'9��߅b��z�j,�Ǖ��K� ���^Fe0#�̪7D�̘��@��]�1`.c4��2��n!�����ƙ#��͋�FZ;ﰓd��ax����w�%���]�\=���鮍���� �E��� 9��a� �K�}>���U/CmYy�j� g��07+�fSw�{��ew97�����2> o�Ԏ�DR}��#u +Xk���P
���}\�����a
XHry�+i.�:mk��k����5�1�>�������;=j���ќ�,ս��O��j������_�JW�(UB%1�1��U�cE1(�J�Y)C�T�'�{��5���w�w�=���S��"{f�zD���:-Ɉ���}⛋�}o���i�/�M�����4��q�N�`� K��٩��� �����>>*��<MRb/#2�߳[��XR]���r 0mi���m��s�}�=��������$'x�޻���}K��jMkx�4�����?}{����Q�6��D&�]�4]�,+e�[ufД$��bth ���?�<��� ��g �)y5@�㈳��V�֗:�]�ެ���Z�)6 �5I� �>�A��V��q���xE�o!c��o��:�_A�ї��8By�� ��-��Z8�o3����}��� <u{�=�h[8 �x���M�j�5K\1Q�cR�{���m��������g�߶ʉ�q�7*�ox�oxa�f��m&YMl@g�F�7�����sK�oJ��ĸ�ux�����S)jxsO��Q�"s�md�9�LL�.��ky��a���=!�O���r�n�K�do/�����v��1~�?{�{� @ N��^�$cc*�h�A�$c%�������{i7�(��R`=�AH1����5#���{�1ތ�*�ikv}k�G��whŷ����O1���_i[�D%I�=O?!KD��6�0���[�s�u�]��T����nP�e��L���d_ mO��h]�Q1���G���a�Dv��
l��ȟ��z���[�з9�J��y^jU��6�nP�.٤	�Q'�ޛf�Ć�F��my�T�7z�a���}�"diD���~�-d�$1(V�^l�Z ==L�"Ʒvo����=��^��eM�\��Q���+/��0��)�zew��͢�q��0� �����V����ȴF��{�7�M������VD���=� |��Uf�V��٬h�ĸ ������@̯1�Z�+����=�b�b�0�X��(��qm��v�#aT,VS��x�y}���5h�2)�S6{%����#|L��'�u�!9 K�$S<����P�-Z��-]n�y�mvxĴ�B�x�ű�M	�%���Б�Fl뵌�������	�5TcO�xd�5Jƕ<�<1U���d�(fO<b����խy�^#r�\V\`��0;V��R��px+u����&ɬ-�쎕b��Á���U��R��p	�8���v՚�5(����0D�af���*]��`j�-���53��(@�m�I�
\+�t*�%t�3]5����!4%Ѵ*X2�Z6%"�9Ud�2��[�j1��lm��l���#l_���>��e+yp� cb5Ѷ�fD�q�L�%m�5��j�{?��b+o! ��c;���ѭ�݅�E�y�y3:^�i�� ܀ޓ��%U�I�LDսt"������:���j���Q�%��8a��`"�4F�ZU���3��0�8B�5H9K�)zXG4m�_��|s�A��V4��n�%{��J�����D��:Z�=NBR�Ų�x={H{c�`A�oqA�`�o��ld67v�}�
6@4b;m�(����eT{u��R���J�y�g �+�t�	�hv�r5U�t4n�*~Ü0�
� �����ñ���;[�C�#�G����Lˁ���Ϭڢ������:��֑ڶT�2�y��S.p�P���M/y�/@���, Z�j�5���WMe>u���`*�8��l�i1��צ\UW9�9��G%m��[���C��BNհN��+�q>���L�X�O�u�d�Y!����X�MC6�ى�zּ��8�z��=� ��{�/$c"1�&2��L�HcH1�<������@	��`�2���k^1��ﰧ�u�oYr�2��S�� W���D���X�G�ڧ��Ѽ�_o^�<>qe]��a�5k�q��s �A�ES�[�1b�	�@37��f���S27�V�)jʜ�K�k�oN= ��P�� <� �6��(A�A��A����B�l�3��u�@5�fj6n��_�aQ��6B ��b&X7��d�܎�3/��${�B3���}�it�p[��6�XJF81VhFݐ�]��F�8�����}�?xi~"y��H �o5��sCG��1w�����m����b�g�(M�A�ql��$̱ڣ ����l�7���H�c�й�1�),� Fs� bE�/���ɠ�������Jp��51��$9Sp}�� {�����t&;����}OP������Ro�@����F�ˇ^���/�ĜC9o�F�H��n�p�+3���N����玎�c:�Z0��>�"�\;�s�x)YrQ%���D?vO��Ú�")|�=�v
��,��ف�^�tA�H���,�F���{O�=-~9xe����v`�>	gu�m���a94o�׭���u���˩�h��m������/R4��{�ǻzg�%ٸ��in�w�s}�X	�;��f�0��{V^{���7��Õ��N�&�#Ƥw��VM�s�F�Z�p��F���;��a��V�}���~���pt�J�[/}��M�=�7ۏ	�}�>������^�I�L��,\=�K�u,��q���aN�[f�e2u��]��&��A��Լ�8��,��/jo��,>X,�¥�VY��Pb���A�B����l+=~�{�s|��6x��P�k#n����v{mͼ�z��/����xay}���gP��O��ZB[��tzT��[.�
�à��3(���^~�}'�[W��.ξ��2�y���}��7�$_�O���|r�H�!v����riW�2V��s�]�DW����ܩ��:�I��|#l���CG���`��I{���=;ǯ�hy�sQ�h�F�{zzN�{�:�=��T���$}���\y�$b+#�g�y$dH<��^�LՓVd5���3�$H$H�$	ܬ	l��Ċ��IV@���2$y���c�Ȳ������3W 	�X��N��3n���#�����"�ֽZ��K�|������Q��� �D O\! �H~�D�ܵ�D��&K�">,����gN��I$��)$"I*T�"D�"ST���Xʸ�&B�	ih��K,���Ç���R$M_�e8!1�!�qBC���w2Z$�*%J����:p�Ӓ|�Ϣ��Y���  �q�2� � +��G�t��4l�ç�T��I$"&]���"e��{�%ED"H��DI$��e�>>=>7\�D !*�C�F �x��IRD�+r���$�zl���{��OG8�t8��yb�! 8=(�y��q�~�8��,�����ӍNJ���d� C��0�	��q<��R�2�qmYӧ�ON��� !��������  6lƦ͛[M�my�}^�>� �
�@���zǚ�m���ɥ/��V5JƔ��V5RƉcEL��TY(�������������}�����p�G�5LT7��� 2� ���o�%�]bb��b�A�K����p���1h����W	�W����+U��2����X[���p���{�ݛ���� �>U�c�s�q�S��Iw�<A5��T D �]0>�H>�]��D��^�B��q�$ɚ~�����ZK���#�1�t�].�qP�!5j�µ4{��q}A�1���(�&X1��5��+:x[>��-ޮ�y�M�>L��A�f�2B@)��83+�O<ζS�#Lbi@[S��,�Ѿ���^�NF�!����ـ�y��T���C��E��u��hC�s�ǉ�ʈ��?����i��Τ���� �2E���1>�L2H>-�t6���y�q���(0"�"��Ppc0vVD�v�w��`,��g�:��S��4ƙʗh{G�����=4����f��b�k� ��ی���uqo���F���m�Ȧ<^o����^-�J�P?�
����UT�"�U1��ĘԖ%*���?��_wuY?E���-	�.�EX�!u1����8(8���+���h�����n7 \�Ϛ��n�+�2
pC��ɽ�>Ϛfuv�Km�ե�Y�ni�Z;�5Vx(:5� �D x�!���Olr�Q��iy]i׭�ݺ�WN4�W�
~�H���Q)7�� �*�r�v�Ʀ�WZb4�lFE�cpe���N����x�(�2�=\���{� B5i��W�>�� D�W�1�Q ����1w�����i 6Ӏ`�Qc_�����;'�G��]Q�߽I�F��§�����������=�1�.�k��mTvb<|]��i׏��J��e#�L�s��7�Q��1��[�ѝ;\"Dg0 �(�*XX�f��q�'���K&�*��M����4m��o��U�xTiޕ�/USN�YW�1O���[�pf��+`�X�`�ƻ;��0:巫�h�"!�Z1�iX�#
-����?��I�!:w2�5��ZOF���Y)T�y��ܼ�l��\���@ħ4ky�[SL�72�7��1��5�DeɢX:��qLM[������b��d�c`
v+-ج�fX�cj2ɥm�]q���.E�6�Bj�X���NB6X��rl�f��h���b4(�4Ks3j0��e�ic&�V� ��4Tns�ܰ����),�n�_S���lcI���a�[Ļ�Ĳ��L���ر�rXF(�{�W����j ^����Ro*��t������w� �9ϩ�k�z�i؎��G�oŹ�i�ԩ�f���KM���oj��X���TNE���n~��WT�gZ\�br�^5I�p6Y�������B� ��<B�%�F�����5�Gt���}���#�u9�Y�oxʕ7�"	i�Cj�[�8�icgш2�VN�n�J�*�o��� �b���nj�RѾ|y+o��{�D���1��ʉ�Pɡ�-�#�&���;x'���Τ���p@#����&x�̯
ٳJ��Ƴȱ#X����D��Yc�K$��� @.,m���&c�橭��L-]���~�d������"JL��w,s����!��<��7^���mP!� +��! h
�s�����tj/F�d���n[�{�(�}>RpB:���v��ϏOAG��5����va[�y.\��=���|���߹�*�V�O"�ʥE���T�&0�d,�U�QUd��&G�痑'������+8�k�w��@ ���f�1XfLf=�����7 ���Q��*���d�Ms�]���GDI�rj��:��x�A��L�S�!���ٺWe.#�A��b-���kB�Ű�1k!ka�b��f,�Cխж"�ū1Ǟ1v�m��m}���n'38��`E�,x�2���o4;���C}�Fy�i�2(��<Be0��[��1!�Md�����^���Y���ƥ|7��x(1i�����m��|B �0A�	,ͽcw-�:�&�-��e��a8���obR/�f�S�=��a s�̆H@C�P��z9��/:��A�b�g<����!���fW�i�����h�niuN�ƹի@.B(�A)���p��s[x;�z+��i@�T����;4g+u��,��Rb	�L�!j`���o������gT�s'�|xP��a˽ޣQ�%SXV�)�_nM��v��u�;Q��n�[~qe��x�����-{�o��Q�R��QV2�Ji၍C� ����[t��c|;�C��A��A�W�$<j�`ES0�h�̆շ^�:d��=d!DuP���9��/:�p�x���&�-tC����b��0�kx��T/z� �L%��
�c`3,*,�n�zݸ�}6�Dp ���x���0�遏2�>��I �����=t��i�����fh8b�6HŰsY�̺Ĕ��>|M (O�Ɲ7� ���O�d����7Å;���^��� �!�����\{�ߢT٧s�$�'�{1Z�|b�`"! ��}3�0���t�y��x�j׬���]8�h���0!� ��#�kB"�:���~yCsgƆ�ep`6��v���`�$
>Fe1�����+�yϻ�0fU����c�-���G�pj����z&O�Pڈ�r���1"e����b@R	���Lk6�U6�n��H��&�9�W�������}�f���wP�Ϋ1�Ī!*�	G�Y �Ko*��cP�ޞ�|g����3D��%O�;�vr.#��Lɇ��g��M$_�2���U��z~�j��.x�ͦ �א3)��%^ԉnx���-cF13ߏ/�RZ�q�If�\Ma��	uV5�]6��vں�W�;��x�oL�C�|��D���w���q��Ӕi=dג7Q^���y���վ/���ݯk�e[n��F�|��0.@�*�KGY���m���G��C�=0c$H׎�Su�C0i�  *�0L�x�^Re�LcG;�y�k�[2����:��	�LA��^�2�%�A���qjz�r�hp�A�`�*o��?F��n�z��!�qD\Џ;��<A���Ԁ"�_/����{\ֹ��21�n��Yn���<H �~A�
�p�"�U�w��3{Y�35�L¤���0nqP�;C[z̝���������rzns&M�'��K%ʲk;���/����\��ɚ9k3��{y"�DU���h�Y��XM	4%
&���Ry�'��ƣ=jxb�F"��\,�T�'�.�.oV�Y����Kh��:i��4��&��-ٌ]�6!�4�9���Yc1c�SKv�3v�B��ll%�k*ʔ2�(�h��b�P��e�\fgl-HX*�`�8�d�f��!-�]��ء[��4���wb;$�Хf��5)@�`1n��bi�fgD��k���yKŮn�������o�%5�6���[���Hb��ͨ��#ao��V�]���y��!x�|�`�L�I��ff��m��n�q��hP���r��"���@AL�2||P� ���'Z��04Q�vP���ׄ��r��Eo�!�������(�7�9|��`6�����l>a�T���V��&�Vn�	2+����G�sPa�=T�xɀ �v@U!��a;�W��
Tp�37��A3=�sl�sS�mpx�jS�u�,Wq�Y�B�L�� G��T	8�oQ1� �`���O��{?{w�h�A�`�L�x�^=;ñ��d��������3����jϠd�`�G%�kv����9T͆�9�N���t.��Wu& ���3)�2�]��#�vv�ۇ	>febZӨ��Z�*�� ��=�m p�BQ�{/��\��
�����opE~�e;�����Q��㼬�`��z^эy�	���r�EN;�oN3��)�e������1�X�5�1��ᩌ.v*Q ����fo��O�-UNu��r���1{��ew�op`fE���A�C��OBA�`�H@�&X3t�l�5�a�WD5�Y������AAL�7��H��ܻ��g�{�L���Hm 8@�,��'�=9mm�G��#�K������� E�L�d�G��X7����ղy����Z���ct������� �-{�4�L�~;�V�p'\�`B�)��rX����c��5�xrT���\�s����\��?h{;��2���"��T0ۛÐѯ�td>�@��py �͛�&&M�����@e�8��! *I�Ħ"v;E�[
�#���f��͝GD��۷`@���T �H�z����t<�l���>!j�[���ݝ��{�X�i��v�x�&ퟪ,lMRR��k�Y�~n�I����L�{s�������������������?�**���HC�׆Xь��5X�ƽ��G��|���e�[��A7	�����UK�j�tB�w޴�����@�`��L��
��{ѫ��w������N�׻;%�>#9���,� ���������W�
^l�}7i�uf]&7fٸw��-�{)�x�>R%�i�ۑڧ�h�yψA��if��.�=����<k��0!�9�bk�j�B%�0ERX�I��P�������c�O���Y���SY�y�:���ֵ�Z�%�`i|���|�y��L�c�!��s��n�\� �+ŀ(U�l�7}��˕�w�y�"K@����0kfo�����_#�L|~�`0����NU��6�\�f	���qn�8I� H�`��s$	t'�/��	�YKA��"H�@FǛޓ�"fv��F��i̤p�f�����G0��1#�����w:?Yh���H�u^������_�ߣkzN0o����.}ߝ��9v�η�G��>Ƭcc�k�7u�𹻬�����|cّ'��DV������(*6I�!�o}8+>��Ϥ�u�oy�D�2�'�"�ߕIAN���~��?,��%�7Y����v�*@ia*۳1�&�e�5�I�y��=?8�>^���N&e7��΋�/��	>7ϫF;G3-�ڰ>H^#��L�U8`�H@����`���")�{@�暪���֭�2��q� :@Jk.2��j#�^p�_���`*�h���	:30r����@�b�n�$��O��Y�xK����c�f"J��x�<T��Y�oi����B�17�&e6��Q��fٸp��� �!5�����_t�~p���q�$"-A�3s�Sr�wgDw�bou�^�ݗ�zi̾�\%�01{ eT���~!���e�}�6�ʘO�*52���
�,H�A�Ռx�A9��.��¨��e�\ʽ�Vl��� ���6����ţJ��}�������+g�ɝ��Y�^��o��>�����b�ocӂtڮ7��w����Yޚ���H���mQ���x�_s��>�ݗ��!;�xo���χ���1��
nm�^lD޾�[���M��;7�2�H$��_X��3��W;�S���f�@��^����,������.�����`��Qx3O�>{K��O�c��~��ks�M��y���<W�v6���}���WVzxY��}�ǖ+��t��]�eF�R��Eq�}x.��+H����mǊ]��t�'�������#�M�{o���=A��=�OO18U�_�ޢWR�9���Ö�^���^e�3��d�7Z�[ͪ�����RgU�K:2慄�\{�3'�n�9y�U�{�7�������{���=������$f��'��5�7�Ǌ��n:�b�\u^���g̅�Ͻ��	l���Y7X���(q��w����Z�P֦zx�{�
n���J����v�Y���5+p$�ut��:h�{��g��h�:�&bמ�*s�}�:��e�=��z��ٞ���S ���=��on�1�r鐕x[�7�8!�nE���1�W��@��[�L�l�F�3D��BLcT�&�bB3P���C�����0��_���t��Ѱbad�Lc0qƪ.-�WR�Hͭ�/G��U�]z>��۴�4'���d���icf����<���z��[�idi����[i����F��[E�-�4�4ūX��Dab4�EZض��L[ű�ű�-kZ,�F0�1��kh��yyZ3^f��Xkp��ټ��Rв[ũ�ff�=��J)Q��vΪ���4+'�	 ���Y�m���m�w�o�o+5��D}�f:p�æ��&$J��bՀ���P��� q<�"9j��>:t���)<�\�I)$�2����JBUHFKt�\�H��:t��ӧ+���	�'�� ��$ � ��R�%I%T�!f:t����	�  ��$� ���!$ �"I	(�==8p�ߨ#�$N� V@��H�E�LJT�BHIN���M�8t�q9��MI
C�8� B��<�#�,�Ӧ�8rD���I%Pt�㽑� $@��˕$�&Y������%Άy���e�31�2�l��5f���+������iIIZ������ڶٛi��m���<=��J���v��`�Ue���IvsQWcl[��3VcK32�iaI\.4�R�q�&�,ɻ7U��ˮ#]��M&�bB�B�-ui�K�]U·Z�0[aq��%�5�g&.M5ee���6S�Z�.iIFj�&6����[D��I���G[ZQ"��Q�� ��Z��sl���T�"��llF���ĦX�.Ks�\�ƩKQ3ii���6������.˶Դ�1�1��.aQ#�#e���Ҷ�1m6� .�Xe���(����m#5�3)�D��#��*��"��&eYJb�r�a�[�p�1�)pE���f�]e#��RR���hn8,�5٢E�-�F%ګbd�e�Xj"K�\Ҏ�h��ŇL����9��"�F0�ju�\LK�J�+-��"c,�����0���[)Y��'
k��� �(�Q�v�c�	XD��>��oV�R5�y�
�]l��5�е���0
:쐨E���i���U��Da,i��u"*�h��CF̩s����SL�f�P�i�]R;�6��p��E�0vWhT�W"]��u4jhb���΅
���1���3Z�a(���ɵK2������(M��ne-,1\�Li��4!*�����ts�弎
��Sa��W���v��jbf:��Ztb���o%7%f���RˎuF�]]N�$bP�����ݨRnPq�Ɔٚ^��ˌ0��D��LM�Ul��Ո��5�Z����mJr2:l�l�RS	�sv��������m�b��vS�e��媗T&WnԹڄeġ�K����@����f�ְ�,�	P�]V\��v̻h5 p-̣6i���a3�+��J�UQTUUUU�K,�MI��ddaMJ���֤L���N�u��2��E�!��D��D�����+2�"�Fk�+���Y@lqɃc�������4vL!a2��ˑu�-�3^՗;�#�Z�U�ë�+v7j(P�x��e��i�V��RXap�+��8лBĖXg ֻ-�e ]5Gi����!GP,p��ښL��b̃a�l�˪��D�3u�i4X������m&�fԽ�a#ؔ.,�)l��Y]U�.����#���z�{�&�|��v���uOA��=�ސ_mp|���T%��x�ܫ���"T��6[�ks�U͍�*N}t�n��{lG�m��A�	�A�e0c$gOF��xc��ކ�/fX7��f����npѯ������;vb�+/�x�x�� ��1)�A3)�����C�t�8f&ؽ۴=��p�>,�5�N�Aj�=����!=�r�����$=�B>���� ���C��e�R��d3jk�2z�
�7�z�[fݸp���r9M� �a6�k�1j���[0 �������v�k�5�l��kmL����A�)b��Wm�y��te�o=0K��^������9{���z��eT;פ�/���S{�O�{6�Ww��=�l���o�<æ�T�Qyڋ��Ϫ�)�u�t�b+"��������wc2e���0��kM���,�G���DIe�r���U]������y�亮�J�����d A,<�L�[m*�S�E��c�$�NA9��"O�t� (�%ꨋ;��6
֩�X��5����7�ׄ���&������0)�h��`����@!�yD�V�q�k�˜�\���[Vd9� �*�Փ�^"'۽�&�*ov���o*H���/&��`��]�ʷ%��.�]���l��K2�W�[�c�;��YdD��g�m��颵�R�d�+s��B�
�p�&q��u�3	|N�'�=���H�2Y��5	�>5I�,�����Ä #�?G�O��Ρ�V���A�a��5H00B�Ցn�gR�'�3�Yzx��E��R�	�^�@L�W	�5�H@Z�M��PA�䙼 Y�1�0 �7��2�N�cK�C��v���9+���}r�;�<c]N�*ڝzL�2w./1��H���!B��0Az��|��X��ѹ���:�#� ���D@�*��e���Ӌ���oY�� ���>���UJH�-���g���$��Ǳ7�&e7@9�CS�J���� �sp�Yqי �8B#7� �ˆ���D��ڊXX>�8�^X��׌{�E�^gL���p�@�,�L՝�5��c��#<`� J`�����e>䭖b1�棪�n��+*8.5�*�l6l�Du��O��e0b$�L�ܷe}���Z7�/��@4�A�뎅�$�9�7��o7����� C�Rr0y��*f��� :@9�6[�h�G |z����N��:�9׊�B�n*OM9����~��y7��K�ъ�zf�}�9�2�l&�#2� �j�h޶C:"�\5C_pw ���8�����ey�����8e� �#
#��ю����g��c#���l}���E�h�1���fq�ySy����7����s�{Tf����2&�����30x�Ç��� D$$<���x<���RE�� -v��n�|l�ʛ{o��� ��7��Us{��4sJ�ގA�K�� �1YQ�h���܏[oN���-,����>��j/&a��u�l��G���J,f��mb�a|{@�W����Q�1�S��4B]{Y��z��R�[r��px�|]��L� �,���-�73�X������C7f�7��=�� aD4�
��]�Gj3��d!`)�� ���C��8 B�Ko�8�X;=��n&��iZ;�@�=h0e $��X3 �������5}�YucC�8�`��L�o$FU����c�=�l\���	�M!Q������L'u0����L��G���1z�>՞�y�6���k�k�>����~Ge�ox�-��*�n1[��8�=2�T�A�O2ư���[��f"j�_]F��UxH�Z^B��M4���N���_n^^_B�nԏ?�3٭k8^[u�m6�lb-k[�f�9u]^�I�I@���'�˦�)Q�X͜m�t�V�.%k��d�2%�n�HE��4Gq��D�.���ɲ�i��ʍ���K�ciu�"�c^Ѯ�`�0)�]N��]s.!��b-�:7bSS<h�B6�#D�]�eĳF���]lh����m��,v�]0n������{n�Mٳ���:���]@��������C�f�e�2��Z�̳\m��lt�b͡��!d�-�J���@i�L�0/)��Nv&֍��ގ?tM7G3�BAy�� ����,� ��=���Gr�}��l���Λ\|���x�ʝ�;z#Kj� �&g2B/z��ē���5\�Ť���<W籹�2O��L�:mw���"1|�y{ S)�,B����\�@Axr]8 �����o�s����J�$7
�)*�,+@;�D6�3�%��y� \���M���*�j�����xDwYW��k���q ��b0��1kL!$�EC� @!"���L�h�RV��&�Jh�L���`Ѯؖ��ԸWh6�uܾg�B�~rUa3V��~��*Vo~ߞ�?n�&��ޜp9�6�n��}�!*P`E�x7��/X
�9���,E@�x���cj{�3�{��-EH"�=h�s�y茜��pR�"�u;���"�*�o��9�s�}���"����7��1�����\�0� �>�A��A��/�����LJ�KT�~(~HS� A�u�n?��#8�[Q�<
��Y�ӶZ��qq���r%9�Lش�������}�[=���p���\�Ae�z5�k�����]���# ��VwYk�ͳ��
�o��̦��◐5K�uL���	�U@�V��xɅ�Dր����2��~�9����ۺ��ױ�A��k���>Ͽ�b�5�;91*]�l��dRՐ[j)	Z�jI��=���B�pv��^B:�f�~����K��x��U����դS}�J��DI�DIM98D���h��\/��a�� �#-0$K_r���jy�ތ����� �42�>��a�@ek��j�&T�A�J���j�#� "Ԕ1��yR�cQWX�̗���[�o��9�y�̓NH_��$�:z�X��z��h>�R�;�/�� � 	 pc�t�?L�p����m���'"�7�V��2^���A�e� �y;t� J����I������R����w-J�k�����&<Y�u ��a�i�ȑ�0;Vڸ��j{�ތ���p��6��,�W�wgk�bB!A�G�����m=��m�\M*�cF�%����0�
�a�G��{�kSE�yx̯7��a�Uv����~ � �'�V9�;|�H#��R�@a�4|��w�.��^�pq��ݭҟj'��ge.�����,!B�0��p�S�C��Roxg#��'��F�l��,�����c�ヵ������h��g��	U��?hu`?�/�G6��xw|�M �pp&��]��bf#�<?�A�闇��ƢaE��K)e��;��EK�d�c2�2�1���W���?U��v�.�7*c �� >*���e���n?�!�ֲ7�1��p�5 EhW9�4N��%�7���[3�//�W A�|@qpfSL�[x�� �> �S6ּ噁.Q�É�䮙(��lc�1�9���l���mM�w��}��z��B��&X0����3���\'��<f�뛔��z�P ����X{�5.	A84�U'��]�og��>���x�&���N�D�G�pV�^)��7&pz3 p�a���Dk�L�)qr���27���7޵ܝ�fxz�O_W>�LΉ���\%�1�`dJSL�lb%��p�.��l��c������"e�GGa��zk�ތ�
"�)R��բ�zo7�8B��	���^��!2��ja�
���M"(��:�0�;���@6Spȣ�U!ׇ^�94��a�a]��܎��γ������6s�����]q��p�}��w�m�<18=�F���Ð2��4�_V�G��/��<!x���Di���M*�5&��ԪJoő�[n����$	OQ����^�q�.��gb�+ؖ�[C�csnek�銘M�Hv#�ItɊ]ɬekn[4���8,o#��%�"�ctJ�f1d	�i0�X�(�l޻�2�����qmF҂魌�TcEٖZJ�p�R沰�q�\:Y��ʹ+�Bf�ɵ��i��]���k&k���l6�ZK�]��p������=	骡���3�|�>���ٕ�Ʀ�&F�%���T��̓��⮰|w��ϯ�}H0�>WLT�;�P"M�[�r3-g�1������qf�N�|�� >�|���j���y� ��`GgD�hi����@�A�_����=[։�����(f�8�<��tJ�6H������u=���M��>�9{�]�~�w�\NeM2����=�>�R�G��j"�/<�e���j���Gt̑�� Fc�H@WlU��ؙn�]Z�k\��s����	�k�ܭyx�ؕ6j���=<���� �i�Z�w���4"�^�^���拸�=�aDx�0o2��H���|�9���K�0A$ŸжA���;�3�m ����kr�5�ͭ���c��3����{��	��2��@(�M�j�Wh�in��� ۞�ez5��:�8���&X	�oI���xY�`����T�N[�>�{c
�I�ouث2+uv�Ѷ�qa�(�wm�}����Sr&�#`=��4R�tJ�?��иT��Xk͙�������Y�M�*>�]���
�0#�W��M�\[�fF�yb�GA� ��p^B$.���'��ة1���������1N���`�2��T� ����F\V�D�bTG����A�L2I��W�!K��x�(� �MU0�����T<ߨ� ����-�|XU/Q��j�T�A�}�UBoؗ�m�v�3���Y��K�%�{�5y fS,T�
j�QDĤw�u��|�`�I�'o�?�(�jm\X0ɚ]TBlKQ��[��]J��Km�������%�<}g�q��� l���`�O�_���E�	�5�;W�Wzßf�@Z���l�⪔MRb,d�I}�|D�Ҙ�<�.��E�	S�K|��@���{ N�B�b(k8�}b) ��	P ���f�2D��{��g�{آbb�*�.��zI1��]b�h�W	����!)����_��j���֤�����έ5:=�������EY��^�	�A�Y�MSM��9��Δ�,g�6�瘼���Y�{`���w_�7�6���殮�w_-w|���3G��p��*u�)>���˝���ݡ���n��j�����8Y�{_��V/o��A��ݬ���p���h�dk�<��+[3+ᳳ�{�g����Κ��JY�uyOk�$�Y�d�/7ӫ=��}�t9W�%^1"FM�v�/}�^�hӃ���h�*�H���o���Q���k��Y�w$�����3���ӯ��"��؇�a����^���3QQ8E�����e��=�|�v��H����}�j�u�S;Xu��H�2n�^�;���c>G���o=�az7�Ӯs��^�W,�|b��yCӞ�W�Iu�(������Cd����'g�ϫ��WM��}��r\��ض�=�l��Œ�����wݑw-�]�f'�gbY5/M}��0ܸ���s
V>����S7�Ò�����4�/�e��v����ni�=B\���'�4t�T5F�緼�.;�fu�N�2��ķg旽��ܯL����}�ܟ��Hyf[�P�jR\W��Z|��|F��8JI�!�|ҁc D������|���C�xoX|��f{�O�]�'"2|�҅��)�g�_�)P�	���8' wO� x�pN�^�!g�gO�OM�JO.���-�ѱ��f�l�4�[&�Ѕ�6t��Ӝ����)$�=Y�N�B���������t�I�K�х�6t�ç9*]�UD{:D�q�q � 8:@�zj�O�mB%I��ǅ�a�����ʒRF��H\.*��VH�B9��{�:V�HJK!f��:t��R)"DI�0�Wع	+�\�NK*����$�����a�G��ǧ+� IFMr�"�$�$�DV��U{.Uʫ��e�h�����|��쫒H��Y$I�sWt�K��C� @�@8;�;��h��:n��%$��ԅ�گ����a�f��k|x�f�<�I�9;���������B��H��R�%t����jk�q��?
̾�_/�@ O�����"���w��Pϴ����#�L�a����ݽi�Wy���BKm4�Z�M =��o7��� �P2���Q�:�nMP�M�nzW-�9Ɣt��爐�A�j�.Q��<���u�A �����'w�UF�&��-H�1#���[h����a�j��y�<~��$z�7��`ޓ�έ���}�/n������Yu+��^� Φ P3)�|A,(���@��[���"��A�sю��f�Wy����>�a�U�#{)gQ�/1{� �K���^r��$�,�&exvŃ�c2 5�a��-L>�.x`%��� ��&X�^a����!ڻh�Py��ɏ2 �+ݙ��:�zf^�. ����˽~v�j�b��>;Q�����Q56��,�Y��L-�V~���+�5�5��,�l7;+�o_��\�{���uy�����$=������M�^DM��7���2n&d�[�]{�w�"X7��5>GӼ-��w�x7��c,�p�"W��3���m�Ax@�`��I�:{���-ΦYf�KqMjmI�\�Q�c���t�x���V��R~���z�1�e0<F�3uB���W0���A�w=��胐��ޢB�!T�`M@"�6��S�#�L0o^Y�ۑ��Dt̾�\|�����*�|:��O:m�	u) �0}��@�L!&P��#t�i��sjb.j�=�՟~�NE�y�doy���l���o._q��W�Ѐ�̀P*X6 �*U4��\��R��<A ����������Oo�U7��Ŗ��ک��16K������Q��C�^���8�W9��ڥ�/��҆��5I�G�5J���m�`��?��+1Bz�S��=�õ���G3&f��b�CHrp��)�C�Ox�����8hq�}a��=�"X�*B��1�x����6��1x1�@�G��e���b�B؋b�/32�.����W����U��c~ns<M(f�;Kh��q^����ڪ�,�m(�̤�ݮCX����kk-�j�da��i�r�\���룋a���-�n���L�]�K6��QABX����e�f��a�V�%K�¦�����0LK�W:��i�1��-��5Ix;d�bKs��hEn�%�����7*٥�}}���R�����	�T3G$Ѧ�˥ku����mA3��H
�=��!`B����K����=��o�>��qYЃ�bE0b7��>���Wh�d5r7P�Y�L��ֹ���m�����7���T�a�A�C�|��d `4���(y�E�=�#�Fr��R:�)h��Uy�H ����J`A3+���!%���j尹��! ��`ǈ@�����Z�;��s��6� �4@Mfֽ��ϫ]����a��7���{��7*�{Z�Ӫ�-�����vk�V���Q���A��Z�RCfX�W������4��6��3�����2�5�t[��k2�Y[+1���E��NY���P'�E% �_0oT�oJ�̺�۵+�^uR�g||T]�[-֦�K�K�����"O��|fPb9��m�}1��0M~f��UA�}��<T�����}�où,wބ����ݜk^Ȝ�q[Zj���N d�Ej��uV2ê�1�� �@@�HF>��~�M��_����3_�]n�1w�;�	W�=-��T�%�n�Er���5���u�oH��p�7i�.@�.g���j�j�f�ٷ�̥ޞ��jFZb$�e"e�s�]@�t��b�x����Ed�����gwjtU�
�إ�q|^�����3�`�&�����6��2)��eXG���$��
�:*�ÿmu2���k�����t�o2��+݌_gv�;�$�D�Y����~>�O�e�RhܖQ��K`F7�����k5�3��`~����o-�#�<�Ro �T������K]Ge.�2����@W�� .E�Tp� Ԁ$�u�6k󌖕�<Gs7���
�h�uN�{���k�>�L ��S�kj۔4H��nS /k Nj"%��� ������*�m��0�`a�)��
ڣC�Fվ��e~�a ��*�{$ѫ9�=~ݱd�d?>�L���s����HNU���[�o�~y���]8��0�"O�V `���� �|8�^n�Rnڪ��( �;)���fl���uM�vR�z� A�A�+�����:)`�D@ �S�4���N!@�|SyST���k^R{Y����m�O_T�k��y�H=� �^ %T��S;&�� �ՠ��vbɖ�i���K�i��GY�:���MW�����Ye����>G�L� \v]-]ѕ�˦�y��k�yi��xE���V/@��x�Z�@,F�@,��;1*�d�a��L��3m�#��n���>�Z�,-�|"`kw�_�;�=��z ��DD�P#D>K�yɜ��˓�=Z���ǀ+�e�9�^l�Rkz�	S���Uo!�O0}2���ܶ'�R�7޷@A��D�}�O7T>�vL�p����4)�M���;�Pޞ\޸n���RᙷK��u�s�G���>����		�YD/�����YQ>�mL�jg�B����y�ދ����4�����޾@��Z��0\��(݁¦�T�csXr��;8Lњ�GK�j�͜K,թ���<��J�r��{������	�A�m U3{Ĺg�W8�������@�q��w��ȵ Z��bMR�� � )��f�hr �:p@�A�.�ٞ�\ҫ�O�0Xy�ޏ���������2$���Vh��B�y��`f��\np�|WU;��Y�փ+U�\�
��=T����>����֣��DQ�
V��E�������Ѹ)Eo�y\ Q�LG��0�����@hN}�x��F�R<PU7��R�j1C���a�Ա�&w�k��7�
4@U���o+���%�N�}3,���ʰ���TO�1ɇ+v������naCvƋ��v��(��>X<���}��Y[jy㙺��0-���X�c1���O��j"Q#����6��DBֶ-yk/3dK�� H@�$�VB�x���H�m����:-[U� ���;1��geh�a�6��Ibۉ�Ҏ���L�]j��Y�Ҽ��X�^b��B
6`�l����!	�M2������!6�[��:Q՚9rm̈6:���I\Kn[5
]��հ%o	&k�KaKbmcl5�0U�M�Y��5�3a�����\X�3[O���S�鉶(Ķa�:����,.!u
m����:M��~NZ� p��P>�Ro&���E�ꫲW{-B:��� }:�Yr&Pb&P\�4r9�)��ox��՛���W����	�'HFeCfv���a:0	S�� ��>�BU0b$��X�e[�����*�f�����j����'蕿���2���5؉/\���>�:b�]1��@"�x�k���\�$�z�Q纪�þ�@�փ+2��tu�<�Ү���|K䤨���"9<)YV32/���Ήh� ��rƊ�מ�j:�e�J�|�oN���L�Q��~x5�� �(����C&.Y��Hcm�sV=���FC�e��b]k��o��|�OߘP ��@Q@�]�g��mx����{ʻ͠��֨��!�'�� ��a ��x�!]� ����Eki�ѳ��-hv����&iq-u1���|��~�����eR�p��p���S��"�dcS��JK[�A����Mh��a���O�xD&�������z��uO_a�i���bA;L��e��3�.���|��1�TI�y��h��c*&Y�A�)�y��5����[X-�E�_4��%�y��j8Nr��d��^;�D-�t*w����z��t/�<��"e��y��zŮwʐx��nMI����=[ q��>?Z�B9W�1��s���L�r�A׺������� ���F���`�����Z������ԍ�4e�1 ������e���[.4]��h-��i2��\>n���+�3���'<�&�ugs'Q��q���/jSV^:�'�U�n�I��V�Q'��4�'<�4�Ӱ����''j���FCjoɳ#�u���yW �� �AL����5Y<���ߑV]_{x�oL�ȹ�^J�U�6[ruNq�̳��)��FX;�J؇��OfV;����V�.s���ǌ����ʇ�7�!�&��M��(њ�iju�1������.��Y!?k���;qt�^-`>�#�>B �-`[�e����MD0E����+�f�8n�]$��.ߦ����܉���l�^�)����3(,���j��h�gJk����T��pd
0@C-�+�(H.ٕŌ[>��%�i	e�Y �ǣ��j)��U��B�\�mF�GJ,er��F�#�V�~>������#���^�T��o�ڋ��ţO�:lD�!@�u0��T��D�� *��{�fg�DR��8x~��e��˷���i�:�)ᓡx�7����J�\�"w�Ŗ�9��^��m�m,nxErSGG]f�U�]��@�B�^i^@̯>�q�"q� B��㘀�V�����E��bᇁ�r�6�$��c�+�--�W��)̢��ֆ��g)ǽ:�1	Ѹ��2d��|L� �H��G�F��H?��H3^����/+��w��]�.߲A�LA���P �)
޴*�� �@����(&����L�c���.��`g=���)vSk{/ği�'a �"�1�e�q�poNqeQ��70�ݖ3�E��9�b���o��$L���0@ �=�Qa��y��L,@Rau��N�[_f.x�*��.7��k0C�zv���pu���B ����UPoPK��纀g�=c��f+��:����2��eN��P&j[;C+�������z<Am��AU0a�]ѼYTw���0B ���'-�,YK��^�A�f�A7i���#2�;n�`���4�T��<�m}��a�4Z�x0���
�=�%T��5�3z*T7?X2��5j�܁�����<h��U�nq���;g��K!]�֌��z^6wuvn�^?b87Ϥ����C~�c�g�����6i_���0=��7߆��w^αh�:�'ý�^T��3��ei��~[��2�R��=u9���u���a���v�n��eCF �Y�v�sG`Y2���mk�.�gqjVJ�I5�;�]�.9��P���B�Ӹ�=�8V�fbqn�����5�Q۞�c䇠��Ԝ��rp�5�7�H���vA�z!r�ݞ�ѹ�|a{��;ٕn��i%���+2(�M�����%�Yyu���{~�TY#��������%{�샙�X�����%'C��X3Ӑ��{=���dG^�)�R�ek�+|�F�t����c�x�i7�F�ۉ�|����w}}}��Ǎ`��$�ǽ�������L�C=�0ͽ�׬����[�bdϻ��<ÄH����s���R���;�?p��I�CfIS'ŋ[�cUNi�"��\q]òO�eٳ�������&Uf��toI���^��NR�a���t�Wb��^f���&kc�����a���A��w�aiڇ�����hs\������?{Ï5;P��<�=S|}ӽ"�?,��;ǄQ鼼�BТ�~�C��f$OX��#��0,�#�}���`2�#��.H�B�A	)�"H-�Ź$Ea��m7 �/� x��R?c�?�Fm`8,�!F ßG���
�<�j���h�C1� Ј�=�� #lj�!@�_P�L]A֨����-o�iY�H�+H�DiZ�kim1�-�4�!�l"�i�[M"�Ѧ�ьb��h�Z�kihF-�Z�E�lF4���j�ѕz�!������, Ѓ
�q6&�j��\�ٕ�&X� ̌"�LF��v||?�$HnQأ�.�E�.�L�(�D����s"�BF�,ÆϏ�������U����L�$�$��rJd�Q�j7)]6Y��Ν:m[���Mʪ��H�R'��D�T��Rr\���K,��g�M�rJDIU*TA˺�/ڵ�%W`�YK�)"�Y*��"%߅�a�����m�{v�r�U$W��HI!�.���%$$�4a������ꛕȯ#!�jVJ$�EH�"JHI"�$���*��fapt�f<8t麦�+��q&J���\�n*B�2'�Y'ƌ0������)%D�m[Sc4m�֞�1��eǱf�������$$*��6V�����b��m����몝H��$dI'é&8�a�%�BIIܜJt�ϛĭ	�cl(S�X��CM
b��J�E�֭�����vqIc%1��S@-ڠŊ��mz�r�2�nu�0j�ـV��ML�˒��ո"]`�G��
��+�XL��WHS)�sf��"��U�G<]6&�B�<=�q���]�$ۅ��PJ+����G5��+,�kIf6��ckn-�s�������N�)�饔j6Wi�L� ��-��n�e�5Xr�����\�Ķ�J�Q��2�U�k5���+l,`��-�m�Lj��h�"j��-!X�l2� �2�;2���u1p;��%�f�R�c�0ɦ-��&�1��͖��I����&�	-,Tm����.h��=�ft)d�f'W�m1�dHu����.�a�3u�\a�h��[�͕��8JiIX�o6����]�h�.eГ\�����В�GX岴t�JY�L5ٝ�q�j�F]"[,�VS��IZZa)�B�R�g)�C`fm�ZT��k��l���G[J,&!��2�å�B:�A�î냊�:$��9���i�d�S�H;3B��cm��#��VPl�ʄC:���Eʵv�z�nM2�#�qn���6u��ClX`��W.�������M�|�3|D"�kv�f
5a-knl����q���Ɣ,s�!�]�!�B.˔u��M��$\���1�14i5���0l��.�������k2���`��iԆ���Tv5�%���5�6ԣ#-���M�$���mn�!�ҍ�mu�ë�D�v�#2!5�բ9�&׬�᫴q���r�\���a�3Gu��TCe���e�GY��T���A�V*�j9EUEUUU[4f�њY��Bi�#e�"[sL�������I�'�>>5�S2�[i���.��s��^�(�˖��r��f%2Xқ�7(\a4CB�6�.͜�Ys5)�F�z��1X��Dή�Ic�t6!��K�R�ؘse��T6q���+-��²�4� ����˸���W����V��% �H��t�ˣk]Q�����mMl��W�����F>�ϟ��/�	�c����X���]1TX
Ǩs˴uv�+|�������"�!΃&X�^��9����v���Ɣ�K�c���%y:��Ħ� �7�Rbu�7,�-�#$<i ��D{q��`���F����CX�TuCt��3q��+���8^�T�� ��� ��կ�9�k���{dة���ч�`]H7��^�fXp ��a�}���|�"Aw0`�^i^M�cw��W�vݒ��n�5ۥ��K���o��(�T��+�L!WM�b�����,>��J߅ K!������D��>���x��(u�;Px��l�TYs{-�б�2�th
�h����^]V�X�'i����$����T��O�5��뼬�ч���)r=�_��@wW��+-�\�t_Tn�!� .�.���͘�Y����8Y�8��f�:�Hh��͐�,H�]"0�T�"e�'���|@��������Tc�����qq��^^egf�B�c'�U��0���{���s�VT�.9�~�@�I�by�-���n�V��d8���2��%x�fS��^��Cg�)HPcyx��
`A ̦��w�����ᇁ�!`�j ˿1�B؂	C�K�E ���&#[D���M�3�:��շ]��x�v��� �Jb�&W����i�H�Ax����}��[����99����䛘] 幙���Ćvα����}�5�1V7���L�k���1��coޖ���Xwg�&�<��e/D�/���ʀ K�̣� �W�	�Qٓu�����ч�A�V���KDG}כq�-��|b}�$ԭ��sC�7��7Gu����4��8��
Ƴ�v��͈5rifT�M�U/Qk�1{s�TἻf>�y��e�ut��o.�x���J"�8�/�翾Վ�o�h\x������Rc��@GΟ'����z�>��ݍ�!�5L݃������߼��"=ە�kg*��A�͋�^|Z�G�/]�!�(�!�\D�� �=���Ǹ��^W?����g�ޫ{�^��5�w������,��m>��]�3]5��٭e�W�W��Sa)4jR��,����y����{�}g�����y^�˕�]��}��w[ NE�v���h�rkBe`L@5K�!�f;Zu���η���xz��2�uĽ� @���$ʙ@L��]3O
O�X�x��^U�z�z�L�L�� *�}ml�Yz�ZhL��U՚�s�p�p�MmG �}�;[-�AN���f�_z��-S+��q�՟x�U�㘼��L�&��d����۝��xȜ�mr��b�p�@��<g�P	����L|n��U0=�rؗ����'j��!��u۠�t�u�@S(L�ێW�bl�o�� ������|_��[~�a���X�3�
B�-e!Le�P ��ut%�H&k|@�n ʐ��3�s4Ǹ]�^U�6�k.�����o<��b�ʰ&��H1��'i���#�eU��V�c5���M�x<˜�z�D�a�R��S6T��Jr�T:���6NN��̀ m�>�Du`=��Wk��KT�+H��i	��ʉ����*�X۽�oz���� ����ި^�S:ϭ���j��3n����MwQ5�HWHezg_e۠>�)i�jn���U$�0yۺ[�H}K>b���:$e�6��H������X%ծx���:����B	�FDa���,�c�#`�\f[r�r�Ryu4��6�1���&��2�$c	���Es�qi��Z�������H�D�OG��f��l(�� �[�۱�Қ �F⃲j�maV�hk�e��"��1�t���eP5X�]���.���A��lt`I�I��ڻ�z�ʕ.#��M�0tĚ���(dZ0��.�ʶnrиqr�L$r���];k&֜�+iK�,	�%m	ph����:c;�hJ���	��_eV�K,�-��G��]HL�V�e%ֈ�%������x�g�w�:�e�V��O޺i�]a��ᎽN��^*��aT�A��&`�GC�U=m�T�=�T�~yW��ޮ^���B�����ȇts�f��Uf�;��[�X��o��Z�E���E� K��HL�	�T��c;�X��S�{�Bs�2�o[�V�5tR��n�A�3x���"�}�:��)�p 	$?�π5T����9�N�fv��G�����7�����j�w��2��#� �!@�W������m������˵���Q�;�E�J�E3�9t�O��pZ�B�z "R�1]P�xu�E�E�I��5���,��� �H8f�����2�(¦e;�8���f𾁍�!0����=�]wF����\�"���aѺ��\=��;A�y�8  " c[}�����?w]ӾO;w�׆� �7owʺ� �����Z�mU��2��B&�A���7K��U��u��S+�+ �*�l����s��>..[j�d����O�Qoq�:�Z�����`�Q��M>�^�S;�^/�ݼ�V���#����^�e՛)� ��j'�;�ħgw,�ԦS&R7B�����4�Y��mSD���_���%��W��F�w
���U� gp�b':�'r���k�q2�O�Ĺ���,��cv2���fɩΩ�~i�{N���B�g�z�p���3���]A�v�o�����߳4=<7}t�Mo'&7C���5�T9���]a�,��?xL�<����L�����o���7���U	*$$D>��[��O���	v$��{���޺�z����򽯠0�^�� U8XzFg��ne�S�nX���1yY}���:��}��DD�/f��)+�V���ο�g�$�r�9�݊�~j�zL���O�@�*hUn;m�v�|c{�0Єь ���c��h��w\kUK6��M�Jݩ�5���U��f	��_X�Z�2�@�2z7jr:���]t�,����3.+y�c��A2�f���Κ烙w0��C-=��{������ߩ��8ƚqXB���!A	y��T�ņ��j "�d6ZѦ��0�4�b��ыZ�[M�F��Z�ҭ���c�F�cH�,��kcM4�����!�h��i��vz��i�=T�2�2@ڻ�n��z�^�ߪ��3ފu�&P��o �UT��ke�W���Ȉ��w��W�/���VG��N�d[�xLb��������mb���1SwG,(��e8�]�Q�ҭ��~Ȥofk��}7z��f{�s�J��"%S�UW#����U��
�g���~�g%���3?j���l�Խ���Ǽ����A�zeL��ឬ�m�Q>^#�����M���l�����׮Y�WF!�9ҁV�e�3&�d��	�ǉHe��un=�=u�ӼW4�����-��P��<G��nj^�8�^*�?v�;�p�̎�i�4Xk aTr+����ǀ�C���32�2��Aw֬�t�r�"�^��5c����C�L��&P���v�˰��} S7R��F���6��h�k�ͬ�:����,�X�� 7#���I`ͷ���ۻ�-��s2y�@�0�v�R7��tgKS�"��-.��6���Φ"*��������.�4a��!ި+�*��{{�n�1����e�-���7""$�7m�kp�-14�ib"֋Ab4��:��Gk1��ߺHXȒO>M�)�wf+a�,v)a�e���M�ʄ�l6��5�沄�k���cV.��!��1��	aV�ڶݓ��(�VRbRrB����R��	.�����y��4Ң�bU���e����%-�ln�[BlCD�F� є�J�l���uMJ�6���7L�Q͸�a­��>?4��dh�5pA�\I�L�ؖj�
[H7��%�H Z�)��@���#�*�>\��|����w��fV+������	���*�E+�;+�����֫��1u=E�<^��>�O�0�������)�٪uTʉ )���6�M�їO
��d���Ε�ˉ��A��e�����t�@C٨]��Bs5�g�˾������&.Mr�Cix�2ޙ��ʙ��緛�D;��mg1���e���u��@S+�P�*/p�c���H:�ÇA�QƗ���Y��ŭ"�5f(o���V�mY�3g�>���HB��������~���O]����Gz��<l	����⭜��@V���I\�1T����8���?f����y�}�T���>�9�^�S-�N6��,�x7��p�횠j�sl/+KI��X| $ $�cLj+��	���g�e�w_-���fwux���Jfe�o�(_c�Αׂ��K�F�Z'p(^Ϊq2�*��U:4lC�齴+7�@�b�*��Ǝ����~ꢤ�l`��b�	վ�L�J���8�U�U\ >�W�n�ƍ�w��y�l��B�VS��O�Q�!S�8�'�;3��-�K�+�f�ju2C��,��e�ɣv�����}'��}g�,(ep��31�����t&Z2)��k���e�2� ca֊x�����h�]O�tWUf?T��< �]*�������r��/@���2�2��0���\���D�_�۷�/���k��G�?c^�����uc	��sFN��秽����)
�bm�{��-����H0��pl���-ߴk����g�=V�k�����a��}�ؖ���A1����a=�zל��e�Կ.�ޣ=��{�R�����a�Bfdd���r��.�<�0f�]��"��n��K<�iJ�/s���ý�3��ᏦK��9�綔)'��	�)繘��{F��QG[i��y�fNJh[͏{l\�^���]M�
s��wĎ�����,�P�7l��KzAo�n���S=���z,�2k�:x���uB{�sU���)��!;�5�`��tG*�=���ޭ�1}�4{��LQ�0�s�n�a����09�����+āR7���6����Vo�w�o�>��]�MCt���$��z��ެ;�w����<:�������Q�zG�2�x"uo���/)��nio�sS�^�l�}�oZB�wo�oG�����"���y>G2A���d�]���󹧫�/{��ub❋�Z��	��v33�H�|fg����'�1��#��N}�-�9�'���8�����ocO�b&{	}��\7�󢑝љ��-���W`�d�{�|�]����H����z�5N29��=��wK_�b��U�����e $ (�y6&�0�e}�{b{c�V���a��[g��!쪞��������.��Z��M1^F��Z����Ϛm�Vfg�亥{$.�q%z�.S!R$Se�a��OOO7U�UR*���*K��I2*�+�4zxzzzo�|˫�t��UY�+�eg�[=e6��<ݗ�}Os��>>7[�*�(IT���*��V�U+Ϫ���L�V%�,���O��ʪ��A%T�R�Jv\We)r���0�ӧN�������*�=�\�#��Q&�j�j\��ʫ�م�l��Ӧ�:�>t�d�y���6�ͦAp���* �*�-],�çM�:m\�q*�Q%U�E2�_G�F�	�FC"�ʻ�;�t�U��Z����<>>8|n���:���@���S�:ȩ%�%.+�!KU.�5p���W$x�ĕ%J�E�<�Վ��u#cӂw��JD�, ��  �0�f��_�e�w�������	ti�����H� 6jHEh��10�����6 S��y�9wF7�axw8'�W�W�� Ң�{&E�z �b��y��ڬ��z�	�2�NS3�d5��<�\�0A����|�3�_��Imv��/�vn�4�M����1)��ђ��������^�Be<ٺ�]�������p.�g!�e����5c�&h�^J g��P�lws��r�6�Xȗl�o�����q� 7�E�]�cL-�m�|�S�9S�����O��AD��gtZ���~�@s�a��B�{@�a`]��3������m��V��A̭=����;�q�9X�<��+��0��1�s���^��Ӆ�y5^�L�F�ݜ��$bʉ޾Z�2y�F�5fu���{�G�~��|]��SOں�ߏ�}����3�?͕��^�����Lf�|"�D��}��zg�r���Zpqs��������o��U-��Y����Zmf�L�*��RͬqH2�ðL�=�]�^�=
����W������1�gq���]���S�^�X�v��A����kP��n!�շ4��_4�ˤw �w�UV⼡�\�H��B�L�3��8-�������"+I�S��^��z����p"3�FR�q�&�=c���+b{u�4�f7L���f͞��@n!�>�&P�S<�覱�+�=��Z�����3�9���.�_�gL�w䵈�X�Cr�%�j���F���"�C�V�}3�������ͯ7����X������9#y�d��P!���McYm��X�3BX�Y,aɥ��B�*mWO��N�Od���O�yu���W��AXlD�M�ą�-�Yf)aQ�R[���G	���a�Mt^5uJ��F-J���phuS@k1s:�Zॵ����<%̳VQ��[��Ib��K5��@8!X�qJ[sl�W����z��,�&kp�J!30J�Qu6��MnWs ��&�XX-	{K��ơf�.��m4f��i�����fM�N&���WHҸ�6nb!4�Ƥm6IE8�p�[��/�r�e��0E�7�*f!�a�p۸�)�@��na�"1��-��D���%Q=����B�ҙN����雺�P/7*�ezo���b�-`%�]
�7|�-�{@�ofU8�T@��=�۴b�L�u���:ɾ�S�"!"��|�A:��'%����O����N�!,�����a�:�u����] T�W�j����7�W����?�^	Ynuc�iA�fa���H�]�0��f��P�_>u��F� !T�R�ܹ�+0�3�?k���l���n�$�xX��u�"㓄�!�b�ζ{�C˄�wm׺�z�&����|�u���n������G3��K���۝���%�y2G�Y2^E�r52V~�o��:B�B!8���B���&���юc8�1��E�P���3���4������fh��x�y�vU�����VcuGt@�a2�UT���������kͳ�2�Z��""#�b,�8L޼�y�~�ɮ{�<Ϙ��z-��gt��T�� �i0UN&n��x;�v�ΗQ�'��B����q3��vfόRr�O�0%1���BR_��@%^(�A2:𹃌���&��մ�bjxS�-��R'z;Y�=�duC �5�k.ŕ/�����K||X
�K�eA�bɜ`e�yv����GC弁]�q{���X����B[��Ҿ�>��Nh�?g���s��.��ތg����R2��R+���m�ͰD&���ھ�_�.Y�-��E�ec-؂��T��61��va�| �� @ UF��h���������^`́Q ���;�<q�X�;���wc��s�fGTw�� F�%�]���y�$�U @��Wm����� C�L��U3Z6��
=��v��-ξV�����|?`Ӏ��(��˂���۶�f�#	H�&ܑSW��}�o廀?���[٩lJєWa��
�6jr��

����J���?� ��n���C]�\�t\�^�g:�������/�}��F�v�@_Z����A��u�r��/���t�����m�Q�r��@5�U!2�
��[�65=���E���Dʧ��'bV���f��F�
��(|G#٧��]�ۜ=���	��}�o�t�����C��q=�o�x�bzN�l�ݑ������ 	��<]5��� �]3���c��8����kh�����m�93_N�˻���?�W2�f�۰��$y�'�?3ҟ,tkEi�A\,a�F�K	Cf��C`�<YI�.pqH��HW����n��̵<�m�Q <����i��xAǇ���f���ʲf��߽�s�3�N�`�A�Sw�̭ev���s��nL�wN�����2���VM�����w�m}��Z�*���#���	H@P`'�Y��M���M*e5흭Q����-��� 0��qU.�S���������L���ڛg��d��6��� � ;0`.�#�NrW3MViQ|��w������W*8��y�7㘩h��.kK�$�l�CLf��e�Ʃ�q'-�����g{���yN� �lH",�3f��oXZ,����A0 ���i��!f��ڋI㿙8$��Ϙw�>f-1��[(e�Y�8��x�|x�C0ĥ�GF�,M0�d!\j�ոYu�h��M4�5�0EW5Ϊ+T�Ev����k,����uc�Ʋ҃{K�n��T�ʹ.�).Qr�;.!n�n�a���5`ӳB:YHa�/A�"�e��ىZ�
\���+U��-�^m��na#� &��}f�p�5�̺H
��qҒ��GV�h�ʡY�c�>%�k��t¹��(˜��u9���B�.�L>�"��T��G��{%�so����@c��������@�����y�gd�D��%��.	��awW�tw9ub���i���^�M�t!T����U���Z/l��5	�s��]�_#'3;]�0%�$�l���g�7��h���r��o}�Ü����h]L7���d���k����`8]�W��5nI݁=�6H%9g��VݻDȐG;]F�R��p�I���� 2����-�jQ�U���&�����JU��v6 ��%�2� I^�B�*�SYN��8�ϛn�0ۻ�4��}��k߇�? ��*�מ[^�+��?";1��G<Bv�]������������ �	 ^�#�=?uw���'3;_Ø `3P��&��v}�`��<����bk�+�0�;�Ss����k��-�y�"m.�	����S���6<���7��eXW��L�B8E�k�V�i�n�s�Ǘ�W��@L��TKp�4�bK���Ft�n�̺��\γ�d|#3@~�ȼcL	�'�S�G��SR]5��#��9���Z�	s��
��ʺ�䖏A����2���k�s<�s��-t�{ӓ�V�hF0 *o���e��J`��� �Y���2k43�ܲ�p�';)�3�K!I��.*�%Ǯ�BeL����`�-�&���pE���I���5��sR$ͽ��{r��+z�N{fƪU��F$�1�e��&�8mkZ��R�h�o� @� _}sן}�Cfe^v/�:��Beze@���5Ƣۤ���pʼ��'q����O	�/(�D䊍���`&e�fgm�:�����;��>�(��Lp��pS���&j�Cj`������l���L촳&��&�@i�[�^�6��ON�{��oo�" �>v�г6�x�7�y�� �v�<@��;��ʙ^*�����+-f�K��#m^���ܧ����o�]�&F��Լq
-�3z�	�=�4B�W�ӷ�R��%FV�cV�r�\ˉ���=���=l ���8�O�]��O��;N,������Aȝ9?�?̼Ʉ�񒞘��d��zf{$GU��2{ŷ���V.0P�9s�?�_&�	q`5�I�^��<% <W|*W��(0L�.�Ͱ�{�
�o<����afֵ�����W����i�������=�}"m�XV��˺aRֆ��""[r �Y��SP�K ���-	�����#�f7	�e�]�Nۯ
�&�2q��[=���>��/�ch�%k�rP�ݯ�".��i~ ���-6��E�~83���B���g�����SBclV�(���.��eO��h�}�o[SD���u!2�N_��[t��U;�P���I�=�p�xPƔͻ�-t������2�#���?9���+F���S
�R���v�n�#!rw��"���ă�_��'_v���Ɠ�i�g��}�x�i�{Y�q�'�#����7�x���=�U2/7R�c'r=�`wylfGsu�L�d���x�[�Fdݷ��{m����g$T�����{3�"���/P��1Q݉�]u"2����sW���q��`�,�=�k&�}���ɉ�
�Q�j3��[Ys7Ն��B�4{��֑��л�d������/�s߹�[�����0i��{�u�x�T��2��Ȍ��aw�X�bY��e���}�.A���>���˶	0m!��W��6��fp�Hw2���?`VC��Q�׌x�FW��}��j�&Z7j*��j���}sk;����؛�Wx����f�Z�}��3.w��7��i�uˇY��#w�x��
ӳ�+�i�[י�y-����o��`�<�^�s�_[��tn눛�g>��=�A�퐴3S��j�a�ݒy����N��ol�������Hw��29YG���E&��4�%�3��x�}�Wc�����j-�=�����{��Y�.��]��L�ݞ˅ʮ��r�����j_n���4vv,�4f���N�6�[�'T��k������s$�,wr��hq]0����h���!�n����wn�P��eX߈���\r1$aI�>�HxX����Θ�3)��tP܂b� j�J�
��xh� �7 `�8p109�<7|=zl�EuA��4�ZнCЁ�?�E��p�	���:$�"O��3�i�X�%��Ukd�/�w{�i��Wղ��<em~�@b�SN�hr�� ��D>���CO���?��@�F��=���:CM��#�F�m��4�a�1�1�j��x�x�#ƖYm1hD-m1���1�i����i�1���ciQ��i��m-��%���:�C��$͂�($��j�`��)��Y[��-A@+Mk&�|+�g�DKro�������I ��2SIRUW��55.U\̕Rd��H��0��>7T�T���D��℅�qqUpH����r3��t��6t�+���
�U-+%T�)̼�E�H�J2=,�G���|��Ϝ�j�Zo[o��ZS�<��O%U�.;)Y�U�h������rT���ʑWw%Q"��%:w��dH I�;�F�xxzzzx��>��y<�b��-#hf�.q%J��d�$\]�==<V�n)qI�d��(�K���Ur�5L0�����l��!M�l���RIp�D�J�W�K��I�IIv��0�G;ORS�I��)qqE�IE®V�ȦJ$)�(�ME5(���IY�qU@��s"JrD�����Ǽ�*�>���p��jͣ`KI���N�E�K����]��^��Ԗ�L��m�]7;�P��m���6k	nJ�.�Y�B�ҭa�Ff�;F��).�ή�Y�Yl�㙜j2�Lh�B��[j�Jքt�"ua5��&%n�U��,u��:้*	p7�\an�6�� �.���Q�Rm�i�1�d���Û����Iu�+���WB����e��PF'f�6jlb�� �)f�;1`ib=t%Ћ2J9)�ha`�Q����iiKz٘D�n%�u��2e]s�&�V�i�m�4��u��\�!��9eW[��if�l��#�!��0��چ���Wm�(ͦ�U�l��R+�-+a�JҶ�N�h7Y(�śqu��Y��V�#���t`T��` ȖZ�fR8�������l��+�n*�Gfn�Y8�Q�+U�L�]6���nZ�&L�\mun�Mj�	�4�m�$%4��ؑj�j�\�W WGJ0���lM	�tABՄS2����.�r\��mL�KZQ��e�e�j7keV#�\��[�(-;=0i�KjU[�3T�N%���	Z�&e%�f�\R��,�.4C��M�u]@�n�t��C-0�I��r;K�h`��9�\�l&窀Fi��&E�;K��kn�0�5m^\^R�n���v���p$���"LY�\��=��arqh��+e��s��NX ���X�]+jL�P!��8n�0),mv�,�^��Y��X0y��0��HJ�	rY���	U;�m�,۔)v�xՈl.FQ�c\����c*@�Y,SMvJ�&�g#����-��)p͆�����	�1U˔j�UUUUUUV0�"#Z""4�ZЇx)���CbA~��$���Y�	�ڹUn�`�[�ccFb$�Fd��B��^�S�u����KF2��5�ۥ.�9ׁ�U�jeҙ��XQ�\�L��퐚:7����1�(u�С��%�ѵG;4�f�r��.���Bk�m�[@)	n� �@KQ��F�c.2e.��p��=�dp���c8��!�~��?�~�@a
�.%j�:ʸc!�K���غIس'�A[�^��ʙ�����`�zS݀u�����ށ�e�-�	����]�]10 ��p=��� ���Ի�����}��-�XL��\jbD���@5�@ ^�^wC@5]p3:�06:��K<^q��B� ���^ ��dyګ�ͭJ0 6��tԄ�`�/�F2��Ҟ�8V.��i�S�xu0�`�p&K�a.�]��;ᓸ�Z��ʶ�k����s3�}�׊5����#�A'���H�1��m�JZ���@�l4җ�\�ɄԢ���	�3' v��4��%T�u�����Й�8�P��#kr��n ڪ��Sz�	�u��v{��#��h!=�wO��|�Y�|&8f/OPO�-��3�5s/�ٺ�戩ɜ��ճdy_�����v�ﻛ�eW�� �.�����x8dUs�Y���w ��_�
��D��C# ���� 	+�7���lt�'�;75+ћ���M7:� ֔��E�A3.ǁN4�F�=�L�U�n[{�h,���s�Obv:��m/U����R��Ux=DC�נ�`H���l�=T����j� ����Z�o9�o�����Z�-x��^i3/���|�65�h:�n��,�,u�e�dH��TRD��S[=��+�R�gWgbಲ��x[�B�gݧ�r�7XUH��T�ڈ\" A�͠R��׷e���{�7�S�r�D�^޿I�k-��:P��2�O��~����S�ԯ�2SH�V*�O��{�q&N���GOfgM�{�G��g'�),��,��~ >>  ߢQڍn~R�~�B�2�2FU N6c�ٝ�h�r ��.Й�����us��0�Yn�Wx6>d́2�虓%�`H�D;.��8+��]�u�t���͋%�o�_��A s>~��?V�j�k4u���u1`��̖K,�F].b�, ��f��D6:�^��±�Z���T��]7`f�禰ϻ BY�2����MM�B�z��n��ѫ{�pX�qL��+C �O��3�d�噬1�Ջ�eL��si�)��i�b�	gε�zB�U!2�����@s��8��M�v��6�J3
y�7ή:�u���7�񞵎t���C1��x�T��t�:�,n�pn�<�����qF�X��5dXz�5\^�}�Mɾ�kԐF*FG�� ���ڧ�4
�J�3£�.�s�K�*��8�X�qw;�p�reL�yh�2A��^>M;)�1e�)�	eRk���K0F�P\\ڭ6r۞.]Ms~��� �.]�T��+����	gε��D��fj��ۜ�Z�R�A�`&]�讶9"����9�Edb���Y���Vݘ�x�zF����kf��5RY�������QX��w:���2�2�
�e�V�{�u��Ck��G��C>u ��=7���`lH�n$	T�T��צ�r/i�@���[1��Q���v�_fp_��W�ɩ�P��cǧ$w�1��s�_��]��z:�%{��Y����CT�̎��w�I��!����yY`^E�!X�d�����^��b��y�ή�1����bb4��Yk�5s3Z����fj����B���m���J@�M]�vPf�57-�b�.�t���[."�SL�tEt�sݪPƪL1�WR$�� �;B4^X1�F�Mh\ت#4�[	5M	(�$qWk�\����l�jVhbܴ؀�-M	v(����cs�b˭z|�Wƾ�6�adؚ0���+4�j�l�.���V��7]�	����?�O���8�٪:�r��V���l��q �i�`ָ��[���3>�+/�[�yw����0��ʙ�1��ݼA�� ޻B�ze�`�|�rC�;֕��;��Y��,�al��U5o�d�=� ��M�U)��Td�e�L����#��f���j�p��\ �H
�$Ux�d�+��T����3*�T�{s�vo6;=�eֽ ^Y4��D>w�V 3� �	�5Q�T�(�ہ���J]'h4U�}��;@5��S垱Z�Ok ��	Z{���'�ݠ0�Mj�&�r隘���v�TeMWvob�'Ķ�1<���]� E@@��y�|f6�1ڻ�y��Yz�@on���L�^���~�2�k���݈�qGM���H3��K��� Ŕ�/p�DDw�\�1c��:LM�o'��T��O=����g�ApHT��~��T��g�����-x�Y�@"-J��v�6���l%b �+\�=T�P,�旃�Z*Ms�zӝ`��̀�b���e�f�ez㊗藞D�|��B�c�]���lj����T�G�z�_�� ~�� ��D �BX��`׹�����[4V�-�*�/�zW�*ߢ>������LP�#&58MQ��.�z����]k��(����&p�8x�}�p�`ؽ2��i��7�s�y�cзw�$w/ex.��2�ʪ���چ�O}����]�ϖo��1���hM��0 �.зV��	����-Jvfe��"���Vnv���]�����zAםf�rYo)����=�32�R�{�^ _���@ �nnaڥ�'1�+>�x@�E��A��B "��h��/!0��b�^�4�u��s<s� D�.�h��tS��B���@��6�� �uR��;��b��7�����Z��	�����e�[�� �#!:�+d�W��s߰M��;\l� j��JP�	���6$f"��7#�HAtPH��~ćz�o�W۶zk[������\]�o��ˉ���^�.io�r�bp�[f�ݴ��᧱p�C�4X@{ @� B�0�y�&�xO�O2�T«`I8]κ�jz�WY1��pxfx/e���B��*���-�V�ܓUx@ml�"nw�d���E[�����^{zx��
�j3Ɲ�f1jY�4�4_�b�2�2���+-�=E���3 i�����rqAD���u���p C))[�"T�h��V���ĩ�j����R4~N4��أ���8����ظ7��yZ��o;���T0�̷{�{i�؎�˙��X���f�cfQ[�c,51���2�J��2�4�b�Ǽ�����|+��d�j����e�-�����2ݰ�6@W��"W��9������e��g���G���]x�ʜG�$�x3���xR(L�"�Ĳ�V.8�>J5����.K�o�	��R@U0z��Z����r�^��Cc�nz�n��U��ib�����B�	�镀����9����\��s�e��y�@�p�
|��{�h2��"���L�)���-l,LV��&�L\l&�~��y�7O����=OZ�ϴ�}��G��~������;�"x�t� �r跚�^d�by^E�>j�C�g�-m1iF�dgi,$&�j:��t��qi�����^oě�˚�eIV�@"��0�l�b:�6���j���0:m,J�n�1LRh� vԬ�D8��sdj��T-l��ڙ�	�6\���mr)t�4v���aI#T��]��F��4m�\mL�2\Ga�1uh@�����hڈ`��*�-f%m��(:���`򰅛)�ӆn�3u�Bh����Z��
 �]*ݝ)^Ֆ:ۄ(7
	Ġ � NC�����@MC��mqanp�y��b���.XHA����H	��$��.��4��0!�P}C1���o*�n��p
������]��2���>�eL�L�A���:~�뚩���Y2���]�/�2� `W^��2���� �o��7��nظy�����i-�י����%R�lz��A�i;�g���g:���n��؜n��@U/L�3``��6K�*�M�o� +����$%�f$$�R�=�{�2��H<�5[Z�e�&U��M�Dl�ӛ��*�������:�=��L��J����N�r����U�ռ[`��Br�)�2��>~C�Ӑ}[��'����ؽ5���*sL�8��t���ɪ�%z� >  �`��d; 0��h�|+_��x���j���׏q��j~ �"'] �Q��jV�<��s�#�t�9l{N��_j"r:�M�zj@c+ޙJ�A:�	�H�ǀ�`�${��q ��휝������S����:�X��y8
��p�M-9��<���Gv
j�KD��ׇUW�k��ɦtێ����Z4�Ir�Z�����$�]Ԙ�h�䮋�^�q5jc`�F%$�K/��g���x
^e�L���[6��TNG_��h�����L̸�S��k�h~�oz�v�͜��z�z��]�3E�X�J;UkQL�A9��x��k�����
�e���݆�5`����b*䤲����l��	�0�;�Ma�fg�W���=�'{w�n�	'Nf}�3���ۚ��i��ӱ�!�:I�7�5�o$�������p����g���l�}K4���y%��hԕ׼���=Tؼ��r��s�n��m�8��!���~��y��f�{{��Ø)�ei��I����3�V1;�c4��J�P=��6sxūq{}�����w���}����.6Q�<Ҏ��b��v�'_j��c�dX&���O�j��ﰾS�x�o
@*�@�@�97I�Ѽ��E��j�b�'	��3�riޓu6m�����}d���FG���nw��w�j�'�_-�;}ݬ��31�N��C��&hy��i�F�]��F��54�q���)�ZS?��0��=l^���U��V���p���L�P�>,nb~ӺS�~W��>�j:���ϔ�]Ӹ:��|#�w�2V/�����"�HS+<oL�̀o%���(���2S��1~9�Lr��[
����������%w��q�c]�[8���T�s���ۋ�lw,^�ov{<w��;g�Jno����|����$��%�sLW��V~��y��+4?nw��M�h���att��4�.zMS=1�x�!���(@;G&�zE3yk;���`@e���]�� =��D�8���$V@��DIܝpN�7��i88Ϭ�<8a�Ϗ�OOCu)UpY9�w���`��D�)9'@�==0�G�����B�$��qRP��*�����v&]R�J$R!�UʯOL0������"�nT�"��*��k�
��Z�T���Qr�T��>>0�g����{��Rf��y���ѳ�E�\e�W%\�j�=0�G��OO7�Ud��UII�D��
n$���,�T��Ҕ�U�WN�0��ӧO�%T�I[+gǞ/7�[6�y��m[)��====7��UYĊd��Qr����	����$==0���gOEUn�M�O0�[]h�6_L�Fލj�ڛZ�ڳSJH*D�ԥ\���ZA"J$UH�^]Uʩ��;C!�
�?|�w�Y��W	�_�&��S3.-�b�@N$1��rK_kF7KD�u� M`�a#�R��{=�|1!܇r�	�
��R�[VZvE��VoO^v=S=W�{� ��@=�U0���Q4�(��B����~)X�-�-�Aj���Ʋ�FWR�B�$Ź]�. ���������&��쵈�	�]8���Qq�@^m�5M'�K��Po6SE�\' ���ښ6�o=�NO_Sz�D�M�o�v�e�A2S烡�3�F2u�E�ͣ�T�h�b{�@3K�e�ʙA ���S�;��e��ifȶ�_�q��/N�]��([�P�[P�8�8{o��߸`y?��b���xY2Cwd3w<�w���'��T���l����
�uW��6o�3��=�
���hU��f���ng��5�9�z� @�^Q.&q�v_oYIg��)y�	���G��i��Մ�[P%ڷ7����V��Ѳ�gw.S�%@�^t.��W��j�0�S���0/���b�1��j�}\���L�CxUNs�o憮���^Ѵsm��/º�W�W3w�unkv}X#�m��л^�H	��v%��x���o^MlJe,�|j
�֊--�g���P�^٪���S��\1�}tj��{;�k�����\7���A���u�.�j�8x5X��c�\k��5 I�#ޕ64�p�6�C4�8���R��b�"6)R�R��wAe��<V?l��}ű�ﴵ����=7*��K>�~@�i�� �R���E���Z�!�F؈bY��R,�P�Pg��z-���2�s��чX�h�.�u+�`��6�Y�E������6��HŦ�p[8Ò�n���V�bkɘ4����kR`X�3��ՃfF]+�V��Z�Ȗ��*�C���4Gm1tqm.#E"]k\$��
�j:�-�i�)076����7��݈�6�5�ƚ�P#�y��Ѕ�߽�~����;S.˪��Tz�j�*�A:^O�%9b��| ���ʙS=��Ϻ/��\d�pz���!+z�j��k�N� ӆ�s��͵-f�`�C&��)Q)�cV���x*��3.�l� n���@�@!T�kFÇn֡úT潩�Ѣ�� �UUL� j^�lJl�t7U���^3��q��X�]|*\l�B���N5h��
�0	��UJg_*"W��c���T�6�pǞ%ٗ�ȃ�nw�;��D[?� �ԿJ����]2hvmq��c2�)4j4̮]�;���<�t�J�`�2��o+��Qj�|@����p~�;{:"�*gl�	��v�`ej���7��U��nY��4ʳg��o[�o]���Z�^m[=	׌���,�S�qu�ݢ��S35jm�3*�S�kE����? ����{�{7���ћ�1�����U/	�9�Y��`��ꨗ �V#
��2��Ӫ��\-�q{�e�3 4��%� 5�ԉ���3M���F"�hZ+�??w���b���X���8�C�eN|��j���1��^�"�U�7�܇��j�x
5D�X��o2���FF=�Y�W�҉S2���LƸ1`�(�	�H7����ƶ�(�����R�"�8ѩ���}��ꪉO3w��Ryێc�Ŷ�+E͡�u��J�@L��f��`ez�`�ͅm����B�нT�KAgc��ӓ7�L&���T˸&;u<%�!0���˽%�(�o=r掫}ڝx7��>��[9l4զ�u:�0�׏Sw���-X�K�-L�G���� ʬ����1��;>+©ze	�&T[[0�N^wY��vu�e ӵ��b��9x�6�z�dG�m����K�k��^�xU/L�Q�����g����sY��Rֵw��3��P%Й����zl���
^�m��zH��x&��L�������������6�Fg`�I���Z�`v8�Wu��#�4c��v�;6�^ا�.�	�	�(��*�dٓ�;w�.*Z�c�ȍ���-1׋H1�@�`3p�
��|轨�fc2oo��;mmw��3���2�.�Wc;5��a�dbS/y�*:�Ce�e����Ь�x%i�ԓS�V�|��C���=��w�����D��r�?y�m};'N1��ݹsS��)ڷ"�
A E/P��I-���ؽ?��ER)L��g���o���s;ET�T�RY�kڪ���m*�+aQj�@`��,�ySbN$4u��dF[��K-.9u-]�=��j�w�ߤ���c����7��X訫�1u�`s
���x\�L��U0j��vS�M���"�s_UNh����� 䦪 �����"P� �N�;�2���L�(�!?`�v�YQT��IdƉ�؄�p�Uqƀ�*�t���4f�F6@�^�^<:�3x�Uw���^V!NϰgD��b�
�KQ�mꖱ� `��aU�X:r7�]�go�*��p2zD�s�����FE[<X�Ƈ��Uu��M,�w��H}:^�J���9�Ixc�w��=}���8m�˞�gW ̀0Cf&A���*>������c�Q�mb"�Ŭ�Lx��0|[�\B�س�O��=<ON�&SMԸ,�IF�"fطSce������h���UF*8���KJ��0��̼�%3(m��$m�r��Y,u�f�&��@��Y�X��(M�R�����K��G�Y�WR��0�Ś�񍱯U�d��rJ�U�u �&��1�����E�q,:�y�J��crf3�-�7]g3FDK>{��>��[6�
����Y�-V�)2aavjС6�1��z燾�����
����3T�g�ə����Fr�7;�c�eB��ޙ�8֓���A��x	q���
���:�`�]����z�L�.�됱xj]��}UJe��$�yK�����}bn25]��o\/
��R�PS���mP�3j�%	��K�E�ɉ��j��1��^9tΫ.��w�e�0K�U^�pyk}�eFs�x\e�i�9&��w��ҙ^/�b��sd$Y������ �q ��r��}~_��e6wS����@"59���QWg��+��0A��8�"�j�e��U���"�D�Ŷv�S�lNSըw^� 8��iB%8$���n4�E2�P���8��*��:���kmN8E�8{�-W-WF�]65��ilKk�����@����7�To�G�H���|���k�71��v@���S4D3�KX^/� ���������g(�f�7���q76ɪ���м.����U4������@L�gtp�}W���h����|-��И�:�/2�ʙ탐�fz���u���%>��i��j�d����!LV��*@�> ��0��P�m,�ge�d&�]5n2�d���5@2�k3;�ٰ@g`&���۝���pUE� �މ�]&j�_g�D���&W�n�ڎ2�d�otl�V����!
�霚ܹ��0U� n6�p*�4�L�`�aر�AvК:%�����N/�W��3S����$t�ޥkSv��?��=Z�n�X�j����5C�R[YX%�e��>��ohJ->�4��=��: �a��U/
�*��[ϣ5��	uᲀ��ݱ��Z��5�y���P���R�q�يe2��`"����s���5�jܾم�n��;9�UxL��I�7Yr�1�%dAI/E�$[�.��
�\RT�B,FY���0U!`P!��N\&��S<@��l5S�5���q<�Ǝ|M@ƺ��<�UfΗ��R� 	f�	t�,t.�m,ҙ>�gx޼�9�J���S_(��  ƨ� �����Fyz��rY�:� �R�@T��:&��e�Z�f��z|�� �<ԢW�W�
�k���9u:�t6��j�7L�|�_x�3>�5g���Un�§�w�P�3o�p�X�g�ĝJ�v���ݙv>��x�������qt-۹���!�i'�|ٗ��gwwB �j�-7L.>����}�J�ߩ���w�L	�����/뽻x�K, ڟ}���Q���sZ�KLV��f�Jj�9մ�M	R]�����}���?t��UHwov���V����|�2�эn�aW[�;j� �U;J�y7��Xi�NR���+x�3��wPԅ�	|��b��B����!��_}m��W���U�V�X�MM}���D�R�����i�9�ä^]���� ݻ��%f��zY�����Ori���l�h���Ez�g}}ƆQ^�4.��P�˖v�3lσ/j @J�3?����?�x��^(�"����*?�!����3�Օ%3����_�QxjT�i,�o@� ���`j!��CB$`jTz��=����U01J`j�`{x�(�(`h���T�@�02A�� ��P00��< `eT��P@J�  ���@`b`jA�� z��T@��UXJ�5P``����^�� ��[*�T����X���X���0^���SP��05KU0����X��R�±lL���KT�l���X�T�2V��°5+ג�baXج�������=�t��ߟ񈱠EmTL٧�t�����w���'ۿ�����_����_�?������?��n^o���>��?�w���_����)_����EVd���W��u�����_¯�_��>i�1AU�_������1���y����W�����_�/��y�}�ἶ��<IAZ�j��b�ZҌȳ���-�f���b�+YLԶ�����d�����cQfKXZԶ���ȵ�f�ڋb�S-KY�cR̖j��Y�֩�,��Rږj�Ա�l�օ�TjԶKZ��KX�5-�ɊږZ�Z��42��25-�j4�VE���R�-V������ZI��3T��Kj�Բj�Z���b���Զ���Y-KV���KR���Kb�MR�Rѩj�MdXԶ++d�����5,d�T��i��Q�KMKd�M(�V�ZԶ��KZ��mRڋj��KZdY��Q���2&��U["�b��R���҈�4�֢��l�6EmT��DV¶�lR<z����U�?����"�
l6�M�o�}�螿����m>���_p�W�?g�>����(*�Oo'������_��k��S��޾}��PUz��?b����оuT^�|PU+�S�ڿ�~�W��	J��'�=}65T_)��������z��%�S��KҿU[P��1M)�(*����?��_��['��������=|_3��>�/����S漥W��?�
��}����?�m_�?)�w����ϩ��������'��|�>׼PUi񱶯���ֽ��t������G�����c ���=�<�ޠJW�w}���\���1AY&SY\P_��_�rY��=�ݰ?���as� ��;Ϋ@                     4 9�� �                       Р o� $R��B�J@�
 �B!"�(� 
�*� �$$(�� wp
*���@�>�n�@��JM���
��#uR:5J6ȩM�;���⪺Ċwa�  � W�z:F��kx��d��:�lQpp��UGA���  ��ܥJ�UR�T���2�M��Vl��R�2��P�uEܓ6@��  ^�t(�A7�Nt2h��C!��!7!\��r�L�d����Q@�T���+��u�Q�![�:4ʆFC���:+�`r�  ����F@3㒷Ѡu��Ѥ��	�D�*ͨ���h�4hlh =� o���*�E(��.��kP��]�����@��C-P&��]ClT� x ��hz5E[�.G#AM@��#��.�U;��#@����FA��� ���|z�
QT�
�� ��@��U#�h�pN (��j��;��J�%7@:�
7c�� 7�'��U@��I�R��:b
h2�hݺ(N�R��wc��� �ݎ���  P @   @ O )J�SF&M#F	�MM ��1��� �C a�d�F�4�j��J4C##F@CA�S�*ER�       OT�Q#@       � �	�dё���F��j6�i�Or���w��./���/����[8�D,}��,y�� ����J�Q A_B��	en��EAB���̣�g��?�q�?X�@	 AW ���j&��
 �E$R��i�� P��f�[�ނ??M�}]u5�=r�3-AФ�`�ʋv�g��W�O�8M�����դP��f�̹�%��J[[5p*�X�����,_�ŭ�lVǋ(1�ml��"1ΘA�qk�G[Gd���0l�fMm֐T�n�aś�.u�n�.�g:��v���~���x%Fm�$RAfq6���h!7(h�B��ӹ[�?���%��S��3O�dX51RM�R肒0�O״�s!+]Aduf�3E�e�-ɗ�d��bڱ����� Y���~���,:��O����,kRkCNP�Ҳ�H����/|<z3�U�T�w�y�1���W��u�n�Y
��ѻ����c��qt���LC��d$Yt���J�umy�Zi��J��jь�hL0<w%UR�W��:�� �����&�f`�q��u�mQ/fҥ&�6V�zB���j��&{�	�=8��A��%l��+ɨ3P�B��7DR�S)��7MH�L7H�T6�rT�!Z�7E�We֍ek�AUS_�Yٴu-�F�G0ڴ�!�1RV���)Uo7J��f���U��b��Ó��x�s2+͖�f|�m f�韖ߞ_<���1��b]M4i:ʯA2��0'��Ŭ�ݚ����y��'��Ê�3��n���A�	UV�ۨZ�(�j��:DO0�X�kTP�	qX��{`����(2a��
�b���e�4�f�IE�t3]I[FM�f��k0�x���p^Y�ܒ�޼Ɏj���."Dn^9�C
w����k�n���qlK�eZܕP��9N�&d�r^��]UɧtP̚���8b��yn1�]��oj���)AJ�Z��\��v�V͗r�-y�ܡY�%
�xt��0@贕��BkqV`���k�w2�P�n��r�А,��ն.�{�[�Ƴb[���w��Ỳt�ۧLZ5�,cř[�AR��n�A3��͂�f����0Vf@�7oK���z]V�t(#e[�{F�Z-E��{�5f^n�UZ���p"ZڰU;�r��5���l�Qe�D�O��5���!��Ud�j�T�K5V��I�6�TR޸�F꩑p+虶s2�,�r���9SnxY��uy^L�9�-���kF��yh���;��VH�j~׶�
��$����mռK-��ٴ�2�׌h��&�z�ו�⬔1ui�X�
9M�X2�� �i3Q\J�eIY�3oc8-������$�b�P����n�]4��=�\sv&v����Z��j�@L���V�=��ʡ2��A��ZXr�8e4s/q�[T�޽�*΋� ��HZ:r2��x6R>c�Cf�а�(�2i�w�%,bOnU�#�@�,TR�ǧi�<5��m��lШ&�eh��(����P�-�i�9kb���E؇w+.+R���������t�	�n��� hQ�����Un��[�ܽԵJJ\��Į�L�rң��M�5r�,݂��H�7���ِ�u�қ��[z仩i���d�ne婗��Ӗjk��A��q=&)��$:kvBp����.Zɭ;ʱ���� ٭a�3*��,=�ܤ3(;�ܹu������D^���#Z/NK��<.�ӗ&�`�� D��;ø���1e�gt�� �R�[Kû���J��:U`��7��f�<H���V/q�-���$���X�R�=��Ѭ$-�ݹ3^��ݬqוz����U@�E�U+�b�����aSkTX�D�� Ōn��1)V]M�xvm�TVTw�0ڨ�$�Өh��fM�A�y7���[K\%����@�Ɔ����]��xAZm�t�s�6�(��}Vuἡ�&(릝Qm�n���6`5����u*��<ڥE��T�Z��P:�i+j��:Ò�+F�/Cy�Ջ[���bʘ�ǲ	���܂���Vk�-��r�70�؄YUm^��5Y��fY4�{������%�jI2�����G,�LS%����2m]m,!lƕVR�v�X���8���E��WR
u���Dr�j�.û	j�A�O*�Y�2F���Vɘ����Vir�ɛ��dc�,V�^h�kqL�����X����:K��r��d��tF����y�<�څ5-�U[��S��ʚ�L���3י*B2URW�Û��eѸq٨�U�3mU+�U�j�݊za�Ұ��x��y��q=�&�7��md�����(k،٣6�i�[�e��e�S8-�b��w��r-Y!yy�Ớ���k��,���>�r�^l��ʊ�ٛX��푻U�����l�d18�wYC�wȺ�#��y[W��.*�(�����W��h��� ��/�V�H��:�*�U��f,n����a�5kF�1�ńh���Jҽ�5���ݪhmIzB�S�H����f�-
#2�+s6�%�AV��/UX����GXv\Y��ly�@2���v���0(��1[�p�9v�<�RW�[�X�ὃ-K7[UI(�[W���ɖQ���2�i�����d�b<���v�n������p��ܼ�S&�9�U�U�V5�y�
Ѧ��3"2�w3Ǩ�:����VC����3#^�O�����6�*Q�7��ck
 u��˧��t��%i�,ɪ�����i5ˇvV�f�uL�&S�Ym�yh�!m<�z�ǘ�ڻyj��wl�0<���.^�ձ	�H�W��f]L۲��2^A4f⚞\�kFb"s	���sJ蛡��qn�Yz�SYr��f���k�5�Ƶ�6��K/=�2�'ZTV ��X��{�zŝ��p2�ޚ�B�DH�1����U���J�7u!evS[G.f=�3�z��(�{y�И�ɵ,V#ki����J�S.)YU�Э�f�]�S8k]�i�5�	��*L-���[ݨd��Tf��[v�u���C��]<[:.�ɍ *	���NVX����xa�J'�x��A��UT�HUN���DI�.��˳�+%e�W3�X�R��2��-��[mbT����UD��BZ�����(T�`�{0\���Y�ZT��D�C\�hZ�����f��ڼF��l��voVme�mګ{g0�:h\�U��ղ��jo$�4�J�͖��ҧ�)�X
�ТF��h��=�/cub��Y4�h�=��m�ZB:��Y��N^����96��r�T��͂�X(9xU���飩4ƪ�ݲ-�V��5�ݎی�ז]9	Ռkp�h$9On�)tŹr��f�����G�,尋��b�RM�	Z�Z�UhB�2�غ(ԖԸ˪&m;�Pa�Ѣ��գ^�xܽ��
٢�ai�j�k�r6oE-��XB-�j����+�(nelWa�éR��f(�k\�4&iA��F�p�ٻ�ô�m8᳕3&�2�6U��5��׳6¬�]�"�T�$�s&��Y�h�Q�e j�u��p����E�����x轣�&-�R^��{Jnx��m��n���u�f�P��-�"��VԷyVCE#���-^.��R�6/[yG0�U��R���[�An�����WL�����**��䴽3y��APӠhV=Je��uݼ���~�*��	Ur��9q�dс��Yz�:����4-Jn�.��&�xrhܥ4Q���z�MaG	�v�+oY��-TP�`��6(��ն6a�D،{X�:/Fݡ�MfQu�t�'7��6j�:�.femZ�
t�WtM�װJ	��ͱX���P�7+��+��Vq�e'\��#�q4�e������D4Ø���#_�Ɂ�����4,cv�<��x�ư�N[uf�IF[��ʷv`w��t!���5Q��iZ���i�m$0����.�<;�Me�Hdq���5zC�z�3'7i�.�e�`��ve����"�ix�p��Xr1f�7U.4a��Oh�.I:�p������2��l�^�5n���8t�4���b����yi-XR;����e����0�2�q6NR�{U���Q�����i�n��ZJv#+��gpUe�5���ܭ�ž�t�:^n[{�(�,[XU&3[
�Ҫ���na��]`�b�#rh)�Uz��ܩ�f�]ڲ�8�ڹZA��O@�x.��onb�6����r��"YA�t��(���A݁�����3M:4�I�^ޙGT֍�ZSNSf�1iN1�.�rb�Z�Ama�(R3s�	Z��9��5�M[W��	�5�e\�f�<lC�Zfk�]i�/V?'/R6B�Ul�6��PIٻB�йGe�Y�S���صfI�(�7"���l!�-�4�1�Y#�Q)[�v��Í����7Vh�f�l[��Ů�|��I8��n�W�`b0₣)]?�wuO^^������*2u������(:�rű���{(,ojUܵ��v:���Э˻z�nj%*�u(bD���9��n��`���b�R����7VE*w��\�v�ަ,
(����!��e�@�Z�� �k����Y��uy�M��j^�����1s#��D�����N�f<ηJ��9)����Ղ�4l�(��Pܥ������y�0ݑN��V�;�QX*<r��A(llW�L�#���36��;���Q"vhoI�ʣB�n�n-�ܚXՕ��)�Lr����6��6��m���ʐ�1x��H��wv2)�ԅ��J�Zl�Y�F��ʗu�.��t�]1���F�Z�J̚e)�nh�dM�g@����k�-�|Y(jLY�vUPbYE��J�{���i�&ҩIlx�U]�J�j���n�_L�\���g:�Ó���J�g��\5�c! ���:���1��Lí���ʴ���5��9,�`��v�X���J;U6�Ȯ#�s-������f`R���U���T�e��FK� c]vN���8%���XiV�39��:c�e�f��#TL� ��ˍ��%��ձІ�eB�I��J�X3���얖����kK�[G�B����ScS"���kVm�Z�-�mZ��k�-��U�բ���X�Qk�Z-kQX��5�Ѷ�bڵ���ڴkU�mh�cmEVƭQj�-E��mQm�UkF�*��b���5Zѱ�����V6ڬmQm��mE�Z��lkj-��m��ūllmZ5Q�֋[cV5�ѵj5m�mF�Q�m��Z�gg�a���v�ӟfnr��T+p;>�g)�UC3*<��VZ5��.]����Q,�hN�b�F�S�[5R8,a�c]f���9���l0e�*
���kk�)���{ue��g4fٻn��.<f�Ba+h�CVյ�r�5h~7�R�#]��Ʀ-ŕ��NR+jɶ4*�XU�UA�n�˪���1�NQYh�M �P8R�G:2n�:'hԳN���{U���&�V/�ɥ��Jƻ��z��(�
�3k*�z�9��ظ���<H�m�]�WLN��1�16��#�jK�5��W�PѺ�ɓw���65�on �3K絛�RÁ�ŋݕ��Y�3���W,퀎��Q'֬����襲��.��0��R�=b���i�j�f�v�q��f�;B�SҢ�3��=ùҨFT�(p䥁�·N�t?d�T�c��� W�S(*D�ɚo���ւ��s!8�+��5�sR��W��`Q'�P��V�
ٱC{�թZYI����卽�]�r�ܡ��e��M�F�
]Q���N,�P���Ga���|���y��)�4WW����@��mXݝ�*An�{"{�d��x����S�ں����S0�+�KL�5%׎�5��#,�ܭ��;b\z+B�`Ub�9d^u�&��f��}U�H��w�wjOA�p}Vn�3�c˃fγG��uC-c�p'�45}\�;��V�3<xH6G)�:�"I��!�k�$w(F�o*⭱vB�dYu�ʜ��Z���m���t��u�:[KK��ҶY�M��bѤv��A��S(k�Y���|�+���U��z'D��_W)K��J袷x+7�$��!�ǽ׃os�Y��3��^�����a����ok&��Vd����Ɛ�5�c����4�V<�ˏKDU_5v'<c�.��$�ݓܮ��3_sL�v8��j<,�9�cxN�r����{�A�<v.<}�.�t}�E�+��REp�L�S�����U���n�h�N��tl��Bͩ�,V�����X�T�;��C�ݼRu�3;�����۱�Bs�j�����К%I���y6�]T�T�W9v�+��P̬5ކ�BiټH0�q�Wچ�9��q9��,؞M]^��J�̮)6�Kt�vx+�v��bm%LIz�^z�UѸ1�%=�ޣ�Qz�/�{sGh���vi�{Ytj�o1N��NSv��Z[{��K����n�Ye�w	�p;B쏎o�^Z���[N�A�v����Q����3!��I���f�f\�xm�Ŧf>ѣ���d���Mv�T��\�ۦ�-PYV줅w{cb�ٸ��ˮ�y�f�����yv�鹹�h��ӕ���)�Jb��P0h�㩹U�\�<�-K6��G���k��KMge\�Q��([�m˺���9V!�;{��ם�$m������2GV�����[�X�������5�9�&��fY�eum���Ѵ��s�7v\�z=:�3v��y��-�D�ؐ0΂8����뜦e��a�]�q��.�
��zKՔt´V�3{$�����Bd�v��1mծ��8�P̋(+���uR^��38�����K�K!w(.b��WvE���G�u���MX��}���k����&�i�aCNi�U��L�6��ݫ�A옹o��cs$f�h���;&�}UO*�U�ԡ//V[��9Uţ��uz���=�e!�[5n��d�n�5k;n^j�r�Z���[�Y����˪��U����T�m�Q���i}��W���wWP�]�;f#��Z�FG��:x R�|�L�f�C.�я!��E�"�J���(v��oAb��b�vk�W	G��3���+wt��j���rUY����=���<��ߪ�2�,���]�pf��:᪾9��S�a�0L�Tt�4/�����=�-�N��{k�����nX����i�1�����}�l�HVl��c�V�_3�V��9XMA
�yd��ܼξ��I��׹��g2j���#1���h�/s-mu�wJ���U-Ü��/R!��ml��˩O(�8���ٮ&/��fK�z]��T��Z;UUf�n�`����M���dJ�VOb��M݌�n�L�''[�]����m�Š07;.��z��0>��*�=|���0R�ż��\��M�J��!cJ�f+����GR^%(�:��o+��I\o\�F
��r�z�f�]j�{)xh�cF��$�T캦̼�}���L�1UR�#��v�U,<Y�r�"�J蠾lr�*�1��;�:OS�=>�ŝ-�=a[v�un+��=�7�<DUKW-[[wmWo=�U�vi5��W]�a���Ǧ\���ڽ��<:]AV;z ���<pi�Vܽ��V�Xsz��
�2�g$x�L���LWb�ڣ�O��P]�sz�7�^l��cd/[���;��Ss:k�Ja"�*��gR;Yϲ�W�+ܕ��uҷ�H~v������4ҽ��3^5��n����̭�� �&�ǢW��w+���3&�|�ĵ�4�xQ#"������9��*	�����;=�n�YB�v���c���/3&�߲�����ɭ�	uW��O(��D�mU�fT.��#����Qs����[�#��F��/�!KY�{��Tz�*l��O���L[;����;@te�q����#-��C;-`�Y@l�&�`�1���x��)Tf�6<,jՉ�zQ�R�x7+P�Qӵ[�{Ζ$��}�xvi�Q���<��=��fF�~UZ���[J�l/������v���Ղ�h��JܼG�����ًi�OM�[�6�}��&�9V��$�IWVV�����cJ?
�
��B`��e�7�@2�mz�A�z0���
V�mpt��3r\~\�B��xp�i�֋����-�c`��_v�*�ʫ��.�e�!*Ş�mY��[u�l�*c=Unc]n^���������Ӭ!l�',Z��\㵞��`/"*�ݧ��M�5#8��M��%�hV"�U^Y�Ms�]�zz�1�� �"��;�xU���~�ee*���0�lz���!�`��MvI�</�]Uz#�փ�,����g���niLK{{ �O0�W5�\9p�����Ӆ�3x�|���B�J��0 �im.�𤝇��XkG<��1ַ���xm�T�3��<�j�Z�2���̝/���˷t.n��*�P5w��!"�;çZf�PvOL��s%�>����:@�v�Tw���6�y�ڣB<7����0� ���j�����`Lە���O<���V�R�@
�a"�=�ݬ:&v�)Y���9�AJhX�Y�LeT�V��c]���wN`��w4�R���t�E��k/��2� �wf�t�Ʉ;�l^�2�smj��n�g�Χ��2���uT�0Bܓ�	,�=xj���=�xW�wIY��_�5+o�t��p���ɀ���-x_s� �d�-]�;�^�9�d����M�i�=-��M�����uoc�0kP�F3�V�;|J��vUv�����U(w&�[Y\�͝�u|��sM^��״i��;V�B��to�S~�p�F�^U�4������h�%����<�b�E8��cZ)��/%ÝMf\\���V�$p�y�v���:�6�[̼�}u.<��pͿD&���9�sbՏ�%��779��p[�1�m�]�{�m��`�����	~�3��s�)�b�!i���X�W�N�l�@����y�&�����7K.^���b��4��U+�:�Z�/r�\阳{F; ������e�����UP�5�o6�G�
�v�fg�H�޴(���U�L�mR�Y�sd�^���o7*�f쭛��Ex�j]k���]�܌�;9��a5�es��%��l��H�$�@z2��5X.��jI-JQ�i�J+̅h��Y��y�u�|ek���"�
U�^�94��6���uɹp��:vU���5Uwmh��sA����0�
Ԩ���w)��FP���|p�t��烧�M��lh��I��2�n���8X������zh�%���E���3O6�Wyz��0+�W|�V���(z��Łl��l�ȱn�V�5R�2eR"ݪ�b��s�=�-��k�]K}�U�TC��Tr�X�$�]�Yu,3V���
8M*)�GP�v5O3Q[���28_H7��^@��[�̮�z�Rʔ9���0���Vg .R�d<�vn9u��]ޅwU�a��eɓڱ��ow\4*�eP}z�a]�䣣��9��zr�]��*�]޺�ZYu��9��ଳ7��I��a�$�eW5��0n�ë�wO�=\7l8j�l�٣V(v��6��n=�҂����w�1Օ��c����;�17B���/2��b�5]LZ����4e���.�+{O[4�+,Vޛt~��d$�J�v��w�OZ��NP�곮��.�o��,�!2r�7;��� �du�VZ_	ٹ{؃�!ˋiƫ.��Bb��Zl6��<2j(4JN�Ec4�g3+��f�p��*5y��,� �S]���ś��Ѣr�wJ��X3��/��2�fcw���q=z�b?d�y���,�wn�ad�'���ν��m!K2��w>�m�b6R�0,�f0��%��u5�X��N@dN�Cu�v_Hm*/���$s�H���R���S=z;*�9#��&7�B�d����~����ڳ�oU�vQ����k�mЛܝ7�Iז��N�4�c9o ��2i�X�y}էS3g�y��*��L�}��2���Ȟ���n�]L	�|�:V ���,�!XZy�c��t�U�Տ;���Ēw�[{���KN�㷍ݻ��ۚ�=y4�PB(���0۷}Y%��	�ܥ�Tج�u1&ua�[��ZU�6MU� ��X�P9نU����K��*���Y�v��+�����8u^)U|O�U�pʫv{t�,�.��g T^�"��H�C�'
Ο!��JC���_e��^Z�@[�u�{\���6)��F�����]�� �d,������)k:翔�I�<��6�L��:�(X�`	��[16�	q�@��(L\Ga!�f�ʭ�#l	��v�y|�0�\M�1]��լ*U%��LV�R����5cv�ٚ��$*ks�z�H,r'X�K����`mJk	�d*�7��22�CJ��������QN:Ҷƪ:\��ٝ���*e��h݉in�Y�RfmP��g!(nL�ed�Yz�&��
ҸM�9;��f�r�x�BY��΂¡73f	�U�����٦@4b��M�r�b��"��-�s-�a�i��j�t���8ݸ�R�ѐ##U��7��2[4X%��\me���,a5�j[t��[��Q9q����e�\m͊I��^a �K��SuA�M3t�h�^����e4��N̪`���с)n�1��]�V�a�mV
�l���(�ql�=�3D!�5*7J!.�Q�V;0�+D��6.�9�f�;�H�J���l��Z M�3-Bt��i��З�`6`�ѵlu��,d�fa)qf�Z�c��
&�轐Rg	�#�;]���qYM�����\�iIec`M�6�,�1e���kFn�#�Z���R[�Sm0��f�8����6ٍj�1ט�3h�6�RF�zŚC�4���J�����ؗ�u��Gr�	{cL!����\���f��F�������jK�8X�݅[H:U���ښ�[XM�C�h�%J�&.�b�$!Z:&�CJT�ݕ1K-A�h
�.�v��ٜ6�	.�W:��m��]06��p�.tU��֦Qf��K-����4p�K�;h(*�3��aq6��u�������.�+�,[6�ż�Q���Ƌt��y
�km&���8�¥!��S7����P�x�f����Sx\+ಓ(8%6�����1����Kf�Ŕ�iCM��K�b�24f+rۣ`�GK��umfkl�h��.#40fՖ�d�ʌ%{J�&;F�3Z���0��R���1��D��5�-�L�a]ͥD��9�kM;M�L��6֗9���p��22���@�l�f��[mZR���Y�"���U(mE�Κ��l5@Ŗ��Ƴgb%+4f+H��,a���eж`�FYc5
�E� �)	�����k��l�0�pѺ���3J��jQ���v�������!��Dc�ԋ��P`͂
7R�BV�8Z�4�։�+���[� ���\f1�ַ-���θ*7mW��EIM�]����b��g����������틐��ڰ�f��ι�i�M珞�E�0]��y���%�E�2!��6�%ի� ���wW�m�cZ����k3LZ�7.�&t�Y�i��y5��0����b����.��5/
#��5��fqY%5��e�qb�����f�����$��2�nS�p�Vivx�2;d�d���\A��ڶ�\�C�qtr�`�n���Y��c��U�t���WF��ke�*�)np�M,v�hkieQ�G,�:5��Ǭe�V�$îe��0�6B�M���it5ӌ�*�k\bl(�&�R-�`�&�8��In��fj�;0
u�IL��f��h�c��H��-��	�F�nl�h�2 WCmtQ1m+bgb�`�"e�#�y�K��fJ��B�Sn�XE؛%\��)SM3a�*�qp������)xmf�ir(�k���.�2��E�X��:�[m���lHL�Y���3	]uqej�f �,p�M���-�6�[ �X�JJ�ʼβ˴V`�����.f�C�&x���qP�P��]m��b5t��e��Aېɵlct]�D&2bX�{!:볘�9��5]�L���ً�mnjB�����m&ԁ�Է����!X�v6����\�c2�!��k���aT��92�P�0J�u����Xb깵Q�#y6�H㵩�.���NuƔ��-�l�W�F8B�a�4�kT���k�bC��ĥ����2�luX�&� j.
[ej���@sK�_<��J�ŨҒ��֋
�[�IJc����Ԗ�Z��.3!U��I�Q�d6�D��im4љ����u-��k
�`�u�,6�����`�a7c!wZ%j)�l�� �+���SJ�������+��2�#.r� ���	Z	bk{C�d��.Լ�(�Vm����a0��RgBJ��뉋�-
�4ks	]K(M)7gy��`Y�Q%(#5�Ϛ�7�V��R:������!lj�٤��*�[��s3VV�-�'j,��f��GC2�{mumh%�/SJ�[�صH�;Bk���-����x�j݈GMڅR	UA���Q�Mm�֠]���t��]2��+�0�����u��S��m�xŵ��ۈ�1����B�.\�Ҝ��)
�0F��Pv"M�^0� �4��`�)&��a��S�XY�	�k�V� ��e]Bb�2mo5۪�
���U	�[�+-�CJ@i��.7�j@���u�Şx�_)�Yu��!�MKJ�R��tGl��#���n�&,X�f��au�n�
	3�^.
ۂ��hq%lq��1��.�n�Bi�.862�lド�HYHL�%��3`k��`���К�h\�ZB��ȖZY���ntr�ݍ�J�dؕk�Z��ks�&ll�ձ��(Ӫ�R����Đ�CQ5�Ҧf�Jr,uj�4��yr�1(M20��Ѥ�2�N���k-Z�,v���6����D��f��b��hu���X�+���X��*�-C�Q��&5�j�X��l�Ʀ��Y�n���B��V���3q+�Qۅ�����JF<]�lac�s��1QiH]1�g0p1�Yu��cn6�IZ�!�1����s,�M�s]z����b�i�D�m%ňEnt,8�ՙeV72[K�ii������Sfڒ����A�H�V����`�4�j�^�k��܆(^� $qX��C&�4F쫝��G+s�c����k�`�5�Q���3����������1�����2��X�Tj�ɛt�5r�[�UUUUUUUUUUUUUUUU]n�G6������nIec֌{G
Uķ2�J#4Pk�VY��¬��L�c��i�q3���+n�m�3@�U�8�ua�p8ˊ�M�n�P����NR��e��.��V��2�RV�r�Tfc2���>���I��B����'�$�cѭ����u\��ו����/��U�XƴTW������釺����w��}o���/*��3^��"	��ou�E��'7LE�j+���u�%���F�J�QF`��o.E��<�e����M%|�o-��罷��Tj��������e�M1�U�I��^j�.��3wq��D|����Kh��F�Q&^v�-��h�)"��w^R��b�"fe�v���F��6��Z4��%���㹽F�F�ű�}]��҉���9ۻ]I���X{��w����>v�Y�l�n�%(sz����5�������|W(7��6��˦�^�-*�%R� f	�|Vʉ�'����,���S�m�
3B�4��X:�j,4[,�Q��k�:��c���m���̭&�umy���Ԕ����yY�-u"�#�Rk]��p2͒b:7�+��0������T�����9c�m�ĬnքC+)�֬�uv��iMDq0���[��,L��F��LE��v��Ba��K2�n{Z�LF���X�MtbG���Z��L!�� �n���D�M6"2�2ܸ�LJ����SF�����&�El� E�ǅ.n�y��X� ՛1[��#�F�ٕԙ�UԵ"���`�ɭ�;^S	�̶�667mJ#b��N�]4M�,Aj�
kXD3T�V!Kn�Hչ�qa���cQa�bS���Ź����	u�� �r2��QqxG!�v��(��M)G)(U��A͂[���V���h�9�M5�,����e�M4��%����Rښ���v*s��`�[+6��&�"���"��Ɨ�mp��%0�Xa�`n�\���IM��`VӶ�"Eԉ��B�K3SDҁX�܉��2�gLCa�\lZRE�h��ƭ�6��%J�Zd��+1t3-e6�S
�f��R!Q�l���A.�\���mXV2�.X:۝�Z:�p����)���t�1h�8�Ŗ�2�%�(2���,e*��5���-!(*���<D%�X��ʱ!�2�/
 �c��B5iZ��J[�+1e%� �bǉV�cU!@��A�'�����n�[�`��*ٮ�4fP�$f�Ͷ�ٖ[Յ痝^8���V��7�^�X#}�d��0���Ż��6�$��t̳���(�=U
���{8�	�/U��"W�T�≟oP��YL��u��sݪ5݋�d;�S�X�6&ΐM�A}a.�ҵ�&�E!-�ׂ@��$A<f��<���kW�����Z��x��)z0C/(>�v�x5�!F�Dލ��w������(���Vx��@e;΀�u�)/s���p��^i�].V/�R��l�͐�/���=���S��KplM�"��;��]另��8|��� oV�Z_.�3�D� ���Yͬ���ݻ�YU��يΚ,!���8�Ь��,NyT4� �A��2K�n��v��!
��0
��o7�Уl����5��D$އ��ѵs�j������^amk �z����qd,��*���V8�6�N��z������LIU�K���&!�~d
t(��6`�ն.FA���/1��lf�]�0�"��d�a��yv��B%�R�d�\��M+3���mkc��k`Q�������S��|�9}�3��}��/�����I���l�\Sj���Vq�!D7�>ULK	�*��͐(���A��፛oSL�BI�BpA�{Ve�yV�7DF ����4����U�����Uզ��'`�ϧY􏐧�\���T`�f��8��i��P>7k�C��Ax����>�ҡ��z�a�A,�|gLV|/��o�?��2��8lB0�VEJ*w�A��]�o`U/+�6}�6P �ֳF��ѫP�/7s�$�7yb��A ���C��Y�Tr��%�Ќ�����9C�t�#���Y��΅��}����	a���@>8�#�a�ދ"Uiq��h�8��P��lǁ�y�A��eW�2j-ͷ�̌A+�<P*���P^"R��7��W�A�&�n4��YD��c��#%�J�/S�m�$G������bv�(�d���B�!�����9���p�zmo���G-w]�����Fu^S�r�~�I��Oà�@P�ϸ����,� ����b�-�Ҽ�ݿ9���5x7f�_ӚЂ��2�Z�l�'�V>�eKha�����H�����o*k���q�4`D��lN�������xig��<uL6F���g��AĭLŁ�A����  �����Z�>�n
7���$�I���t�n,�{k̃�}i�q���`֤��!1��K(��W�u�����Di��<�Q��E ���A�@�^^>C�����^6P=a�
m�Q� �M���^��!-�а�Hj�+���϶}�=��@G�%c��R�4h�y�1ҮZu�U�$���&�7�vk��0��$K��z<㒋C�P�A\�ݖ�4L��C��$(D�c]���b+t�L]`��[cmh$�t:"	]e�P%�T�D�Y�LL��iE.n�)��،a�k�hWR�K�[3]RR �6�V�a��M����m�M
,B��'%�,�hU�\Yh�K�m�1x��m�˚m�ҡ}3�V;:�N30Hi�mP�j�4sv���.����:�Җ�	��M^�׶�����&"�`l�]
:��.��U����b �x��̋/uM� �>A����p�A���o<����Au�*�_[M�2�*TU�������K!(/&X0Y2�7�uu�G�׸��Ԁ��U7Gvm��2H���W�D�EH�CT�iM�$�D0�Z��[d�t1ci�cf����Q�	��� Q�a�M��:�#tl�3��9>)0!���mK��4(u4qn�_����H6�1�!*ojU�V�X�ق��`�Cj�jX-!L�a:ȱE7��5��*���c'��;Y(L�|m֨���B�{9�ے��.bK+����C\
����ar8P�͖�Ѻ���s@�B(|�W�n�RgoA��$!�B�&"HDB^�BcY���յ١b���:��e�V���L�F̻� ]hMv��At(�VD%�?���q�9�K�ױg�g�\�}�P �t�2ޓq��0�
�����e���!}#��U�"!���gwK �L���n�%u��ͬ�8s(�#����Ż)�hб��l���;҇+�� A�B�3�!ģ��FN߶���5o_-����w��Y�.��~^ݡW�����'C�5�	eP�O�56�bP��� �U�a���T>���Fr�l�m$Q"��q>�:o+
"����Ē���}a�ްA�Q�*�A�a��BW�JScB^�0iz�#��i�1g��g����inC�[��i��6BT�*�U֣�Ĉ�B����������^�^�,ѯR�R��=��X����+�K�I��$ɓ�����He�)XR,�O��RM*���+ٵx0n��z��Jy��DYB�R��D�e j���r��K����C
d*��E��A���a�t��@Ҹ+���Q�*�������;oSc5v��yC���>�A8F`fB8��_�� �$�fњr[M�oQ�Fk^���6���w����o�өM*��[���2��i5��[<�L�)+"b�K��k�ƍBb�2��{@�oE %U*-++��t����[b�: ���(�'�|�^�n�]n�p~�C����M��.�Yfy��dF�/��>��B�Z�B���Ӓ��c3� �^HW��5-�׈"!/D �
 �(\b��#M�&O����}cg�	�@4�,j�V�S�0��A��LA�|�C�5c��iY��,�G��1s�,e�k��)ZeuTA�A	A�0U��a�w�|�G.�>-���A�K�h0JK	��ނ̱�X��>�y}w�w�6/�z(:u��e�7y��{��f��ljL<�*p@^�mԼ��`�U�����(��:��M��	hgƜ�x{fZ���E��$�j���B��M��Kgq�<̥���X�d&s�&�B2�p#	�ViRƮ���tH�l/j�X�6��a6l��a85�qx�V��c%
�Tu�-2�-ܳ"h2�)�dS�ز��ˇ9�p��V�\j"P[s.�]�vv�>�~-K, @b�eQ1x�c5��Wl��B.��{����xh��&"e-���F�Y��
e�G�BΚ����Ղ#�8�-e�^ݯ"1]��G_-��˫�@�+l[T}�,[�@g-ذQ�9�7WY�n�c�c��4-�X�00����B�м-�j�k�dJ�cv1��i����tަ��@�uTZ�� �N݆�XCjQP�%+����5ڧb
a�h�K�ػF�kW�B�Ax�`�c��K���V�@�%a���$�2��u&����hKՕyg3\>�Q�F�
 #V@��>��n̶8��/�yY=$�@�/A�K �3)���R�
և��eR��c1B]��&K]��dʌGϸ U`�H<�}>�V@�t�4y$>��|�qC8E԰���K����>�4#�b\a��a��K]L޲@�/A�-��`�p�on]^E��4֦ ��2|��2Q���6� "��A��������6�߬E����R��^V��L�I혴�Z.p�1:ٲcF�La�|>[(E:V��Z��'-n�����-_�tη�-mM(k�+K�4/��ݢ�>�~���{�Rv�n�3jȸ�i);���E�(Zx�RYx����S7W���#Y�2&4��[���I�����!? /�2<4��W�<�iVn��WuJ��V�f⦉�b2mu�ӱ.OVY��-�k��;�g��o�36�-����J���w��E�b���E�X��ڪR�.�����]i+T.����v�ii9���l�0���-���k�X7yܢmb�
[u�|�v�6w*�oK��+sv�t�x�ѽ��գ+��^mrj�B^L�VP�%d���Λ��^�4&���y�ҕ�L�|"	E:�u(����껹�ΡnS�
5T͹w{e�$��^Zs��p�n�Rw�$�i��B�Yg,�j��F��6��*Ø;[6+P�&��i�H��a�}(�ֳ�[6�bY"���?ۻ�M�2��=�bnok�B�c{uOx���K�H�V���x�upB���ϣz��vU����~!�*�C��Y��*�7ˠb�
�f��]rk���v�^�$ݛ�ݻÐ�H��{�mʗ.�똆BeYN��W��rb^�^U�kUv�5�J�욬҅f����%I�Ϯ)�&�ɖ
�!�z�Hl�T��n���P��9��CgD%y9x��˃&��~�=��5�r�ɣTj!0[�/w���UsE���-��sr��(Ѩ�[�͊+�p(�.c[��{���j��*��uΣ۪�~��^wusn}nm��Z�-=�,y]s�{��(�A��6��̖�7#|]$�r.���X�ɋ;��bƹk�Ҳh�,h���&��ѱ�J7���ȃ|\�6-S�g}q��w��;� ����m �lF��#h����E�D6����JA�ֿi��xx�k��"Bbc��f�f^�q�h&�8�����@�"q���Z�]6��1`$��h���@н�C�
�� � ����<<0���VE��68�9�tv����X�&b%Dze � ��M�U�����r�l��]0��hU^;�b�*^^��Z"ځ؈�z@1�q�T�|�v�cq��x@�D��ŷ��I��k�"M��%�#����b-��5փE��7b��xa��u ,�x ܟ�̫�ƻ�o�
�f"b b H�3���rj �cM�h���j"i�Z#��P19[|ъ�k�ɹ���FTM����{��D{�����(È�D���H"%-�Z\f�tB��8���q�x <O�@��T�!�2n�F>��_g��%�#oXt�Xtȇ�Q$�[�O�N���&���P�(I�Ē��ς�mC#1��R�n6w�U�~��w�/_��QUtt! �J$�t�'0(�Y[W0��*;mayfs�X�m�1%�;��uD����$C1���nP����Uz��s6��S����A����m��a-r���;�3l�*@�v�����`�[8�Y�y#=��H�FT�iX�[:��j�f/F�|����w['�' �a�hס��t�ql��7/5�"��7�'`�f���~a	C�T�l�1������1.�[R ����Mj�bٯtsɊ���R�0'�ƥL"&���آO@���éI���[���K�4��2\�hp�Zdt]@��̮`R�k-R�#�\��,�,�ݔ6t�<���v�LS�A�������u�i���
�͎IQ���qd��By���2:YX#�чb��`����ʮ\������e.�X9�Ch����mq\�321tS;���DTCeM�T��+vo7򽎧{�vj�6p�UT�.�g,ݩM�(b��ѽ/WS�Eu�*���-.#��Q�7U1'
�vT��s=�����(��A��eW8����k��@�h�[r�l�o��|�oی�Ƈ3M�R-����ݬ�����́�!IW���9b�����f(�AŒ�؄�9%��j�Pki�s�����|���;��+c�Vl;L����_5���S8�iʛ���2�wu���V���c;B�a%��+�Z���j��g\�������z����tb��W)}�y�)ҡ��U�.�����$�GK�(��\o./b*ސ�()��+�(�uQ���CU�4�w��jq�+6�2
�N.����(#U(�2�o�ק~e&�(��U�z�r�m^fWB~��̭����ʯ,�M	`�Rh���s�jX�-�,�(�&��?]d��7A�iy�<=��-����|nԾf4^Î�T�����44���r�Vܵ{��*ޯp�ƺ�K�ӻ_��Ёt���c�mJ� ��N?:��X����ݜ�����d�<z�T_+�v3z�F5%	H��9}�fJY�y�Rk�}�ʁ�� ��a�����S��l�$�]@��;ӣ�|��]J��Y��X��a��V�mz�	������p��m�ʎ ��2��.UYX�E �3�rɐwv��7��5�H���m�G��;wn�L���M�a��C[ےq�"���i���l�}��R)�R�ZxxB!��'�m��5��3�{4Q�7����2%l�%�������b+"6-۬�s��X~�������g(E_�}�.�<�{HN��Z�[ήM��J�˛�FS�[�NHE��j&� ��xy��A> ���"P��H��Λ�^�[ӌ�7$��۾�>�33F9�������]O�'��v��ˮ�9��˱�k��]�O>��>^��{�S�ﱸ�_Sֵ����qX�3�5-v����"ٳ�1�M�\W�����d��R>�B?0w��C��髓�L��>~�9*0��.&��B!�jf���w��c��W�Cm�d�D��y<��V�^N���&���2�Ł� ���o$B7��k+ī<�e�/ɣȧ�U�����^�7i�^gdN6SK�Ô��w3-��tW����"d��]˴Bi�����ci��
\e���u�VĖ��j�
��mA�-a�t��j�bib�M��J����'i��a+F���!r`����)��9hXi�Mxd,�z����ڢ�m�%[�����Nl��8v�;mo�=?7�� ����n��-[q�F7�û:��6T��𤳹DgE�ؚwݝ�%���Fe��nq0��Y��k����Ѥ^=M§�n�S�F����њa��v�(ؖ�Q 1���թ�8�����"���Zn�gZY�asWˣoN��>٣�Ѵ鶩��w�"��.e�L7V��d�e��͌m�<68=;=�b�n�C�?:~�߳١l�ivbl�B�1fX.p��X�Q������H�x���.��6�������c���d~��;����uK�E�<�LF;)�%��l��3_ak��=Ӷ�
���_^�����
	#�{޻���/�)�����|�*����$�7�P����S�9��#q��yU1.��J�r̈́ˢ�xG��w�wYػ�b�V�6Wmǉ���A@X�a1.��=F�-���B9f�/��<=���@I+�co�aW����bZ�N)i���5�ԷM���V�V�Q�}��Y7ӻ�g}}�5qk4�hҚ�f�B|��Y��{ZLʓ�|��*��`���W����A��k��t\��%�_�X�ݣ��_2����ӧ�aζ$�TF�ȧ���Eȼ(on�m�woq\�:k.�t8��\o4urȫ�![pWh|<=b��Uw-�~y�W �%k4����;u�p��W�v�O�0��p��n"�~z�;��qaJ1�;��� j]�*���s�r�{e�D��~���b/֕I�ț����fE�v)Xkc�΍H�R1�������s��p�P櫆��6_.�v�ɜ=���n��&f\�UM�=R�{��w��v�S�rj�;��2b2fn��"�]����w-��/Z&�B���-8�L�3d!�N�H�Zw�Z��;V��}�\���Z*ט��>�%lٸ�h��<F:P�%���蒟u�U�zL�nTK��_x{�r��^��XuK
0"��F~y�;E���=���Y��c��W[�A'����;UҐ^,'�ՂffU�$c �L�h�G&ť���;��q��!y�����}��\�.t�)[p������fٖ��[=N�0��嵜9z���i��jgzו��!*��0*Xj�b��	�f���)�:�Z�`��� Dpʁ&e���(� �C�=�F_J��V D1���|�fB>6���;���sd�n5���kg�΢*TB#������� �5�Ŗ!a5��Q�K��YH�H�w�_'��t��~�#�>�b��Q�	u<�=�,t�d��r�3u:����f�́a�l#Or9�2N�އz�ee��^�Ɏ�Z;2�CϤ�Z�f��.��_K���ݕq*���m�œw��sfv���˿-xE;��Ǿ6�e�r�Ut� m_]gF֞Ύw^u�a-iu%������N��{ݙ�X%��b�6�H�j�qP�K�ʼm����Qts��t[~�j�ɡԆ�y*�ݍή̡��Z�$����yY��B�TA�{�`���9vh�m���zU���޽�E��n��#3P�깴��)vQ��H��f���<��+%��Z��i�nݚwuօ��,��M�u�8v�:�y��U���đ2������̙��/�(v��2ݨ��n3â�)��kqM�U[4��`s�s��d9T��������:�e��g�2�af�!���qӳU[y=7GT�ػ�x/h���6v��=�v-�����lmR�Vqgm��]�k�6��s֔slA�����v�Ҕ�m�=���7��Oy���x����Ch�����fYh36�<�p?}���D��8��	b�%%�����k�-�7���("�T�o.b �����yzP�[���`�d2�廮�wn��]�ᤉ�Q�n[��F�2Ywt�4j0Q_=�Rl��;�r�$Z5�|W��1��ۆ��~�y��gu�l�RB�ܷ��w3��N�"c��	.�-��a<�'�dDHk{ï���a�����o�B�t�Nm�7b��5��il6t#v��f]eJ�B���u���ۜa��n��	\\]Ue.�.Ps��E�F���]�܃p��Њ�i+[N�4@�ٰK�l��l�l �:6:Y��)�M5�&K(k�%�60@�*�G��KӠ�l�N�L��X-0@l3K(��J�.Ʒ(�U[�l�\T�)F%^!mIhPR]av6]����Ҹ�<@��t��X�/���Y����"it���7[��g�;;9�W7T�֎c2���e�.[��&-�0A�it�l-�J��&�)c4j�e�A��@�fH�m�%�+�2)�
:�6�� ���2: mU�[ЋYCK1a,h�C/6����<e^cC9t.��4J�5�d�6F��i�6�Ōֈ�"6X����eG^����֏��:,`m�İ��9�Û�49I	 ��C,�B�ƺ�+���X�%E��j�ݒi�rbQ��e�ڹ��D�h�t6��b]�L\���h����ŹW%�c���j�EP�	��U4�Z]���F-�)qo;`��T��e�`�X���]T�(ZpCi^r�V!R�m��L�إL�\3&U6�Pp��6v�*��0fa�G4u�].i\f�!Va�!�r���B�!|ܡ��5�\�p7jK���::]Mt�q�gS:�!eA-�u��)I�]n+�(�MR�1����Mp�`���x��v�6������,�U�+aK����.�6`As�e�����J �Q�e.0��+r�Z��=����K��iWL�54P ��X��.�8E˿�ʿO[�`@"!�{�[�8V:�y{{Wz*�n$�S�;@��g;���ɸE��?Nt�<:q��H�W��A�#�Yl��D;��w;�R���ؚ�V�����"�h�X�Q�"��U=����_	��"�x�Fo�>ԌC:Dr�Ю�Cö�ŕʱ�/��7ҧ<6qD̀�By������2vӕ�z�P̼��Ձb]�Ͳl�Z�t��c���G��?A�y��#�xۻ�͖��^�������q�;g�2�3�Z��5�������_�_�\���]�v�h.k[�L���r�7ծ�^`��l��pFذ�W����|��݇��_�q�
p���B��~�AA�D��((�ٓ6��hv��;[-�q7��z!�?'"�b"���MM�[Ni���ȽV�[�U�j@��8� "�TA��3/ٵя�Fp��`��PxL���:�F����n8#6�rڑy�(c5i��r���ۃWxa�%��ݽ��Ͼ��1bl6�*#ZO��nh�x�kzˎ޹~�u/z=5����>��t̍ZWͱ�8���4������Yn~_���s�{��m�����yJ�\m����
Ɯ�K�4���'xy۶-���Έwp�2�:��-�b�1��B���z����v1{윾l���v �Ι�4��zj����U���>��y��S��"���!/�!�rpێ��������L��.�,���"���q�h���Ś�8�i=��w7Y�L��R4�%Lv���4ƥ�+P���$��z��a�;����dJ�,�z�d�=�u:.�oeӺ��T_;�Xqv��tgF1�� ����gh˘Gl�0���K�T �j����;k3)�mcN[8t1G����Ҏhҏ_Zv��"�<<�5���� Dg�G�g=S�b>O�on�u|׷�� w�al��h�B����l��5f��тfY��%���L�ɮ�pP1f.�'}�7!�����Mwmev�躮�}�gsz��&T��f��s)wo�R��V��]�>�q�#������(�S��kJW�۪qL�zff���T;G3E���w}��oC�M&��ƞ�wG��A�����wS|:�M]L�M�eI�e�끏n����/��[���(����䗚�z�	+G2��i{;�v���TV$ql< ���]���w�.�	�[���'g����ն@Ѭ$�Y2uP@����< ���H�l���+Mǀ�d�I�$���q�58��Lk2`�"�B��G��i�k�l�1�a5)a�\��f�ėb��]���We�ٓ6h�&�	PѤ[f&�f�k8,�ka���r��ц)h��6�q��˶/;�{*��1MլB�&fh�m�tTt�;��w�)�LʙA3�l�ם��q��in��[{�	��ޓ"�:͑��n흛�ڥws{�U!�)c��N�}Wm�q���Y*�b��{�5
!C�dn�EE6NAc�\]��i���;��> �'XI�o5�FC�@I�D̊����w���ڥw}Yޫ^�����fB�|�緬�<�!c����X��X��+q,Eei�s)L�%�v�F?��T�gt�`���`q�n2�r���V�ت�!����AUR��gh��3�(RRYQ��=#�W<���^��y�P{nu+n�Xn�������RL���of�8��|s���*X<��{���S^��8�^�C�umw{�m5}R��kx��3-�c՜m�}��؄�fި��?^�����'g��cd�P�PDD�Z��B�{=�؎§��}���ӭ���3I���&wZ�a�2��J��Ia�@K���v)��d71�C�\;���q������o�׻P��U��])�W9��;J�Kؑh�`;Utk��ws	 vEm�E����%����q�~�U;x��J��Km��x`s�c�y�M[ĳ8��|}t(���Ѯ&f]-ALF_9���*r�K}�G�������U���o���m]�ʮ��-t�#{.�^�F���1���;�r�P����zv4��7CN��;�6Hꦻ�P̛��I�v���R�eU@EW6[=L��{z8!-eFUB��`V�F8!�t���עdj7��*�����ǳ���b�z}S�{A�a�q��;Ք�)1�o�]s�Wn�D��2��N�gu�{v�{���ߛ�<�'��Z���;�"τt���~�����ͯ\�"���vv36��6A9���U�l@���W�mT�^Y�����_R,m�C�*J�(뤪�<��� 	G>�y���'�o�(<|����4��dk�����]�ꪦ ����)1�w�%�(��������\M\�6ZE��E&z�u���!=UVU�ƣ/U�l��������n�I�#��~��nd�05 2Y������fm�¸Q���dΔ�-�w?a�$�=���S���~��^��l&�dw[ג�.3��̪��31�n���'�z���Fm�ah:e��Ո{*��e�ɜ��M��j��K��n'g�r�����4���xp�7ag�S��q�R�~��(a'`���c#*���T]�C�k4�y��46����0S7��+g�N�:Iw��-�߂-q��6]��#�[X9��Cka5vv�m�1	W���d��5�����H��g.���K�30�[��di��v�!lm�G3$���4�T	�
���1�=e�帋�J.�m�֘��sx�*t�X\�\�j�>}���!ٖh�e��j$�Ћ*�b�fD�9v����>$m��m�6��f&���{�سǫk�~t٨�I,.dA���:(�/v��>}���VZ��[a,�g۹(�6�i_��K���ih��Cn�O��d�z�p9H�n�����I��S=�����1uoS��2�X��k�wuW�fZ�.���v��񕋾�B]m�]�n����X���ʶ�g�$1�`m��-5�f��
]v��ow�η�w;��;���O��uG,�,R�qg&�f��X��^�0~uB��׮d��\���%	��:i}x]OcI�_2�\<�31T����Xp���x �����Ǝڶ�躿�8e��aT	��l�+>�Bf��3,�"s3i�\��xi>N�A���h��D�8�������k���h�sۊ[h�ʟT�vOFf��J��e��M�7v�l��_Vvb�3,&{��'3���U��ϳQ�u=�T���8�u]\&;���"�L���"���H�*�oLu���O����m��þ��7�uz1P*����p����^���*���#if|��Y�
�i��/z����/��~�����R�1���j���-Dm���ݭ�ۍur��ͣ��u�H��[{���Hˠo��"����[2�s�f�U\˸T�Ql��D���E��H�rR�+ދ����9v[�v8�R��3]�B�"Aue1�3E�sĴ�oI�C�i]-w�*"�z�US�XS�wnde��ۮ�j%}	�sӲ���#�gsH3n��e�|����e�b�2 x��1�\iZ��ڝ���r�x�z��36��}ļ!օ�����Ӫ���EF�����%�h��of2�m�h���b��=p��'s;y��d�qY�/�̮W��=����=�,sZ�v.��ie��3kX2�����E����I���+�n~1��P�ݛF��ss^%sӄ��pצ���e�ޛD����6�Uݔ)mU9�5ǩa�����;R}�� ��r�:0�q��ۺWzu�7-���wooQ�L�9[Xv�y�ud\&�a)��?mJ��H��*�a�������I��� �	��׽�H�B�;���ι�����]���HDF`cO��&]����f�I�H)1R���������
>�)~ˆ~W���$��g���s�n�_�v{���m�$ ���xDR��LI�/S�n�啲^8�M	m:6���1��r��.u}��`�u�HE�L��������W^���]_���p�I).�_��{i���=������z)�%��U|#;o��ݯf, �X���3���ۛk�[س��*.[��3�
��d����U�k�bI�3�[���-2�Zme.թH�;���GU3Ҿ���ȕS�W��KX�8��{9~O���ߌ�����刌h�����[)z2's[ &���u���컁U^X�����ӭ�8�!�)
�a$UVtx�7T �V��ݸ������5;u{v��B�c��j�^���#5|�l�W\�u,��f�CG{[���8��ɈkXf��e�iC�7�����_?N��\�K�Q<Ƥ���o&���5L�8�b�Wtӕi��`�C�����X�X���cn5� X�vd��<����_���z�Z��z^V��m��(T��&#H�1��
�~���A%�L�9��U�����_�7��#U����[��|�v���8o\�N��c.f�}��'��ݫn�t�Wq�n��_geo6�͎��o��k�h���3�Ji8U�g<�}�^�S�=[�F����fq�r��!"�e��ܥ����gFiy����]<�I���V��b�v�2a]��c5�iz��V����$��-n�xf���xT��v��փ����Sa%r7��,u����(ݦ�W.[mY���Cv�e��*��a� �+�ʘ(�7ЬB��ܙ5�kk[v5�h�Rm1����L�je�7P��6k-�us��M=�>�yC��1)�˭��A94��O�w��}��T���ͼ�:��.���&L�l�lP�:\�h��;|*6�`n���sd�TlNS�Úm��V>���w}���J�?�^���K�VD]��N/C�T�<�#/z&�̎eC����!�.w{xKW��	"'7t�e��w[33H����-���k��d�|���A
�7�ݧ����I����m�X�X�ٍ��h��B�ˑ]m������r�B6�z3!�u��G��nqEz#�
��1]���e5��в��e�r�z+�
�9u����޾t��n؝&*�b���zs���ș讼n���[������v�ek�ǏI�Z�e����Kc�����Z�0�B�L�y��7�
an<G��׸��rw�>��y��B�Z���T�Hݱw*:k����p�����DR9O4Kjz�Z�N�d[�O���i�mºh)SD%R�w��w�}�r;H0�R�@����Ǫ����g����b"�Dv8�^�����,�C����n�<͎�������U>$�۴�^����ƘRDF�O�!�WDHtJn>�����Ώ��S���ʇ�\s�2qu�Xe�w �����N����W�Hl�eS���w�c�*�9ٳ���#�m��U7^��%��t�k�{��ٸ��bOzL�2݇SAG<��C���ܘ��̇Y������������e%�8��8�1KmGM�&�eڥ�o���[߇|�}��l�UX2���C��]۴dL�hM2Ǵ��fۨ;���y=9�2�[�<^�q����	�팊l��3���'�݈\s�*�3�ɝ��v���,�S��}Rp���=m-h��D�t:��M��>f�J�N��C���k`2^,t�.��WoZFZ�kkj�`�{�{͵{���Uv4�}�>�3�ͻ5A
Z��$�mCm�Wp�����d!Uv/k5�1����=}��V.���b���ᓖt��rY��g����gb���D�ٻ�VJ*��8Npmڮ�DL���ҧ�*N�	}��~�8v���R�ܪyUa	vf���u�!������i^�7^N��dI3�M�M�)�}|SU�:���^uB���vvr�GZ�d�QyHf)1��zџY|�kUh������#ٹ�	"��gg��!�K�]��.U�k�����y�ҵ>��'��A��j�����U�������F���R�C�c�BT�º��Wj�����-��2�s�4�&� \��1R�فx����;^uɁ�,IfØ[�(�4T�h������v�]��т]6��Ǜx��r�s�Y�,�٠�#�K�{����F-B�4̣��vij�G,�I�vd���+��(L�ޘ�m�~��O:"b�S����ej�����"�ي�E�̮ݻ��f�l�/K�oUv�ӏݱ���u��	n��S�W�����9z=�y��^�}U�h���)�!�2�����`2���M�6S��N��Y�wl�YO/٦�
gԀ��stT��V_[e��{�i"f ��2���}O��!N���]HmddL&C:t�x.�b�>���=�^e�1��An��X����̨�T��ԥ�f�KQ�Ó�0��Ʀ��DW� ��ݖ�:���m�1���Í.��ڙ��H$��#+��E���)��'|.�
f����9Ct�d.Y��	�n
�x��Q85��p�S3/2�����.��6g�;2���me���o�<��>���E�|T�B����^��ѷ;z�)��'E���ld5���z�wL^ᮩ���S񁤻(��h�ЫCT�KnEtq�|����]i��|�z"����Ө�ƻ�����:��'	�Ge��V��%��¯���f�}鑨�k��>r�����0��2f���.��mV�B��Y2����c�Ř�a+1�e�e����
�6��Y�b�i{aV*�>���7�;z�Oy<*���lm݋8�L�ݪ�ǝ�U����X��k:��ӧ؋�ԭ��91��i4ʻ�er�]����f����􆎰�z�����D��ԅ4v�mqff�h�6�������<g}��d�seDud�k��v�Whq�
�	�6�L��݃�]����fE�d"��+�j�A�4�_5�h��6mډ33P�*�y���s�k4Ey{g��K�zn�q��t�.�n��̧U}x�QY�޼�W��<cCj�e�?&���L,5�v{fYD�:=,�ؔ�(0���;s�b��ͅK��k�m>2j���+�[��˂9��M�4l5h��y��#���_q��ߚ{�O��C����a�%ji�;`��J�M��'�������Z���f�n��V��5��k3'��N&kN��U��ۣf率�c�'}7�s.���dVc���d��m��v����lG`�j�q�^jTER���v�����:!�7�43t���&7[f3y�(>�3�χ�D׽���;���@9�s��O��k��?���N��z��X���h���%t&]��&n�K�R\������<�`
@/��C��6��uX����p��W�Q�s�H�t�2���pb�b��U4��$W��x2�V���\-^RŻ�:��dW+�F]x������(�
>�w`�gP�x\�����7�uS�q��twJbXj	7�K����R!D��	�72��=�u�S�Q�*̎�:��56Ǔ�4<��Tض/E��������WPM�:��I�˲���L�匍�Nбݹ����Zj_;�
���g��2��+�Y��R���^aS#��U�#�eu���{/2Kޥ8��9���C2�)��8�guX�c���uY�]�n����FWUv�M�3�;
��Y�o��1r�s//0�O=�{�I���ݪ6q�u�z����Q�xv�s7*�^�̕Y(�<u�c����:]��c4vj�n��3S�PC^=�ʧ	Ux;#A*{[�gfa�wj!�ɮ��M��G:z��a�����{ܮ�9J��q��.���!������~�KU��M��d��_>�,c�[-�׆��R��HmQ�]˹0b�>ͽ����x�m+"�ܬ��";��D�4��fE��7M�ȏ3�,#�k�xn%M�{��
�w��(��cs��]�l����wAc0��+%��,"$��o��X�-��ƾ����sO���I5�ɋcTT�vܐ�I~"�߇��bk���&�ES��>7_{��/�&'pHo����V^S[���o]YgQ�N�p1�X`[4���Bcn����.M̗4�@�/)�dab��,��֒3E-��f�����l<к����ka���3j�J�J:;�5�C
[�D.�C\�s�	���刓g~˳�m
����Z�l�s�At]���q6�5�M+`�H6�
����,�Yq�F�]�CR�^�����\$,��l�"W�	Hbj��,�����@Ί]�q��12�梮��-Ĺe� "4�ж:�/V�x��*�[�[0�ƴ���� X�I��q�f�Ѷ�P0ql�F(�B��ؓ!��["�Ү���Z����A��e��h����к�Sj�m��sl3il1���l5[���	Dj�����eE��6њ�%]0[��4�H��XX�K�5�]�`^S]���$DX&�����"�]��ɜXu�a�
A������օq+s�YR�T��Җpe��J9n��$ڈ@˲��tu��[���]X����W�cdb]u��5,�*��VD�am��iu�M6o)���E�`5v��u�qHh$L�� e��Kc�����-�
�vw6z�v���K4yS5���ڶ��	u�^j��;mjd]��۳���r���(�&��U+1�(�`ꦚܱ�Eت������_ͦ���;���Q� �q��^�/[���f]�nl�Z�v�(6Ù���2�ƹ���W\<��ibi�Ր�C7�l3M۴%U�1I����WYS[��x��u2Y]��а-JE%�i���k�[[�����1�������$f�p뀩t5�]�p�˲	��:)��=����laƝ��*4L�ּ�N�ck7�U`�|{>i^t�d�)hқu=��۪xU��p�B�����q�����-�5�3�D�Ef��e��������K�a3����~�n�P&�t�T�1�����١-��%zq�?�_
�z˃�bv��I��ȼs�S��|#��Y�SO��ۜ"���Xa��+�[u��ɥ����;2vI3���[D&�J�3)���k#_J�ѓtH���g�s2p� O��P�ϼ�e��*2�r�8�u;��v�G�Q�_�]�R����ÓuF��uTO��MO�![�O��x���ٰԱ�ܲ����;3������W^:�ۡ��~'VJ�槜�T��ޙD="d����v��V{&��7h-���מ��ѓ{t��ot�Okww�(�X�~�lc�y�NjhX�WeW:���DD:����Ҍ~��-�r���܏
m[R6`�C��u��O����'���/�x�Sݚ碧���^��g`�Y�	�:m���T3��)�~���f��OT�><�dOet�]ٝ[����<%�X7�4CDFz��.Ԥ]1�A���·�d�
�����Ƀ6��5�V|�}�r��q�a�f�$7�ϻ�u�5*ת�>�R~�j"�_nF�����4���V��"b7-�<l��JŰ���]�R�b"c�a&"ˍ1�lU��r}��}+��D�����k�����#6�'.�f-h�*�4�Mak��e3Wyv�jeO?�]�L��v�f�d��u�m�?P��m�P������ީ��;��Dt��γm3��M?�m����߳(7��wS�Yӓ���\�N�$��f^���YhA��w�8ϭ�|З�q����\=lf�zf$<���z�%u�BB�A�w��:gr���˺F,��3OA�䪖F��.�:���y�RZ��5C��&�����l��N���A�Nhk���grTə3J���@�ki����3L �w.�w��oL�L�0�׃�[�γg+���aq��iL�E�v/W4�{�v󎴉bM��]y��uw�/��0*u� FKY[BN��[���Cp�Ϲ�\�	}�TsL�53Jg�۽�&��3(���w���~�lѺ��a�ڮ�e�Uʙ�US�%���j����m��w�5]!B��Uf��/;�(�R=/�w΍FE5m�����M�h�v��۹}G����ĝ�EC
8%�(��bP����(��-����r���C0�����n�6�
Gk���G^CWC���l�C���˹R+Rݮ�0J�\X�J�ݵZq�F�6�����KZՉ�ne���(�Tل�Z�lĎ���;�
]����^Gh�:���8�:e��}�~���b8�A�uT *m���N�oN�6��d���E��n�l��Y���i�ޯ��$��	�~�����%e�O������wo�ո�T�+|�]U30g4z�v5p�jzY�̌ ��[��`R��'�)����B�{�S`��W����~���1�ġz��]�j^2��d4Bpm{�X��X�wÆ��3;!h��Mܛ��n��v���0`�a�:"�r���JΉtS���]���$��˼���hYvE퉂h�ފ
e4�`�hG�ݑ�s\�s�%hut���P˙��f_p�W;���Ǖ�>��on�m��RUV��H����G�[�g����.~��Z������]��:~���*ey�w\�µDّ��k#C^/�����Z���A�N� �R�A��]�B�S[�ƭN;�_�Cf)1	�f��̳�e��9g�:*�a� !��Hw�m���N�mC�[���t)�::�c,v���|�oy�O']{w��Z�5��5w
�V�:�b�q�2��טl�����ʇ�&�
�ΎO�f�F�I�ü�M"�JL�J�\n���]����|kD�x�v�`�$+�A��6Iy�I���n�)9=�������]���E_���Ϊ��4*�芖W}5�Pz'�j|���ї�2��hޱ��n���#�(k�=U0���� GMN?a|��}�oz�ʈ!�&�]1�[Nŧ����!	M/�y��!�%��fKy]��w���݇�rY�,I��wY��i�[����x��۶\��z�EBfwB�K�B�q�Փ���I����Γ��W3�;fWL��dlCj�S��>Y|��| �:У2�B���o/�4�xiT�aT��7����F��e-Y��f%��5Fj������{%�n	�3��y�e6AvMvN3�?5ޘ��3Ȇ�L�5}�"%&˩X�1���Ѹcf8�����w��|�����O�ms�5D�93��k֦홚����?6!zF�־茣w��=�Sm���&P�G��6��k��ey �
�Ė��uz8�uQ̪����O�[��fR�.�2�[B��;��-V3ž�0�j1|��X2K��Wz�>���� �y���#h��q�CX��@�,������3S�*��"g"�5�i"��%�0]h|Q�=�=��]�y�rhJl.b�5Hsŗ������.�x�sl�d��*�I&V�F��[���h��u��،fWZm�[���?;��[�o����P[+w2��B�%&���X�:���M,݊I���Ե 9Õ���N�4��������G�[4��xA�M�!nHFPbf�5���F��a��O�������6�����v�Tꘚ���.����v�̳f?��������?:��meڮ�-t4F�-\�wh��}�"��JA3܉�}/���^y����\֔�c�����v�Wo��Rޫm��g+�R�r����V�]OU�ų}���,�tV :V�=�.��[�
NuWF���f^��}�5k)���y�q��1\�z�Pw�꧙dv����78����Y�Ј���N�U��YyQ�1�e�ʬ�c�%��Mi�n%�3Au�5��d���q��>��U a�m�O��4�jT>Ȩ�§�R�XG�ډey&^v��{�Xu���������,F�O�=�!��I`��Ihs�6�;�x�8�4�z9�g�5���Y.�����mמ\۝��	�2��������v���-�{� ���/N�?�P2�Q�V�� e��P��2�t�=�MT=��ǧ\e�NO������w,֚*�ҽ�Օ�)x�a%L�.�e���
[�u���˸�R�����J��ItS��f�>�Qނe^�c���j�\�io9ͫ[ѓJ�{b�©"�+�]���Z�Wi���_+�i������c��,@WЇL��`��8L����<�xs��6��=(BVE�nut��7˞n������r����QLV#�ºn��]u�~wW״f�����y��j��J�_}��dpcǢo�[��u��/:���.f���S�YX%m�n�
<�]���Ʊp���v��^yjT�kL$�T�ѱog.���D�>�$���oh:�b���&�sn���l[�5��7,�a4���hޢC���q#%]ٽ��V&-����&�>�c�h-Ju�<38����҆��ke�X�������پ���4�Ef]Ly�W9百��_��G�:e�S'^���Qv�������Φr`�u�pHNeq���q:��:��M=�VqM��m��9�Ψ�޽+I	��f�z_K���UJ��dZQ����1�vlCb�C�{]��:�V�XbU��s�p�ygE�Wr,�\.u�k�WP�c��0j��c�����)%5��]��僕ֳd)v�#V�c�		bF_�Ѭx��̭���t?5d�:ke��K�b䱍�L_3�6��2TY$BI��=�I�o�\��6�W�ۖ���r��%%�+��������o9���j��
�>�Q��5�m�\�渕6��,j��}��I�s�E��5�^V�X��j/�\ܺZ�m�o1��W
���-�5z�ۻ��[�ͷ���X�ϯ*�ȵ�A��\ڠ@�D�T�?a�xʹ��W�\^_ߙm��'�
�U8�7��'�:C&�]
-�A��qs��S䔅w;�Y�̉MP�i��5Xm͊���*Պ�b�l��v��+��b�,la�"!�������hYn���a�6mR[^W4�~������9��U�&�ݕם����{iK=W��b�Xw��E��n����{�N;�Cm��緪��}Z���<�8u��y��mU,"5�y��A��V��`�Z��!?V�ް��w�w�I�Url�y�Z����&�6�m��&��`�\-\_#�3*[�a�6��[�c �fXK+��˛�(�a��I������Ɩ���"��,�����I���(7�Y�����[��.�e�	%���ݰչzϷ:6��뉞|-�f��xy��?s�[hϬt��k�aCau�Ke�����}��=��^J�	��ݶF����«"�k2x�[k���qQ�74���-�x`����gDLM�̆��¥�T�T�U���F|ۛY"o]��L��֮�L������U� �D^7�w�c"/WG��@�U��j�5����߄ܻd��z�a36݄��1��k�����@l쿦kp�X0�g��;4ŝ�K���lʥR\s+MV���������n��y�LYD#���Mu��=<P���r¯"C&��g3n��bKCn�룠�Y��1,\�TR�h%�A[Q
�(�hQT3v��:��*jKʰ�f��0*Xkp劖�
�[���Ŗ�m3WB,l��).b������暉�r�l.�t��w�����$uv&�`���ڕ�Yl��e^Y�����D{%%H����r����k3S_�EK)~^��!�^}N�d��˜���z�Sn����F��5��R��-6���$���|�*��ı�u��_F�-�b���fN�=w0�v�g�ed>��������O3���R(L�^��n혢�V�;m�t=ehF��S��ƵDY22x�o2!��(Jf�65��16���˲g!�b����J"��*�3�m��O2�����֪�n�.��A�v:��G�ZH����j���z8�L̬7O&w�/�	J����.����WS��^�H��TN/�-xh(߮Ĉ�Mv�D̺��T��a�T�7p��Dt̨CL��:ػ���N�m�������l|[uT�,Yn���G��](�o1f��
d)��hnN�꺝���fN��U�6�o�3K�q�!k	�#�j�ed��V�F�x�wf�u��ox�'ȉ�&�����D}4WѺ�r~��Ʒ����H�	ؗ�4�v�)����nL�3[�����L 2�ۗ�Z��cv��̻����������m��TQO�c	̾�}Ž�DG�8�wRt;("��kr��Qy������dfЭ�Q��]�#����IR]����o��O�]f�n��;��zY�[�WV��	���ʀµ���xm��z���Z�rr�.��m̬ks�}��C�f/g!1�l�>`��2�=An�f����kH�`�`�M�I8!�L�a��P���N5�R��7vL�eVܱ8�.b�c���b5&�v%�P�z�U��wqsp���ڸ� K�"�_�·u|C!���:�.D�D�Y�z��ﳗ�Dʸ�"�6(��������̓;Y7���f;#to˛F�.�Y��f4yfs�l�Q����d���묐��rqj�'D�mG��6���F����/9��B6"�o��j�R���v>�[�f���28���������y�o��	Y;���L+M,���<Y�L�v>�������<y����,�\��OA�"�q�`���B�5U;�YCDD�oQCwXc���Z{d�Vuc�^�3����bi�tK
nf���BC�]����z�器�}�>���x��b�n���Y�vA�n����� �M�ֻ`��-�L�����,��1<��vL�f�*�r��&eJ(�H;9b8�'�bi�C�X,�)�2��]��Q��V��zEqk.t��GXu�d�v�L�� y��� �Йp�M.�˓�)v�P��c{55%�2��)�U��]P��rÌE˭lf������4ѹ��f%F�%�R�y�\��z��n.��3(]5v�X�f��׶�dЬ��jEU.e�����}���-��&�aC7X�P�m�\�����v,���c��2��p^�5�4�����^ɞ��˺W�+�����j_e�⿾S��>�����.z�X��B��a�����_N��)�&sͦ0n�D�&�e��TMAzu��y��Ѭ*j쓘���$��D%��Ư�F(��w��l��v�D0�����0Kjz�:��~qs MmКf��;6��v1��l��k9Ϟt^�~|����_ӷ}��x���]�{�H����Zܶl�Ƴ6١j��f���:4�Z�|�36��*�6s��كS�W��:ͤo��������~�hQf>��51��!��d)e�bV�Zے�|"5�yy�����3Y�Q���U�N�Lă(zfP!���b�����8���߄�}�{�x�O,?��d�.�~�n��-�߾&Lf��������A�>Z�$C�h.��hED�V�c'gt�C���%�0��fX��*s�cu��Udԭ�]���y*��G��o�s��WF��+9��7{�:k>���m����(K�fHj�
p ��mC(m��by�un�_V[��9ӻ�����z�ӵ_պ�[�k)�)����q�"���[����S���霪�V��%��p,ը�����l�����@�ۃ�+lf��,!y�4̱��{,�^��se �"sqc�˽�PDB���Z�7wn�Z*r�U�%�I�I��E��K����U�Qf9Sc���0�Be3뭛]�M��7�#g�y2��d�zj�`+4��"8�߷W�����fs_}����ݶ�iǪ�}^���eLo&~����\~I�YO���G�PIz�%�nsuu<�i�U��qt���v>��� �7S;ol���ƿ����v���)ayj���Q��dT��;��Y`��U'��8o�<�_�S7�e�Ҙ��&�����[��5�w_t�S��
��ۑ�slA�p�I���;��(�ff�J3F�4�v�{{�� b)$����:U;�W��Le,T�"�.�]r�˺3l��A�T�6�s��N�4�ԘG&�h�ғ�e���qp��d��Ϳ�t���3i��*��2NV��5�ջorj���ʽ}x�'���=U��L*�R;p�r[u��0�r��޾�k��i�Ŵ�k��<.lu��t��IK@5�2�Ql��9�su������g�|&��$W�bstr�qUC4&k�[��Qf����/�^ۭ���y狚/�Ż�
k)M�X�$2�<�UhQD�+
k�ʞkY�������7.1�J�`�8�	�A�^F�`�|�������Ϭ�c��D��/��cx�{�)ySd�;Sef9Wz����u��W.�����ޚ@ɤJ�ն���/ ΋9�[ckN]_^������
��y�sT7��#�u�@�K�����S�U]\�hxҜ�
ǂS���U��ً2dv�'���i�×�7�;���K���/�}�-!/DH����8����{h�=OOZov�<��hf��m�n�w>��j���ONӛ
V��$A�5JeC�Gc7W�3������[�z�݌��n�+�^]�]m�Úve�]�q8�X�7GdU��V9eYF��by�5�����*��y� 죻��O\��g[��+[�u,�P�|�����#A`Y�q	q5�L#e3���Hw>y��=�{����<;�h���Y��Mf�]���iD��m�K��zb�n���1�yF�`�nV�����ʍ˚�k͍xs�\�lk��h�Ɵ:��Dc���;�*9�pY�cQ��\�Qr�ssi�h�+b�7u�nh��o�W�];���M��W��m��|V��(�܊���FKr۽�\7��v�������nk�9�s��u�����5�\����]��W5o-��ݯ,cV��W��lZu��6��yl�[8��p\�K6X�`��.Yf.�iX���q1�3��C]sNv��@���m�v�,V��e6����\����0���U&,.4+nr6�t��+s�Xj�1H����js2�ف�B:0�����5P��6��b��	IL�BcX�Դ�cP�+��`�	���o2��JH�.\�[�7#���3ca�ؖ�	n�������.���5�K�a2�B�u��(�`�7��ĭ��c�]��a��DM���d��CV�E�6��@�D�Z:d�,l�{.��YXs4n�\��W�5�z�RەE-l[Y�rEJ����ŕ��a��j��
ĸܡf�tV���,�+��V�c�T#T�!+L�[�*�Ѹр�v5��j�SgxK�%��i0M�<u�p͓�s���(��0�[a."r(%K��u�Y��Ͱ��Va�5�����Lۭ�	\nVˬui�����X���Ke48��^a9�1��ed�&E&��f�7W�h�k���KL`��ܡB�-2��cT�)p�6\��u��[U�%�n�,���\���L�vsЛ �%+S;Yrj�� �p�m�����c�"�e��Z�]@�Q,#M�ps.�p�p�ev�iR�l�r�!��\W7*���Z����r�f2�5�fcbl����r����y5\E
�Q�
̺9H!�rD�X)6uU��bie����0Qh�k��,j�ח,� %�ɴ����sk��bb��I�JS;cF�����]J������7�<���ki��s�.��J`��l]K�:
ݕr�,=}�:��:3�l��lBTj��v,��O���3)�\D�]�Cn>,���gH7f|�X��/7e�A���Z���U�h7L�rb�t©ܫ�1yb#Z���6���|d���-�δ�dh�c9����}��f`I���=�0�s�,��"��n���ϴs%��15�­��H�M7����[U�%�-���t�>f?�s���(������z��'�� !n�q��&�H���sEes�ff����}<��\뮮�n�s`��[,6������@C�e=T�S%�{��j�Leuh��9�9<'\��� ��a��=�
��I:s�r[2\2!�=����� ��I��5��t��A�ŵ"*eԟ��C�E�_;����?�w�v���*J:Ю�m��謠ذ�`M�އ�����<���YV�vW��w]���=[M��\-O���{!'�zӯ������R�"d���qfrvT��Z�"�>ggNAI�2E)��Qq���o��{=V̿�K��^)j���Ӱ�ro۸.c��0P��O$��Я�fM)�$bg���z��ՇNεRy�gzhD�~4���|���^������1�w�9�v�,e#���S}oՎ)��e�k��ǲ��S"�"�˂]�� ����g._g�oW�j��^떝�Z���Bȁ�7����w2�� ,l��"r2HS5��m
1�"�L�ك���,��ڋ���Gb��*2�A׌�yt'HssD�]B5'�¢0�v�Kf�3�aL�:ͻ����i����~�Y燤=Ss�Dtv���V��w��zO��Ռ.׬������{_3�y�s��L�{#��`Nj�&^��5W���a�W�An��h����>�s~Z{Vz���8f���� A�R�%�0(U ݑ���#Z����PDO/5SN.n�dGOt� ������l�9�!��NL�)/�;�g2�D�=��ʺ�
9�v�Yqt$-�P�{���Ѵ���,�}�`�z��k�D��ze8��"��E ��~�϶���p���W��l�7k�$��ҕ��/,.�U~�$Re�␅6
�-�m2A�笃�)m& �0cE��]|{�zc8f��^�Yfx���#�~R^�NC���pj�����RC�0e�iv�l�IFj�*�F�u����x�&�$��ty�m��!C����/f�Vh��0 ֯If[�e����v�Z�%!�6D);FWfq枙��\Cx�W���ks>	�1�B�z��� ���Q"=!�yP��[�=�@�\A�`�H+)���@��:=�Ɛ��O�(��F��2�xBq��+3x��7�I�0��ո����nR���v}D2oP�ߒt3|�VR�۩��W+�(��8*�d�[jl���f&I�n*��b�M�H�:�w
J�m��d�jl�dh%��c]coR��v�+�P�Q��&!�kBbӚ0t��1h�1���5!6�-��+)c�5ڒ˨:
ܪ�ʹ��z/�`�`�1-.]�صk�]1��ҰՄir�Ϥ�_i�T�^��wc��]9�q�p2�3F5�.�P�m/5S�e	z^ǎ�/[��ŴIҁ�;�{�����9�w�{�@�"ۋ��M]��ϹT� ��?!i0,T�&q�L6� up0'^e�"�������:��_}�PD�+�3)���J053�!�h�����C[Z-�#3_�
���p��L���Fc7��pv=L��RorHp1k��m	[S3�������	��8�T��H<�2ͣ����D��$����<뺎������tm�_��`޺^k@L�?�X'�:��3�'��Q��_%��3X �R��n�*���]usO�-��x�f�Ѷ-uwU���p�-���%��oU\>w�����/-1��� �z�}�8�x��k�nm��f��de�p�"�*�s\�֡��~�`Ҵ��l�� A�3�&eD5�E�GcWuu�9�u
:@�C��L�HL��#%�;+|D�Dn�U!A�Guk�D�t�$��>GSV[ݕ9�=��έ�~2�`�a��e����l9���{��,�*3���R�A�ˆ����[�@a+i�Y�"��&�,�?:TK&�X���JciS�bϽ�Ⱦ�5�zH*Cmu�]�7y�tY������$^("H�AT0 �!���\S4��Â5ׯ��$ �8`�&��bg�^� �0`dԾ�v2����ڕ5�C~��EF��J�"�8<��>�ׇ�P���娳��B�dn���YZ�Z��3tE1�ei|��q�Nz��T�ȼ9��9�gͅ��!Ȫ�;��0o+�l"��b�A�oIr3)��;���ẸN�C�,++�j��2��̦ �!3v�,��g���3Fڸމ��<�S�`�2|��W��;�PY-���dp�BN�!���m��cÀ,�r$�o�`L�"�2�j�%ff����b�L�0Я�KĈAx��oT�\�s��M�W���!͟ �Y���5c���@�!*-�81ɕr��=����`�}��ƌ"�n�Ϩ7a�AĹ͜鸙��մ�q���4�$T��	�e�4�b
1���i�j����l�y�q���j`C��7ۅ������w����[�w�����
1�c%�a��V&��	8Q�R���V��4�1�?�?��f�ߛ�|�ey�Y�&L��l Q�L�Q���s�p��޳�3��V6�{��y�ց�b�vx��y{��w� �����Ĺ��	-��s-���v\M�G�}���/��T��`�mGu�ڞ�>���F>}�0k���uD7^d?� �xe0�J��R	N]ӛ�͜/P����
!����-�����>�*�(02Q�ʭڞ(�ia�QVu�4f?8&�DM�,�
��
RbЫ��un��X�J�"������'j;{� ����v���J ��x�z�m^`|h�B^h̧V��zhڑ|;y��������#���"����R`�a��������g�̝C��8���e��z�+jU��d�4V
*����u��u]�/g�A�ӫ*S�:蘕��Fi���M�4p~��˶�H��̚�n֡�6!�tRX�-j.�C�i-ՍF+�����]tJ��I�َ6�c�1h�c�� �&�ԫ�KD������L�k��:Y�Yme�ˎ�vöv�߿����2Bf�KYa ��J��k71�~��;!y��1��&e3U��~�<ם���;Tr�: �c����-���^sV��Nr� LP��KQj�D�Gs��3��/�*���n�^Ԑ#a��Hm!�"��T��#�9ǝ�����v6C,�{�3��2��v�`������T�͎���� D.z���ys^w`GY���ƺʈ�~�&�1��]�"�y�[EWA�y�3�5Js��Gk��Ʊy��1����3�BV&U�=�X~��y칊K7J��`¦j)t�v�?o���ae�5���6�����e|/x0!�lHqӥo�.�s/����^�-�7�u�vn8l��2�S]�����7.��܂��Ae6dԨ��4a.ID�x����	�M����?s^p���,AlƩKp�l2>���_�U����W����Ja^Ucz���_�s
��l ε���� ��zM�wx�O�f�n�����["t���u|/x7����ev>�V�o�-Qb	�L{����F7U_m�x,���G>��;y��8B<f�sT�Dhb��U�|C��謪mS%�cBT,�ѱ�.wY���z�+�״:�IwdICZ�S6��;�������j���}�޹n�S{�@ �����`L��\1/��,�/5�������'W��3.�y� ��8:���{.�޲hx��Y�Y���X˽�^��C�"}���གྷy��3�of-���V3��WYYe��@���Ih�� ���,�uR50�.�I�m��=$]��E����3#8�9[b���O	��ѣ��Ѯ�D�R�����㫻[Xy��м1F]�ikOR�E���i�5Ozf+�Ε�_U����_�r�Z��z��t�m����}�X��˺x�µ��g��.j�I�rD�����O�Y�S�ˎ�I%e��^T�|<�9��¥R՛/a��]��U�q�4��9�� �M��#���'x:Dn����@¶C�*0��];2��Den]Iֲq��rJ��x0_aO��>4�j�u�4{�	ʷ7;0��:o��Q�4,n��h�Sc|��Y�UA����4����J�����4C�R5�<jB�qݶ1��6��%�Òv�G��v��,�{�.���yq�7/+��n�l%n����s��劇+N)��v�%e՚N��b[�����gQ��m��u����[�Ι�<I-��O��S�Ǭ0C䎷��X3��Rf�U��/wC��+>�8G�U����-�GK\�h�S��w�����y�{�����o��W/�d�+Fьj�o6��[��S����W9��[�co#k�s�UҨּ��^m�U��5r����	-�mך6�����5�Ov�z[E��ʒ�Z�h5�.\���5��lw�د5�r�z����}�[�ֹGվ{���E7�  '� "�Cf��;y¯�7��A�w�|[�!��	t�x�N���"��m�2���/9���c�k��j�^c@�nְy���D D��*��ʪ�f��Ac=N��~N����"��l�T��Wh]��=���nǌ��bȂ���m`p�]�Tv,���%�9;1r	Fes��W�xu�
�*lT!��@> �1zH+���W�k�3� B��^q��"�gWW<Gl&�gX1�͎q��ށ-��{u���B ���2�a(sL�i�a��#�[S�ᚽ���Wy����P�2Q��u��X�ޢ��I���Xs�u��`N;�é��P�D�\�ѫ������Z�f!�ܵ�	م��;z�.�&�d^�k���������1B��T�T�@B���s�:M+"����]v�D}�@�^�C��� ʡn4�׀�w���bR$��w%L�H��mL�\�6�g�Am��W���T7{X����$E���������o�d�2����~u�,�Z�Rg�m3xu�
�oi����%D���t�9>��+h0ޙA?��1͝ˈn�<oS:ف0��EeXy�ƻޥ�W� .�g�9�����2�7�7���Lh�_O\�e0�]5<3�u�x���/t������;�;�i���\�xX~��ל*�X'�(����!P�Aa��&�j�vh�ͭK�����~����|�9eը�<��n}�	G��t/�B�L���w}|'v�����z��d��R���Dڶ�Q��I��e��WF�\��ʹ��qhᄖ
��(K�XP.�f�^H�
,7R�QŔ���ң6cIaqJ��6��d�L�i�"�u9�B�M`�ښ�r&ׄ��f��#i����Wgm��ߖD��b�[İ�b�:�[(%Е˳b�~G��hb`G��f����{��ݲxs.zw�[2��t��g;b�kB�����<�C<��yĠ��E��t��ou�("&n��&]z����զ �7����	�Ws��C՚9�Fn���s��>^)E<2��D�AJ>��m�N� �Gu��!�
1ϻ�k���ki����nq3M�|gjv޳>.�]�b�uqjP�s�͚�/Fj�z�D��-�����tNlﯻ߿�FW�Ҹ"&K,��+���%Z�go͓��Y��>_/D1�Oo�kn���1�:�x*p37]��,�u��� �Nr��ޡZҘ��K^\Þz�xQB�H�X�]��eL~����'{�q��m(�gTηt�q �����ߗ��"6F���r��I�X�Z���/;�$0��Zp��`� =�	���^�CL���ۓ1}̹�E��^�\I2�"ey�X6*>Q:�E�o��z�8Q���5��&��o���?@��B�2�~:��6�Q~AkX*׬�3V�_�Lٌ+�Wv\3v��X��L�V� �(�¶nt�V�nE�2���������4Y���t��g~k�FB^�`R`E��Mf%�<3��F�k�6X������p*�y�Z�5/_����lո4�X֪nV#w��h��t��L�"�7/Ӧ��j��o\�0�,�L�����A�/��jӺڃ�dL�\[;C��vf�VڠM�� ����(0Q��~��	2�r�'��9׷,���s��Ex6��VP �ݤ1��xx����J�B�I�����7M����K����_$�Df �������W+��zL;�Y��G`�S���g�᳚2W�� �0c2�$tg1�Ě�g$Sm�'�u����iJ�(]t�Z-����'x�Ї���"eze�[�7nY������]ʣE^�oE�� !5����7~�L\��-h���h��7P�s�PDL���Ԟ�$����(Q>�6��ݍʆ�(�>P�
Oi�1W�g8l��o-Lį0��yi)]�s��=v�,��LD�����{�,��x��{:p�Uj�����Z�R��\i]��C}��3f�&�q�g�Λ�v������Y���� Ť�C	L� !Kzem?ft��1Y�����4n-<sW��� �ݽT��v�4#�	G�y�RXb���E�`!�M��p��b�V<�W���'�fU��1��ᱛ��a�����r;{1zH�(b��J���(F�,�n��o7�[���=���p��jטN0�Tc����NP��[_�H�A�x�!��7�R`t�	<��	����p���dzQ����Ʃ�>�Tnu�W6���7Ɗ�*����]�:/�o��3ؐ>����:n���
�G�J� �"�F2�@�0�a3�{Z�m-ۇ�ox�*#'�fVXt��f!��y��m�B���݉�҅�kTI��9�M�la���[I��u�hm3��u��c�i<�>��K�:�w�y�Ͳ�Pi�Q��P��L��8jL�Eܷ<�bڀ�L��E��3Z�����)�A��h	��`�T)���mvS\ڒ��m�e�����F�U��8�6��.a45��0ᅚn]s4�
�a�����Ui�}z����Il%�5o.��As-��&u�*}���O�}�X�̦"HT'r�^o�kp�Xc.y���֧{�H����`����P�%X ��ǳ	�FJ>�MS�CZ;xt��8�DS�W%�*�o	v
P�v��b�&]�fXm�kw`���̦�ym�<p��� �7����u���'����5D�oeࠉ!o�Z�;�8m��n�g}���;�c3�O��ڲݱe���]�&��V\X��7�5ˈDE2'��J^�����f	'I>������\!mpK2����m�?	�_���HY�y��u������{�sr5&�5` �0cܘ�j��n��4p�E��O�z2z�ʥ��E�7h��v,�c[��j˽��*Ǝ��;w�"h����7�n ��՗�޻�ǹ��ډ��=�4m�`A�LA�˼9��:E��S�j(d&"�2Qj�٫�fvs��5?^�����
\�")n�v��h5�nEx����V�$�3a
�U�ekeD�n൓��%1�,sf�e�A��Ї�;=�]gA��SG��f�1n����kA㺘�(ER�ze�����߿������cXM\̱f��C[��N�⚱W�>�t�������M^�j~�=�5�f�uԠ�ZE�$I��LA���8�0�$7��`æ���sԿv"�D�'Grs�>X����wC��A��L2�mլf���M���LY��0���L�jf�FV�øUJ�����
�B�����&U�M2j2O�٨�X��s�;���"�+�2��ڋ���g�s{	�A�����	�M��C�7xt��<B!�;�5�C����%� j��5I��DL�p���1�<mU{�VN�waD��xX"��8X@�V�z�D�Oj���)�^�w=��U�`�\���,ۋ7�pt�1Gk�|ߙ�����j��R ���V��sF���`�a�I;��T��QoU0�?���;���o�l�v�\�u�Gw���5.!D�3IN��o� Z:���2u�n�[H��/~�K������.�ͯl!r��"�".М�%�H�A^0`k��9�q����8ަ"�;�"�R�ݑ�Q�XP�Qn칵!d��5��V��Bcŀ�����c���(���;l%�����-(	�fMΞ��Lp�,���z{�n�l���}�m�LA�7I����W�g���<%-�?.�PI������� ���3�&ߧ�ϳs��,���v�!��4T��l�]�x��p㯑��̪ ���9�O�Ž�������Mi}�`զ ��6��F�ѹ�of� �e�_F}O���؛��-
��^>�Wd����4*;�.�l�GUÆJ��,������oj�W�
��L����s˷L�b&f��I��@4@�[�A�bp�`A���R|�Φݷl��ǞT��sF�7�V���"�z�	���	BO�"Q�	�'k�3Yeexs�)l���0��PB�P���o�C����vzIC*�����vZ�N)�7%��F2_d��p�y��fL�aө�Z�Jr��M�n�麽zU���j0@��f��:�w3+Yv��Ѝ�������=GzwJ�[�/f̴0:����^'�V�S�t�]�R���q�z��5���)����'q��g,�&�B�+�c��yh�����or̻�fvΕj���{*m+�n3���+�lCC6�� f�5ŵܬUE�cjl�i�
��c��_���f�/���WlG���vH��Z��I�W[YOr�mWM�̮��eb(�N��Q��[]y��媓t=Q��&�F��_S��sa͏.Q��t=W���z�jX�3�h>�w=45������ιբ�l�酻�@��]�.�	��.�L���\3e�{�/2^�7jU����^q��,�79oJT��p�R�,�e�k6��e����ǃ���R�.S,�7XӪh��Y˜�|�M�3�o�,�.��]e�*LD�O/ic�;��{��ih�E���LU�2�u墜W�Q΂ȣ���k��uF%���T�� ��k	�1v�z����нi����z�wz,öh#�����~{��r��y\�ض��y��5�k~�r���o6�6��ss�cyF6���Zܭ�|���\�9[�W*q*%��+h�(Z#PCh��^TE������k����V�k����-o+\���nj������V�כ[�6�[�����N�`8;�����2ZY��,����:��ʼ\J� V9�<�u٪·UŋYm�
gR������lj�1�3)������׮���sE-�-Ѻ@��M+�6%	i,���KG&V�1v������hh�\��n�n�I@(Ũ��Cl����$Qa�I�����\�B!�J��f)a3D�n�1�3XvhQ�l)h�+Y����Y�I��lk��I�E�ƙ�  ��k�r�J�1���M�Yo��(y-Zˢ�l&"@�.�.�l=b]Yh��&e�4����\!�4&�B���%�,��YJ�S��.����ʺ.�E��q���ƔѶ7sB�S"Q)�!ٶĔ;m��ٛu)���]��ݓk.��2!.&�V�;0.�5h7����f%��g���4�*��u*���b6�[�Xdµ+�U��F��(�UI�����\�9l�Z�lZ��H���Z,˸�R5��K�F�6�e��`C5b�֫.��/]��]�lA�C��t��k�\ +t3 J�ؙ����hm5IYlR���\bU�,��*���,�KR�lô�X�JQыm�n#B�-f\Ƃ�].�h��-��f�j�M!�iKxeXCX�s�@�p�7L�"�]�h��nUUUUV2��5��ى�m��Ƭ�]�̹��R.Gm�I�<ۊ[�`2��@i�.mQ)��Lhh�QM���c�8˂-u�. ���ga��\֌-��%u*�.S�e P˭"im�: ۋn�グȻ�׀�73����n-�
�&Ҩ7����aasTsu�`����)b[h[���.s�09k4	��2�\g������(֢�}����L+&��4w?]���0l���m|@��㺘�%�ª؁N���8���{�^a|��1���Wn"WS5
��bԆ����¥�LD���z��f)jh��7�wSD����2��T`�{s�Ӎ-}��>�f$�ER��۶[=;w��{H*)Iv4�8�&� ��1���7k�H	�z�y]�Gj"o5v:��݇�>�LFR��4P>�Q���θ����y�}#�X&�Z2ѱ%�m�\ܼ��Tur$�?���e��Y��ͳ��#h��Ԛ3x�����c������^i��G�j8ቕ2��r[MNGT���3�V7�2m��{����B��D>bFئ���	�g��eD^*~��kg�ۭ|���G�V½�#�[3�J���/��G�\�`NJb�2��;2Ǝ�0�mQ�sl� ����[h�T���F�Nچ��wS A�מ�*#��h�C�{4(<VB���o�b$�}2�2�$�ꪏN�B�P���Y�==u���x�QM��R�
B��(�g�L��o�Y�K=s+)j��ڜl*�%j�e�q6������������0l��8��8�V/T�Y�4Ը���.Aeu j[�@����ng��&�p�\^�(h��7P�se,ESp�*ݩ��^�8A �I^e�|[�L��������Ʃ�*fL��gӔ���e��G^�+g�zu}�|�O��Vwn�Kw�%�����U��2k%�r��3�)������wh0��3j�4��`�3,+z�eB��Kp����\J��)�e	�N*���rVl�Av޻SUNQװE�,+;��vp����Ŏ4��v�R܏[1��s5����!�{:f��\:m�BRƺ$�p6�GG;��~�-����X�^�q���<Vu^��~�������S�Y��2�ek��	�^������uZ���w/���{���LK�U=�@ojà�:E%��"�Kb.vd=���óX8u1R��o.ŇD�>�yoJ�������04}��O]n��讹��� _�v�4�SyѫɋrؓyS_lt3�:ݐ��R
�mf�R��s�Х4���N��`���e'�/:N^S$	���r�اz�	���c�ܻx��Izq܃���}2�j�t�L��n/#��b����6��HZ���%�#/gC��߃O�����7����)����}��3k�ir�b���`�mF= W��p���&D>@�)ˮչ�;'s�!6�2�!��dX�
<�u{5zH�&X7�Tx:@N�N���3>��-��Ӌ��n!²���4�jB�9��$�!�P�6������՝�vh�C�b`F��7l�#v��a��3 �t�2ޓxr��2��=	�U^g3�MWG�8�%"&W�J���M���N_��ư����pq��ͮ��٣Cu��}q�r����&�l�R�x ӱ�~t�%��k���O}v�R`���F�M� �V6#xe�l��8t ��`%mֹآUٖ�	�U1u�jX��e#�ÀA���c@Ⱥ��fHm���V:�J��eb`��KXk�Q6��l�����7����7l�<���G8�:C�y�o�l-�jE��CFcS���F��Iӿ�������d06R��2���;��x��^ʞ��PGR��ꥎ
h9��a�����z� A����e%p�ó�����LFϚߏ���C3��yB�I�^i�h��s[��@;L����_F�0 ��2���aw���T!O�17�0�F[�`ި�Vغ3yuq�^�Ö��5�IG���-��`A��`�̭i�/&E�tʝĶtvp���\	
���b�a�q1eò/8���X���fQ��j\�	���-�.�uD�Y��	{NC��󑤚�Bw��oGMG?�6��Q��$���L�cZ�kA
f�v���v�:5�0l�9!�<�).Іb��0h�U��is����+�y�ŝ6u�c���N�Ɍ�k4z���^��64��.{�;G� ����y���`�a�z2��ES3)�r���>�N��4w%���s��o$ D���������1�F[奎ڭ��]ѱQ��7�K����<֝�4�;���!��`M��&l-�Aڪ�1�<��n}�=g�&�1(02Q2��.�[k`[�mHe!i2�;kKZM��\J�+"�lL������$3@r�/I�M�mó��0��M2���e ��Ax��L�pd������ٙ^�e��Y\��b�cF�0����E.H]���'O>q����;9��Q�����!�|�_X�lmTJ@�TU�MV�˼͟�J�]�g���=fu�]��l�}	��?���Z�Q�z������8рA2Q�X���ig�#�[��+�҅ �b�h��6�����7Gf?ul��/�п}P�>���$�e�����'�����Y�w�*:xn���X��	�1Ph����Fz�ț�Lǈ@�@�lA���*M��Z՛6/�8��pU!�E��3�r(Vb�}��{�X���ijwVA�yqeJ7DȺ^�*�~�jO2(��<l��=����٣k�"3�}(S!U�?G�R���j�qv��䚥���-ﲧ���Fjx���03)�2�0���֋�;O��iE�7�Pm�#s���� ��L�N��M��e�I{�ibV��K ��u���M�!���W��Ƭ�FuIO���X�W�jӻ�0!2u�0��2�$a�'�U�KsF�r�$�2�bXotuf�z��Za�sj�� H˂9F$q�8���u�U�#h��1ߜ~7��w�N|�A5J���޿V����Z-¥ȠD�rW���a���9�Y;.C���݃H�^�C@��|��h�>�Z��af��kk��u��(Ib�ud2L�����ٝ�8��CY
��L,ق9��Q]�/�δGk8Q�e0�˼8�=Ƨ��0���"#$�a�LOUd�v;pn��ʲ4�!�?�S�$m�R,H��nѦP�/����� h�>!ܠ�_.�yLP�6�uv�g1ZV��]�S�����*�m�����\S�ͪQ"�c2Tmȹ(��lٔ��||x|J�6��C:Xs��LCJ+fh͘� �ax�QqP���5]�Qj���$��.a-��5#�cR�6I���"�%W�e�[�kqbT���7J��WY[1���$h	��n�vY��hlds�s����z�+��S:�t��]V��7j�)\���g���$�׽�4��H2��	vu�f����yO�M+�@�޿X݃���6����Bm��?{���(��o}\*tf�5��Z�\�%S�yHh@�޼C�qh/T���awQ�&x����9��>�`��@�fT;����on�OW�۽4ʲ�w����R�A�M͂�9_f��om&V�AF�<��7��a����4�2j/j=���x�GWSO�oq�#�1�^���S��4��f�\��$ҶD R��B����	������cS(��^�B̋��F�^�A�:�)B��D��%ߡ�퐺y�u(<kv�KSl��R�m��v�_V�Vŵ�>+�����m�ӛ�6<c@��o9�[�4x�v��%^��(q�	�A��&]�x��}#I&i����BQ���^`l��������}7Y5:��w��@Q��e1PZ(I���0=���"J������'3yh�3��ɼF�`�һ��O��R���Xh��&��U	z�CW�"]	Yd��W�:6��f��d"*��"e����N���Vv�'@E RT���J��ø��e�f�g���������Od�۾��yѻ��N� ��D\ �iz��B�A��^k��uoe�t��4��Ej�}�xt>�^��3��n|�O)^]��"�Cu��["�a�h��cn7ƻ7��!u��_;k�u{A+���i˨9Hq�.��K��[�W�1��v}��m�4�;���N����aݔ���hd��T��XR�{�I��_�za��l�ť+��i,�3Yz�ȧ.\�e�\�ε��10��\�w�O����Y۬�0ت�`������O��_]W]��ֻf*-ܵ2�%]z����F����f!���{.�������Tc�gw;�+h�j&�$���Es��bmu�x(E�T��nY���-2��h�������7��w�ӆ������V�?n�ͪ�6�wI{.Tɸ7��Ю��t�� �7��u��-ؤ��s����.���Ÿ]ttԕ�4v��Q�;�$�حt���	zsv�t���Y�[�Vwvٔ�[��t�n��D��K�Ąt%���z���u�����<e�펛Ԙ8�N�.��TU׭�U�UD�������v'���Á^��	r0�u�e����͕T7������Wg���\�A꾝;�~���Ռ��"��;8�!��-hQ���_9�E�I�%QV-F�j��U���w�oѵ�6�*���r�cj涼ս)�Z�sb!x+�!QV�1E�Z�y��|mE�ck}�����DlF��U�k���}꾫_}R� �!kP� b �7�^)x2�$DY	D�s�uƒ[:mZ�6y�3���A&W�P�%14��
�׬���np�^kUs��`O�u�8'#����5M.��ey�( D�g4�s^{�
V�oh�� �.t:����R�7Qjԃd���R@�׉�5X��P��m��З4*qmT���m�}��?Kݟ�g��O^y�$Z
n���s_g��Q�!�iDJ��ݍ0��*�:lp��?��Y�=���W��jy���0���L�v_�G�
�����,�P� D�/�K�&u3Z�5U������&�u�:������xn��=��Sg��"�ъ҃.���lێ�\����8j��:�#�ۮRi�TI�
��;F��!��_l�)�Ɲ�WPY;1@��ư�^�A�QDҟ��B���F�e����Vg(�h�������������ZٓLO
�q"�XE;�-q b�C�[I������{��J��,�1, b��;�9�3�Suv>V&� DS
����]�|a��	�C��wk��� ��EZ�9�=�6�㶘eD˿��O>`���T(�e]Ш�p�B���C[�G����=6О\@�^�RD����M���U�]����[�&\7��`� t��-à� ����w�3:M_�4Y¼}����0p�?��0�S8;6�}��˕�p>��g��i"�9�DU0o�Ԓ�$�$g�F��S4]'ƫ�7bq�;�a�3�!���ʎ[UD�9\;6ڨ�⡄�ߊS�<�dm��5 ��I/,7�x���!�2k�Ca�V�:jm��X�Qtق���3��W][�4 #���桔j������ih��
v�[���	ZU���fU��GcAh�kt������N�3�@n�,ѻJ��2��l�:*h�-�u�h9���K>Og5Ѧk�ZB�b�L�g)�2�Qg��Y�x�K���Ϡ� �z�͑Ԩ�&wR�0�Q���`�ة��\�-�G�d��^���^�RCc�	�{���6u��dt�n�Ǡ�$֮���U�!�!x�&#1{��n��IXD#�}�Y��aZ�~z�3F�7��$	��aLOF����f���p���(�eF�E�ٝ�Ѣ��:C�ht��zE��`m��i�A�ȭ�̕B���`�E۪ΌӰx@7�ѨA��fU޾�;e�A��U�jGa�Vd��]���%��(�E3����8d���`Ʃy�~�Ѹkn��n ¢E�m����S �ψ��b�c(�T�#</Ϋ���]�g�X[\7�j�]�W7#�rjgx�i�`�J���o�Y-4~ܾ˗n� �܏�>�>�Qӱm����/y��� �7�Tԭ�Q�$�T��u ҆x3�©�g�^ܧ��f�ks���#O����GO�������g��t�c���H �Sիt�_����?�5N�� ۯ$�<�aJc(S�,1ql�a����wc���O��:B �0`fW���5Q��<�ǜ�0�%��۽�����s4��hv�Rt�.;\�W��@�RD�金��to��gد[�Y�2W������s�nz�D=e�-�͒�A����7��=��q;k�C�3y��,{��`k�"���m�.AeW޺=�z]5K!�c�y��Kʾ�O���u7���V�uGsT�Ϫ���Ur��--�����^��DޙPA�)�����5뺙h��e��8}x��8��ձ�t��<D�V���{����~:Q�R���d���3��y�������?vn�~���;�����H"&Y�@�a1^��Fy<���>�u����q�)�c%�K�b�Ҋk�__G�����2P#MR뇭�sɴn �A����k�. _0�b����U� �&#l:�/��VC�`�"3�c���xA�^a�ޒ_.Dv*� �-"�C�d Cxz���0�҃`�������|��ѻ�5��BL��U!�H{�=���/j�U�U�m��v��8`�BC�#�E���y�<T�{�qO�rWk�:*��_uW!u��}w)vu퇧z�r|�y�Fi7 ��^�PA��h���̅����m�ˠ��/���_��*�T;��D���m��^KtXT��kB�-4Z�mM�gaՇ,����Rb�53�����F�X۪H#Do]��~g �k�b۩��3��F�҅�Nލ���n����J�!C�T�N��N��/k���"P���1�N-��(���`��J�c��u�b'ߌ�p"FuY���?q�սo�x A�^��f���zB��V;hF�XYD� \�&�������:����^��D�"ez%z�g;��#@��a\� ̖*Z�Ĺ�7�/1�:j��!��À��v����Lcu�:�-�Բ%+�-�G*���P9�(�����4�pkSA��E�v�b��Ŕpa�+X^4�i,:�1�8�e�FR	G+��٣v�l6h�Ȗ<Ɣ��9:a`�@i��)׵l�pZ(9~��7MX�1l�F!QfK���t�̗�m�3�Mg����qM-�V���R�pDfrY�w��p���e��}��źytv��Z�1D�'ʐaC�x�͵��A��u��la�LF�U[ŝ�z�F���"#m��*�߳U�<Qǥ^P��,�"�ﶏl4�o�[�x^�`A�6T��L��$k�	�K-Rբ�x� c-"e��{��-���T}�PѬ�Ԋ6Q+���	�W���*�����5z���h��X��"����,1O�������~��g��y0骒��JKc2u]�\�C����>��K/(s1��`�\��`�n��w�	{��H����b �D ��?[�Iwǳ�kO�<O�j��/,�&d��чR��.÷��-�{��BM8W������|��X��4F���ˤ�8*>�@�1�2�*��؏>�A��0���L�:U!����y��l��PQ�LAP^"W�@�D0c��䦼�,�&%�!�
1�UC7�y�O�8�![S�	�X���� ҄�����\�!
�5,D$2Ke�Ͷ�m�����z�"Rl��|5�5�:K�r#�08QY����̎]��5��C1���'&����l�"E��gET2E� �Iz�p��!�Ctt�A��oj�� �*�&�d�Tt����!ab�WM�m�"��;i�f�r(��s�+2�SJf�a�����C�|��ؠ�tj[0��_�����f�Jn�w�wA�̬�jl�F!�Z�7Y�4|��`u%IZ�@�D��Qx��LD�����ƈn��yz�1�E���^7l/9�� �en�1�u�Uv��:x��P���ѣ7�D" ��B�B;Ix
G�ӫ�>�0T��/>M`��7�b�V���&�h���)�o��RD��W^f3p��>�ll&0���1����oI�'��1���5I��	���h���:4��ݯ4 �D_al)��-��h�D7���d�K��|�h�yN�4f�9Y��fSh)Ax$>R����2r�8#HDRRB�`j��ֳp��<>4P#��Q2g�������%/�(�un0N�qd3c�B��{��,��N�\�ʙ:�۹����7��@�	t!;`��, fSl���Z�s������xo Mj�B���x��?�ޓ�0B�l�_xMZ�µ�V�kA0��E�^�d<`��� ��^��vѣ7�'u״��~�kL"fB�:`h�6�Ҭ��|�2�Yz�ã����,1�,P����܃A�[vа�2/%�g�
@ �A�m�4:w�g��{�[V!P
�^)X��͂1t�U��P�E�Z�ϓ��cg���{C�pAD"$6���ZW�u�a�Qj��VD�S��d\8��\�67꒍�|D��~~;���k����ӭ���H���8 H��J�QABZ��� ����ܴ�
���I���m`�X)�k�DS1AT�,�i_#����2�
���z����WM�j�ζ�ZPXAHEK��B�T�db��(�x�4EPZ��"�ECH��I�s�>DDm���8\	Z�}�X,����"��yNsI�M����3���#�]yh\���޿����d�HfD�d�"d	$�IfD BS"	�	 �BRH�� �	�@�d��2&D� I�)Bd$a�$ ��a&fHI30��a A$�$�� �hH �A	0$"C!	�@�2H�H			$$���$ �0�ȚX$�c&Lɓ2#"D� HH$��������G�z�5�{�V�]�9Ԥ�%�t�%�;s��9%	,X߿���~c	1H�e,�E4͛�I���&fY2cc4H
ccI�K3E�cI��T�f�eI���RĚ�R��e�"Jd�h�Y)Jd��f3E*+2Jkh�)�6Y�S)��!4�Sf�l�22P�,��5FFF)1�H�����d���I�??��e���(���ח�>�/��	��E�AC�DO�=�%-�[����up~"�A�/�@D[�+�������t$G��
((j~�����w�Đ�q����a\w��_Xџ�l^ v� D]��[���ot��[*@�gi���v�5���X=yd��DC��ԙ,
((M�7�}�V얟��Uj"�>�*�� *�锂�p�� ���K�"�B�`�ZD*ŏf|��ey���Oh(���2a �s�PD_5�>(".�����t��.��B��ŝ�!����t=K����}����u�!��G?�
�
�
��>Htϩ�||ӧ�c%�>�t3֬�@�h!��W���ϣ�>�T0�!�T���rS�g�x�ϐhvJ"��D�"@��{�Є���:�K�4�}�|(b�"�X=`����>����c�E��Jv���AG+��650�+����YUPP�d:لH��6'ZX�P9ɢ�����b�����2���S _�n��J�q4��E���GА-�v4`���[�0(
�|T�Q���y�O ��w��
�����@�WϢ�������9���jC��[
�����z	����bu="w�x�|H�B| ~���Wi��/��ȥAC�y�q�u�E	=�Tҧ���@�'�AO����Hh�jI6��mQ��V�Z���Ul���mQ�Qkm�b��-mE�ض�EE���Qlk��l�VصEVض�Z�V��EmlZ5��V5����bլkQZ�-�Ej��m���V�֋m�UQmhը�U�EZ���Ub����V���Z�Vڊ��^����f��~�pD]�c�����Á�=U��oѺ���"��$,�=�w,�d-=4ys�c���׈3��������[���tD^�N@���C�  �&�>�8�b�|R""��*"���s)�n�D:>���=�*4��v�`�P| ����0C�X��`��^��E����uv��b�����ĉ����xxRa�
CR!�-�y��20�"��!�
��]�rE8P�|T�