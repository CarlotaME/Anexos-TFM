BZh91AY&SY&��7Ԯߔ`p���#ߠ����   bF^�@      ��5j��k&��[,гj��(��
�lT�f2�$P�@a
JTZ�T�l�$�QE"���)%6�M�6�
U)T��z}i;������L���V��Z��ij�j-�֦B���S+5L�j�4f,e4ɪ��cld�5a���mSR�k-�SJJ��l�� �( c/.�[-�Ih��{����V�fL۾7/F���ŵ��Ξ��E����u*쥳d�6��k,ԚX���V[[D2b����"km��Xc[4f�ji�SJ�x�s,�%j͙|  n�j�����ӻV��ve]�����[�tNխ��3kmC-IV�J���UW.Du]Wm2��N��s]f�f���v�f�Z��T�5+L�3m��  ��P� �'j�iZ5N776áM]F� m:��Gl��Gp�@y��[t:ʅ�W�N��C�n7�:B��r���� һ��3[F���.����Z�p  ��TQҚ7�k�QA�M�{���ӭ:�j�޺t�(oJ��h�8��� �{.��IS�=�U�*����w[y�= ([x���z= �kmf5�����i2lf�  vg��hSF�j\�^JZR¯.uJ� ;'��2P{�<��=��G��]�ݍ4���掽څ
�]����eM�K��Ut�:r�t;���w6�TE�ɩ_;��3cl�گ� k�z���{�@z t=�W���R�Z we�u��-��W�CM��P뺗N�J R�u�r ��V���8��f(�2k$kZ[4�  f��t�s��;��t����`*Ԍ4kRj�7[��v���Ӗv���k�� �i�SZU����tܭ,��+7��=2��i�x ׽ 4�q����n�MPt5�v.ڹ"��s�5�t:�;p4�c]ݧ] u���k@�� :7qph Y��5��ZKv
馩�j�  G�P�t,E
��ZG7)F�F��J��p 
ͬ��v���\�tq�E
���:uZ#vS5V�Փ3^�-�KZ�� wx  �Y� t��ݷ�h��v� 8�Js��4f��n���4]�
փ�;��[j�A�kVʙ��R�O  w� ��� S��Q@(�P$���
�����w7t@۪q](ѫ)��sq�
*��  )  T$�     �50T�Q 44  h *�b����ɠ  @ OɈJU( 4�     "�� ���40	�FF�h` �@5BcQOГ�zSdɨ�6I�l�4i
M@�RPC��  4`��[r��8�3b��b6L�����_E)�Mo�M�ϳ�n��g0������� (�9����PO�@AE~�������Ґ'���~/����q���@Eg��U_���ª��ʨ ������G� �(����(�
�)� �:@����"��i�@�����4�L!SHQ�@%SIT�t�L$!SHA�� i"�@������B���#��i(:J����i
�H����i :J��!����i :@���i
�J�+������ J��*i
�H�����i��D��*�B��)���"�J��)�"�	�i
�B����"�*�B�� i*���*i :@.�"B���i*���*i(:J��:@H��#���
�H�����B�$U�P%H�t�%SHA�t��IT� t�!HT�U4�] �E4�!4�%W� �:@	���B���b��H&������� � ������� .�"i.�#�PM$�U$@�t�M$ �$I 4� GI�Tt�] HA�p�I4�)�� �� ����*�"�H/	E�%GH�t��P�t�$@�UHT CSIQ���B#��@t�	!�U� GI�t�]!I�!�]$IT�4�]!SIA�Q @�@t�M!�(�J����"�J� � 1:@����(��@������\!�!�M � �M- �4�H4�It�H4�I�, �]$8@i!��G�L$�CIt�I4�H4�I4�!t��]!�M 4��t��M$�!�]$�!�] �H4�I4�I4�I'J$�!�M$�HL'IM%��I��@i1	���!�&�X@i*$S	Q� $SI���9�O���_��!t�k��|o��V�J*�?� Ƣ �g�zb�s*D�m~կp���W�P\��RYܒ�oO]!���qѬ��b��u�W�R�ۡ�Ei .��+��i�z	xm@^5[DS���H��-��I=lZpp��W&�6���\N�쬩L@U�GkChh��]�l�ģxF6L��0�-��qm)��
����w�����ssr�O#�*�=I^��)3�-�8� ��#A����Ƶ�T@Z{�����b��e�lL���e����	��sR�:����,ڻ�j�4h9���i�׹f�4�,�
�h�m٠���1H�u'K�o�i�;x��ф�轄�q�A7�E�j�Z6)�9#���tT6��c�v�4FdƵ�ܶ�e*�Ɲ�k�A��Z�n�G��r�NS��Z-fL�a)�W���iq����M�Z��j#��:tp�m���+a56��wf��3/f���`�yU��M���(G�5k�{N��-�Ma@e:�I��;��݈�R�&t��F�T�C�qZ0���-�g2�)���G �hMԳ/p���&�I�\7(+g�U�f!4mlUwV�m^.b��>����V"h��.�f���y�:��3UCEY	Z��TL�r]�c.嵖�be��VPi/fd��3�I�p@)V,����݅��B���J7l섳dl���2�7�*G�a�D�Hˎ`��Ȭ��r��	6���ǯ3lN��a�3E��D�ED�{���:f'N��0�u�O]]�ݎŅn�$q�ɚ�|���m�ɸ酴3#cq�j���H�܊��A�JXI����A֍MB�p�T�d��/aUf�ѸŠ?Y�`-"� �tҀ���*m����9z@�����f��tS2n��t^����@jLQ!��5NZ���� �aC��M�n��N^�ӂ+'�U̘�n���V�ю��N�O������l�C讜����ޚٌ�e˺g�Zuk��"Vn��dkZ�Y�vS��O�iX+�ϕ�����F�C��t��M���s�y"�or��E�LV����R��'�i��v+u�ӵA�eo蝧�J�r�2AF�0n[ժ�"��)����[�v�t0�(P.����l�M���W� �X �F��"`�t\�)E���[�h5eء+&E����� ���ݻ�S.&2�n�Lf��٪�n$�c7K*��7
m�XhB" �Z1e��2�lͱ�8��NJ�0������*\x�*�uċ<�+�ѧGwz�
��'m>���F�
�*�۱N�W1�l`��*�;7H�#��G
�V�ɰk��d5�������q��kL�� ��n��
X(QGF�S&��X˴⽣B�3�u��	{�F$ݿ��a���B���"��6IN`�X�pDh�iËQ��g@�b��,�x�m�s+�qV��Y`&#����A��,^XA۶�f��Z!ٶ��,�d�a*�EU��@���&=[�01��|Ν�afDt
45�[P��Z�Ů"�SvR'f��SoH+M9r�f�y4��SǊ�,s�,�H��.8J0�%�����d�7�㩅FD��-�rbI��{��Z���1Mi��Z9Mf[�h�o-\V�2��`;�$˖��,V;ǔ��N��fM`b�3����]�ej�U�]��L��p�.H�[��Q*���i\'n�P ���;�U�j��3/5�Z[�!qj7V��V�k\��eD���Q�CˬQ������Ω�aưf�7W��d��F��C�UX�o
��3_�X��Rډ��*5���"�b@Rv\��m�wUdÇ��л�wgU�6�[�u��Nu��A���NL�����Q��V45)cP�{�٧�M��ʏ��9Va��ɵ�6ʗy[K"�wu�eA����ĴF/: ��cl���\���搥���W��+���q�3Pdj�h��x#cD��n�b�'��JL�'��M[7N���(�P$(�X�`�اroz�Sz��#�Y��k
��e$VKh%�Su*��p<p���ɲ�`��N�F�b����RX��C��Y�_W+r�f9�CR-��[��cj۬��ЂT��f;U�Þ����n-xD̻�(�m:+ �R�M�2e޻�l��0*��ÇpmM�J}���Q˿����!��C8-}�wp�ַZM����ǟbaRDz�v��r�A���(�q"J
�ޫ&̈����a05;�/˶0�
�p�:T�"�fR&P�?�b�)��]��:��=�		Ǫ��]`'i��n�n��K�w0<�?H�1���^��jt3/-��oѢ�H�5��+
��m�/,d���e����V,ն��]Sj]�X�*!��L��An:?�e<#-�x�́��n:��9Zi!�A,�l�'ݡ +R�p���_��f�s8o5��=#��6�V,\�'u�Z� [�;ߖnm�E���CLe��'d�	�HZ���9u�q��ئ].����Fj��w����f8s��B9�
L&6�����0�Mֵ��c;A'Xh$w�Və�s�"�f8i���f�u�h:5���N&���S{I^+���kd]ót����`.�߉4ȷ/T;�JQ7��[[r��ȭ��{��RB��)��.!����3��bG[y�ݬ�,���of���u�ZJ�cd:�C�U�D=�E���q��U������Z1e0B�+2Z7��z
�[x��!g
z��Lm�LU�P�u���
Ò�Ȃ�0���p']]�4L�� .�
id�����˽VT��d����٤��K�f�f-SvY�[�u�cZ+$�S2�M��-9��n��b���K�6nRi��Y�,�ƙ�����; �FcKXizTلM�d3.�s/JVMQӘ1��OH�+%x!�3�2�좵���T���5C5!R�34G���:LDށV!˺��L
�J�2KPQ�RFGSn�]#0���	CqGQT�b0�(|�m=��yl픇E��L���c:��KQ}��Rl2N�2�/D�܈�0ܤ��f��[7
8M��z����l#Յ�%��6�:D\�dV�����n����?�}�6�{�v��L�X���2[�"�T �N�L����^E����ܙ�t��袜���(aו>"���fC���Z�ݑ[��=X��$xAO6������Ɣ�Όz+%����V�+Ӡ��{��7����l�MiH�4H��P����YJ��V��-S�\L�-q@��6��%3�Ϭ�Dp���*'��o�%AѵZ���J&�� ^��Hz����-�<��YM��q}�8�%��0V��G%K-�u�G0U�Ivte]�T��!�gY|�*�\V���Xq	�{t�&�h�����3b䠊��8Cү��ֆ�z&�$w6���bV�2 �Ȏgش�)5,���]��v%�\��l޽	Rͭ��$]`S~N�ת�k)�(k����A���#�FB" �#�ҳ�Զ�/hzSZ�V]J`�W����%�í�sV`�CGnl�{��q�ˤۧ�r%���z%L76�D��tݪ[P�������ji����IIh���5��WO{1�p��
m+r�V�]�d��ڼ� �����
�5dlǷ����z��feA���r����5YM�rU�@h^@��%�`�[D��[tvh�WV�kUbs$�L��wY��l�Z���9�f\�Yze�&��lj���5�ٌJ��`��m�֝�c�����1+F��]C��MP�zY1]��ӷp*�473C�R��c��AnXbke�jԶ�ͬ��RE@)�a{6��ss-APܢYs�d֔r�Ճ<�`�ݤ�r��m�z��DK(a\�4��w�͞(���s����h6-
���R�U1���^Y;���f������-�r)5�p��zN���ɚڗ2 N+4i�"h6!9t��J57 +73U�/�j�,`B�;m�5n,d��A��d	���
��� �7ԙu��d,[�%q�]e�1Tn��џ��+.�:�&��2�B�X#�T�֧zoF5FK��������P�mV#�a���(��*@+EBPԝ;z�藺�P�7�������k{����.�*�-��7���4iL��M�W�T�*��d�ȹY�,Qx!f��J[1�Shk��)�#H�Z�0ll��� ��T]�d���kU[w��ֳT.��ɬ�f sN��AbU�`.������v뱺��x���2�xN �u��2�(�ZP���]�hbw�6�KT��aŶ᥸���I{�(1Rl4mǴ췖d{��!���R�n�Y��5]6-�6RTMG(�y�Ln%��K�5˱��׃#�-�Q���0t���Vf�*p�*YDnm�q婍6�C-ldVj^H]�U&��%���L1z�U��P��������c�괓��(�aQ�m]�[%��QM�RKM�Ťn��3N])��l��L&m�g\N"�ܧ��\�J�4�&T�X�}h�Sr	��ӎ�b�7�<��d�ɠ�q䧥�H*�K���a��-M�vsS��iFmm���	�ʓ�"���ta����]F�$�!�ѽ+W�/m��yZV1֤��A��΋����0Vml۷��IsqV6���2ޫHm�B�P݂w�[a̤V���䉫�t$����1ff�<1���f`?N�{D��y[�<���N�nb��ƅ
��1��+,�R��B9�`�D�Hi�[P@/�Y#��[�N��Dn���e��7koM!�R
:�N��U���f�Ū�C5u�	�N+Եͦȕ &�%J;B�.Z4r9b-�"P�V�Zz^m�����B���$���=����:"�H�4Ĺ����0�Q�[Pޚ�U��M�N��@CRV�f4ʏf�`a9�Z*�\L�*�T����_��!B�݃^r���� ^�x	E�&���=V�[�J��ق�����]�9��  ��ehe5F�Li�ZN�X4^Dk@��1��Q�������C�9��6�J�e�fS"c�Ʒ�`�6��l��u��b�ѭ�F��Xӎ6��ƭ(\���K**j���$�xӫ�
'S�Y��l�

�쑌��t��D�n(�7��NCm��fJ�r��Kj�KW٬]L��7��
W@i-��T݄%��`wK�Eg5Z���D$�컶�{Db��ol�X� ��K+wԩY�ǛJ�v�Ń3BŹ)<����aAPS4��$�j���C[�#�"�ɴ��۲[��8��89|��;ekvt��]e���@CH�x���Y$kL����ڑd8���J�*j�P8L÷j��4��
4�d�4�9����K�sd�xҢl1���zʛ��6�k]�v��s��i�*nf#*�9��`�P
ά��47p*7Y��&��2,�{� k�V��[�i6c5&aGp��� ����E��f�y�f��P+6S<���6�*O�f(3o�WFTYr�GI����R����W�Lcwf�8��2°�-�j����i2+U��
i�wi�4h�x��j��GH�"��{q��-JL�SVȰ\j�QƮ�a{�����y��2�?�-S�
c*n�4&:(��q���,�"ә��¤w^G4�SRx��Q�E�FS����e,r^�o,�AR��Z�U�Ykp�l��Da8�7J�B�jZ�O~��KA�@�.����S����hvҾgBկ��;���ɔ��I�bX�b�w�(��	@m�[�C1)m�����ZA�c{��@EPQ�,��̢$��Rn-�r�I�[�6�]��ɵ���8�6kh+qY���G^)��'X�>M5{�[�V�����f��>n�[yz�#�LSG&á*���[�����c1E��Ǻ�������&�(MT���n��y�(DR���t�24M�/�i�l�4��C�TB�Z��<ʹ�2���j.�c�Z96�J�-=ȶ���2�-n�Ɂ�����5�[��jIi�^�+��E�sv��VkF��m��ЖӨ���Բ�*�e �8V`"�ܭ/s�[b�$u�R�u��k�)�[kV�Q�F�٤�8!4BJ]��������PnшA�J�.e�wXf肋�$!��fő.�Q����U`L����/rVm-�@+F�MT�=�A�Um�*D0�ٓ,,JRcI��wP��p�E@n�֋N��Bp���ĥ� ��46�����n������Fڠ�iO@�e\�C�a*ƀp��YZ�R�R�F�Y��Ȩ����vK��	pM7�UmԘ ��=�w�[��� ���)0U�cш]�db�N8�y(���'��d�p��e[�k%M��ȥKJ�41Gr8�$�a�ٵ�~;#�R�ثq+��+�^�r�M���� ������k��XoQ�
��T�i�cr]7MǊ��kbʐf��z�++&
!WN��j�kn��%]��o���(=�6��Ǐ$7t�:T�K�j��7i9��*�iQ�F�:�J4ãӁ���p�&���zz~8|vGG����p�����8x`ǧGG���vxi��Ɲ��������2T�b�4(h��$`��%·�����4��a���p�C��L> ��=:
�!�B��48�B�
���=4��������ن>0�4P,X��2T��F�0d�����4��8vA���Ў�Ύ����HÄG�g�a���aaRI.Ib�
(P��0h�C�{���F��N/�K^��^<z�x�LҔ�Kq�FKk�����L���*JZ˰�f���w�j�]����<)�/Z�׃$S�Q�͸K�r�7&���v�e�W)��ێ�l"ڸJ��4�Mk�t]�,�`�`R\���V��6���zJ��ٮp�6��X�:a��&S�,�˼ڨ���N��f��|�>0U����i�����ݹ�рT��"$nv^ȝ�{�f�n\�wCh�/�gr��
w�}�O�g�������}���k;n�Z�3v����4�wd������7�k#]�9ߜM�5Pf���nb�]���iN���z���h���ڌM����_^,�`�J�)M]')ۻ�,��2��=z�M��S��:_�4�8���p������C8>��|�-�띙�U�=m��6�o��¶L�,�Eh�¯�j9ݵ��n׮���JZ��'%�!f��M������LzUn-���ݺ2F�FG�멭���Tnk$�W-��}�si�3�,���+���ȇ7�L4��J�B��4�qtUZ�U9Z;v� kB�ݭ,����n�cYFZ�ڱ[����:C{oj;�<,����7\e�e��nޔ:'vr
dC���Q0t,�D�ԨK�5��1<E?�������v� ����.�ly��HI�:+3����;��x�t�E��f��}ܿ>�ǐF�f�ѣ��d�*������;]Ϣ�*Y�aa�s;�̵�����uY�!�v�)�n+��X�_�EL���r�^��P���Shk�DYM�h��Kc�V��-czj�`5���UZw9���I4��j���ʼ�u���s��pziROTo8�B�}QQr#[:�Vh��K���� �V���$hl�����'�+Pm��砨s���s�B������jX`��'u�[Gާ-B�uz�:hM=�k�vHJ��6[AKʊ��ȴR�|�>)���SC�K��D�0	�Z?�p�Q�r��nf=}$�֭�WLm�[/'T���@z��|�n�R�q+/L'��*b���U�q��gy�b�b�; ɭ-��0BwYv��ۊw���t�s�(Z�q�*Z�+^����������C[���^^�R
�m9��7:D�5�/C/����"�,bn6h��m�l��fQ����"���:WK+/�o�8��6,��gQrֽ��r�(1
�suN`u]D��w�+��9r�f�&!����]ժ�+���X�� qZ����@fv7��:}����+����򘱖`耷�)Vr���e�q5$J�W��:�<�Ɖ;`���w�d��2֭���]�����'i2[�.���d�L�+y�$�t;�X��]��сKrt�+!Q!���齑qW+�^frYR����=�k)���Պ�k#;���g��1�ɂ�������1�غ�ْ��v� ��CJjwUü���s3^�*]Uȇ.�+H��ۜu�̾�X��(��32����-p^��ueEv�0D�b*��(�⋅��39t3^�[W�!�R�5�xƑ:8����_P��q̽��J@�s �5๵:�.[��̾訊֢�f�t�Rߺp><�xm�~Dh9�[I[�[N�V�۳z\��gQ;G�Ęx��=�gK��ۚ���%m�D��Y�B���ׄ6��meaCf��\W�5b�VY�\��:�E�[�@�����veʶ;_�2�:�/l���4m�K�lol�$]F�&s5 �nJ$�+=e1�5]Y�|�gSÏm��u�x���x�5xK�	�kf�Ũu;S����n��Ӧ�R޴/4c�'0V�A�n��q �/�;�[6[kuԇXF�w�l�]���sBK+��;,���o����J}o��g�� n��s�6��݅d���9_*�Z�O��&γ�m�]Y�dl����\�f�Y]R=�'U�����&h���x��4�=Գ�I�sK- �ŢX�չ���c�oP
��c �
gfD��ʃ���'�;�Ṗy^�^:��L����ncSp0H��\���L�X�WM�ͬ(<|�C�n�WK�k��L���Nا.���!��B��k�0=�B���A]���V�Շ��*seγԠ�]m��:�̣]V1�Z�Kd���Q'�߀��T�
�M�K/���5�`{P������t�\j�J�/�7�̯y��׺��=����;V٥i��X��GwC����1�Q��Xٙ��N}���w�ɭa� �x.}J�hޘ{��:����	i�i�3�IfgMog�ҽ�r*ާFQHhdJ�3!Q)�⛗<�b�I"}$K��ٿg5c�䤙��8i�o(;��_m.}V�C����q�
��6��#vą�k�5�����Vތ)X�ةBV�oB��ꊖ�+���B���T�����e&���(p�8�K��D��ݒ1I�*��=�f����^Nr�=�����WG�˴���T�n7�jd�N\=�3��I���ͯeLd�yk����4��ފ;��-�X��(�ُ�*o�Q
ó�M��`�ժ@�RK���Ig:��₯��+�e�Bp�]N�2�,it�<��|����]į���V/o� "�dΫ�"�;�
��"���(��A4v��)n�9J}�Z's~�\	�M�9-�٩ݭ�"�`a��u؆�������JU�Bέ.(�X�sX�(m���P���X�{�0h`���Aڀs*,�շ!=w�$a.h��:�o�o�trt��N�_Kl7� �a��Y.��%oIز���6����p�� n����-Wm����lc6�j�fJ�O�֠�^u1��V��ݎ����2�b��F�u9�^Ү=ٖ�,���r�C�7y�q����u����J�lݛR�/��k�0�keP.pt�(��u���sN��fr�uͥ0�pA+��X�����/��$/.�w�i]�
�9�9��5.@�<ZhAJ��;�9�+W;�����j�W�*Y����k�ݕ�.е��s���㽂�E�1�a���^�z���yI��)Bp�e	A{��0�l�֘�x	�����> ���p�oMr���0n�aڭ���O}�?ҥ�*ri���k�ȣ$�����Z5]MxP�!�{Mk���ioY�e74v��Z���S�j"�4Q�­�.wO�����%��v�G]w��g%N(�V��E��4��_[���v�վ�;���]B���㶈������n.�_4�@^�}zk�jJcI��,=��0+ԳZ�}J�T�J
�Jlg3�M�%�:��p'Pa��5���n�%b�q!�tUuec
+�������8��s�p�g�t�
�:��;;%}��uo4��ڍۆT���d�t�̼�r��L7EW}�{iJ�v�*M����ݬO_'-mb[X�����)]Ѿ�N��)+��7��@�Ep�����z/s]���f\�����%걂�\<��)[]�	�v�Օ����ǽq�t�7"��	q��6�+���ny��n�֘f�ʹ�F��&���Y/J�Ε���2���ɥ-S9�͹���Pr$.�d&���@���@[RQ�M�Ўa�ߧ"���B�$�l̤��۝h���)�*�""�q�/�.$��;�FZ�(���^�̮/jid�A]`�ӑ^�˾�(��/��M�\�wR&_�
2�=Ty����REl��v��c[ [��{�����YA!L�pWg���iD�sA>�tB�`<u�Z��EU�P ����ӳ��� ;R��J�)mK��2#�R]N�4@;��T��7��w�"�l��:��a�36�%*̍�J����MC3VZ��A��ʰ�Få��^r�W8��mո�<|��[��|�n�EXP]��qn�_o(s'�NU�=V���V��\�Hg^��'�l�v�n�ٷ>���8��,D�"�J��b��c0��x|_WD����0�̝�x�Uծ.���eB&�v�VB%�Qmʓ1?���<rBഴ#Y]w�W�R%����|����M���[j�kT��𬟻fɓ+������W������+ ����a�4�b��Ei
��c7�E�]��{/ �
��W��k�d[%+dj��2�[��5��e�⠭����Y���t��ԼT�j��v뙽����)����9��p[h�[�c�+܅Ng6��ƌW��U�8R������JXޝ�� 1m 8j���7t�uu��lU;�P�A=��Ѡ�*��u��%��G]�{�2�=K�쀭�YY4�:FRx+i�u7ϋL��Ϫz?Y{Rż�'rR���b����~F���%�"��5���P޾��K3��VY��U�ʅ}��-�z�E�-�w���Q� �3մr����Zv�x�<�]9q��Uk��n��f���μL�#x��i���6v�&�E]�Z���S��J�Uv6cuq�jɛ���ۣ�XP6�J��npJt���7\z+�[}�"�V��T�2ͥKwL�&���ט�wn��m�f��Y�_�p����%D�9�j>��gj�/w"^^aǵ8�1���r��Q��&ub��s,j|�[�"��cT��֙�Y<��1�n�4�8^,����vD���쫫�B)+ڱk�y\4�|�tU]�^�vr�a��:���,
o+q���;�N'M�*W'{�P���Oo\6Ԉ�q1�yѝY��|�{VF)v]�B��3����Jn:�9�(闪Vʇ��Z5�9�`7Ʊ5};�j�Q�U,`6U<KQO�{4e+Y�l�R����|ݿ_�\Gܦ��/�97��Q�&hJx�����ւ��a<��_ײkZQ�X}s��;��ܢaZ1��~bZ/�:Ȳs�wV�b�qNJ�wc;%.��1�7����.�Ɇ��{:�D܂D�fa�`W}{9NNE�!M����M���^�e̗צ�4�Á�j�}�+bޕ�m��[���./x��R
r�k5����X��e=)�2�)ړ�ԫn����1��֗i�Чx�z�Α��<�ث6��bņ���{�N�sl����1�GWL �����#:T�}�ffm�jK����p��>xW6ر�ɺ��w����;.e�N�ZfZ�s��s����dlHѶl�`��|�R��H9QV[�GN�;Ƃ�~g����j=1@i�۝ȵ���X�Ue*�Q��*�]h!�z�fЬ�*�bCd��ioqq�;��f�r}C'�{W��t�Y�,8�����t&l]�B�d\��vlȰ����Gkn��$M)[Q}q�nE2��Y��i�lR�	R�X:&h͋�����-���Q-���2S�FNF�m1�(e�+�Sd�s����d��B�ky��"*�rv]�v��X�ٙr)�4�hq�y�C/]�׋�������A|К۩m$a����	�J_^�j��S[�2^Bi���B��ue�֌�
L
JN��Ή*��8ll|k���!�]z.gMu1%I������~�[��[���B�Sr��\��C���J��;����j]�+V�'w^��L#[�^Tb��ny�$Zs��9�;r��EֱQUw�⯸R+-R���`�����\5���Y��U*pWbl<7CܭFUf}��d:m�%A�wox3��v5.�t\���������}B��U�,-��%���]���EU�;���Ρʒb�&�B���Cf�h�M����r��R$�#�h1��Փ�1
���U��[�S*��2t¹E��icX�T�v��o��Q�n��9���mZ����t�M�`�μ1iʎ+ns��V�-�:�:W��A�R�F���L*�T��qޓ��f��.�K��u@�ժ�15śC_T�or\����L5M��|4�A}��\��y����q%�:��e�M<��[>2��l�r�WY�}F�u-�9]u:u�ނ�$��[/*T��w3]v3�	<t]k��:ʌ��Zۃ/UlBD�3h�����^�rࣖ�폖�hk��SoLlg��tk19�����}�}p{Ұ]G��-wֶ�d'3z�b�ik���hg&TTI�M���:Y@b9Y�37溻_��
�.��b�1\���qf_K�>����YPy�Y�����Ƣ@c�\�5�^�	�5�Od�G������g�^8뻎��ڑ��+�����&��%3�*���K2�������8�v:�t���] ��U^|�v�,�:�xH�.�:�*���Ћ�}F��k����:h���3z0�f�r�a'w-���=�;��wt�D�V%"�tΕ�[�����Nc�O����u�;E1Wz���p�%�Y7G�g�l��[�,[^s�}eYn�`��F28�/��ƹΰ�>m9�gM%E�7���:͡��U�qႋ��s-�,�8�K��)O� �]K)n�&K9AY[e"2`�1iWp�HQ��G�>��Iʭn��9���Y�Ps&^��^�`g/��P��Ȧv�����<��ʒ���o��f�r�C��\wnDl���B֭���BS��(Q��t`�V^�q�9Z�/x�5�ٝʉFt��$�GlQ�!�����GO����N��V��xm�Z�V{F��Tkj�49N��#�ؒ�]�$�E�t��1@dI1����Sf��3�n��'"}H���@������C�%EljH�/z9�f�T�)%L�˄V�/�W�5��왤�$�I$�I$�I$�A�c�M!��뫗G[�o�(����X.�F�0)&?�R�eIJsP~�(;��f�U~8aB~$4��]s�L�(����n����L8��+"Xa�RR�\�R饗�}]��մ���l�\��:����/���V�tn�rƚV\m.d*%ԃ56�q�j-jT��vڂ���ۣ}7]�9�����E����uF�r������m<�(ַyw�J�Ἣ*t��܃���۴rY����+���5V*9[��E���'��#A��iИsV<����AP:� ����Jh��-jT7�P�9�k�B��[�+�9��{:�jΌtZhث��q�l��vva�B�$�r���R�I�8(}ZP^ث�]w̴�v���LI�Zs)��3�;<Wj	����Z�����^"�V�Ði�<;{��N��wJ�^�W1��K�dܘ�Kr��J#	���{�є�,�j����^Tk�S�k��.�.*���d�ܫ�]w���*t�el�_2��lH5�;@�V(@w���I���\j��Y� �e��ה�W��Z��6�%�e�=w�oWSeտ��o>檂�CZ��mfӶP��MM����ۖ���U��'�,�q�4�c-��n��v��6�*��צ�S�R�����N�X�:7-�p�RGԐ���K����G�����yj���~\/T�G������u(�2����V�)l嬱ٮ� c�n�B��Fw�n΍H;���Z����#�P)p���&�.��5�&ԍfv���M�i��3��b#o[�w��0��	m�m�	����J��E��n�K�XQ�g�+�t���rp�r�.�����Х3Q��[R�ɣ&�2I$I$�I$�$�	$�I$�MI$�I&	$���I%I8p�Å��8p��8p�ÇT�����]]B�K��p����`N�n�L�J��R�����YZw�9���w{PN�ْL��Ӧ�ío^�5��ɩ�|u�T�P���dV�su*\�&��g#ٽ�M��zɀ��{3)�%��/�V�jfiѯz���~�������tV1(@���
͔��䥩Oi;��rs�u���r�19���!
�.����ۗ��R����g0*�c\����^�x��P�\wi^P'�u��L�ω��4��Uk�2����jV�q(��6-��[@1�M�ڭ��)m�ToB�t�p�d����Q��θL������ۊ�u�Unf�����E]ܻ��)b�!e4G7��s�뽑�vf�"�SMs�Ҭ�����Xe�ݛ�ձ{w4$6�:�Wt�TU�����0V����ou૨c˝��C�^ޑ|��s���i:uvn���D����7	�`�-�@w[�&��g~�+Y��p+J8��>-��
{��WQ��Ok4L�IՍj��3�)ua@9�����C���vi��kkj�[I7%��z��gN�e3�F%a���n����*�v�6�{��)��	+����9*�Y����B�_�6`���1�(1U�z�,�oP4�V�n�e�U�.��b�����d].��*�Ʈ�P�x�
�l�I3�+G��-`!'؆vI��sX=�M�yp�����a��,h��G
8p�����������������������������������>>>>>:>>#����������>>>>>>>;>>>8||D���⾔5Cu�[���L�*��7t:V��l�.N�����Ԩ�+��I M���"ʎ-
�	�U3@�T��I�RԪ\]B�\,�m�J���R��QmP�ŷ"E�!�9d��B-�%S�K[�.�8Mu��#ml��o5�Yڟ�g�t�UvwH3^"]bHl�p��+n%ˀ��U��dF����_j�����x����H��|��唸�o���p���n3AvJ:L�1���[2����M�$�:��άl��g�͒�Su��i��R�^Y��R�Wb��:T�A��x(��+͎,��n)���k�]���5׮��'�q�a��K����np�ǐ�7�����c9�,DYV�S�-RNY�ߝ^lԔ�zct)V�k���誢��7u�ҷ+����0�wˢ��T	�!RD޹q��++a����/��4��S9K'�\�L���S�*1Z��3NfJO,ّm�@Mط��;U�l�j��S��kWLR$y����]��G��p�׮H�vC�VS���^k�2�+�J�Y�:��@��,k��Ʈs�xkj���-`��6O(]v��pA�Tl�|�㽉�ۏeƕˬ1Lk�S�/�b*-UxB%�XN%s`���WJyN�A��SsS �gE[�\r���ŷ�`�cF�4p�Ç8P�Ç	8p��G8p�Ç8p�Ç$$�I$��I%�$���I$�JU*�J�*T�R�:�*T�WZ&�!eX�b�}@���t"Eu�0,;
`9��m��-�4�
V6SZ��(��v�^ֽ�]x�1 ���k��E��Q�6���\����c����z�e�v�����-�v��U�^.�l�K�T���o��Q��al���]���K{M���[�xE�j<8v�v�-"�>����V�R�Λ��'�^V�rȣ�/�w���6���ǡ
.��Â[�l��7������oT�p�l��E�9<kk�Y,��w��R�5dw>�1���a�u�"R��%'�S��c%d��(�Yr�Z�<���r�--Ȫ� 4�t�\�����4�h��܄�Ԛ �ā���{!٥�]YU��V��ϒ֍�2��``��eqST��t��#�=�S�e�D�#]Y�gX}{����v����M������FAy`�ʀ�q�T$L�[RjC{sr��+$��2��^��ͻEB�ˇY9@ftI-c�7s��[���
N�v�TÀd��)��3{�9D������۾��T|�����4"�m t��t��,�dp.�iL]�z/��eNy�V�Į��Q�`��ɚj�L�m�v��xYp���f�Cuk�ǫ/Pkv���]i-���j-��G;Z���λ����ay�ؔ�e�������������g�	0`#F�aÇ8p��G8p�Ç8pqÇ$p�Ç
8pqÇ8h��8p�Ç(p�(ԩR�J�)T��R�6_.E��@-����2��}g5�A#q��i��F̇(�kT�U��}*ͮ��k��GP�K���X�ݬ�Y/Ip�X�:9:�m�)����rq9���S���:�g��[4�:�YGF.���̵u8��WT�"\� 8�e]:�5�ٙ�O�g_kr�!*�� [x�U� Y�9���-h��l �>�c��C���(0lw��F�R�c�H�1N;78=X��u��v�2����@��E�[[�$U-Ӂ�t+gX9�`Z�����
�Q}[V�����Q������=�ܥ:�꽂(��pTSS�Yc���;��o�:�rtyB�[�(8dw����P5tx���Ro��[Չ�T�ˌ�!��ߋ[F4K��P��[2���ү���̘�3��R�wwu+)em�ۗ�uE��<n�nb�'k惇Fm��+Y;��Ի��T�����ԙu���u��������̞ف�^��r!D�):��k(�`��NB�o3��-�>]�R�h\d=3-ř"Z�u5��&�Z^U�&��E�®�ɪBj܆�AК�L�jr���g_Z
�`U��왝���\���V1P\�um٣5",�ߞ蜾+zL<���9�ߦ]�ݲ�m�L�"�m�݅V�s��Ր�1�'M4;w3�c��|>��1���YA�E�f����@J��{h7����#E=+E�f�ٺH5��]q]ز&�+AN�;���т̤�ב���ԙR�5'mA���U��q�&Ժ�k�����n��1_ҏ[�L߁�8S	3�W)�T��1��/vwL岋�̣�%�g�l��B4�SO������,\�� �Fݯ�!���e�kd�v�[�V�yau$���9����%�

&�7�h����6,5�(��0�J�8kTs*¾���%��r����l�S|�ZU�:MuG.Ь��R>C/kΟ�}�@.(�q�+1}6���qBy
�u����rܫlWe���f㱃��"v�T���c��"ӭ� A��	��6�6W"3���� #9�� a;8�.�ZV��ӻ.�B�%LW���
a�a��\��������^wT���B䭻��=\h"�ģ����ϸ�N�r�e�Q�W,��p�Z;}z�E�T���I�F��Y���kD[z+3�*b�ͩ[yt�F��4/�1بɪ�r!���iP�;�df�j%*aSS��=�w�P�XaKjM3;��:G�մ�cy)�9�d�k[<?M�9�K���V����tuz���E5�-�� �{�u��t�r�եx�˺+[��PU��sO����^������u;1Z�L��	�9R��.�w�w��Pa�8ha�����q*.���+-�W����ޮp��aN�iq꺎e.�o�mr ���,�ڕ�on�Iؗ��1���+�7����Xq�Ϲ���f�$+����C�P�LI'{���:V��f�)�Ht�w�:B�V(H;o3�4�ֵ�����S�1�0K#*lôɺ/7���h$*��=�����J�J!\�D:�Q܋�%�|4r\\�[6h�b��٨�����n\�:fƥ��yi4C��ñ6��6Z�͗�C�R�́XS�o)ؽ8i�'�1�N����{R�����\���.²�&�t�mؙ89s/%4��"�M,��ڢ�+0=�J5��1أ��RY[��[�����/OqI�+�P�XT�ERS]�n�,�VO��}N:�#'Vq4���ۢ��f�_u��Uj(h��
RnL+Zn�9Nccw��g7�1��x��x���]v�շk�R��
V�럝p�CfS50vs���Ю�1�݅+�5-;;����-�tn�����f�s$����,�a�B�m�Z�pS�]�",^���&l�fg�ج�V3q&��X׆�k�V�=�Q��lR���{�x�eVҤ�G�gV֛�7(�$eݍ��vqw���mV�WSk�[*���*����� ����ܴ���R��kkp�,��h����eZih��"���ѾT��N/�qթ�v�x���Y<1-ݲ@�����ݔ�˧�h�X��	Y�����+��͎.QTxC:#�9�sq�ŵW��������ʭ��w���uʙ�!r1����b-*�r�=�h�z�	���iB����-V�y��B�v�]�s(=��N��`�B�jV��ͧ1{�\w�6�#�ΙZ6Wijq���N�[m!WdQ��x7��)S��ٮJ���	V�r�6�F
�qI�.C�n>�F�|� ��3�W�}�Dz����pS��Od�b�/hس�*Et&0 �˂Cz�B���	;G���:J� 9�� V�`�6���XY��t���f��[����ER�a� R*�pݥC���I׶��Ӿ��.^����j��Q��Y�:1��X�taγ)q<չ*��V�m�~s�r�Ij9�%����O+2m�3������2}��W;r|�(^V${(���r��n*ǳ9p�)��n��:Z
Iu�g2��[F�mtsmΏ;�̼�<V�2�+
?Kڅu�n�r�ҽ��2J9Vc��GV��Q�e�X݂�TV�����6u�����w�68_F4ڟ<p�ZW��k@fdd뚲�B�@܁Z�}�⾌�78V�-�֡[q���c����Z�&�9̽��k:m�\{r�S!��E	Ҷ�ҥް�F�c`��m �@[��@�/�_�刳2�lPC�A�ʡ�y1V�w���s�e`��XLgh]"?#IT�Z�P$E_F�H��Jv(͹W@F@u7l�Y�F�*z�/$R_\�ϒz;���{|�+�5Pr#{��[	=V�����Z��Jǃ5l������#�;��?��:��	O��G5�s�0�����^�WM�Sf�M�MX�@��}Ɋ�+X8�Һ�5�ݠ\|�1+]2P��V�T�vkU�u6��,d�u)��i��T5ū��d���B�2�n�K˔�	��)@5�o[��������vт�N�,OG���J�=e�6;�l9�L�'7a��\���X^�f�����&������~Ò�W�k��y�q#$� ��눮�C��7�޼��{�Ç*�xd������y���͆A����E
��(��� ��zsi����C��e��M��PJ�
�nL�+��k��@�-n��.����{cH��t�M��Rou�Z�ݨ�vM;Jׂ�F�U���-1X9æƧj����qg�hR�e�vyӉ��_A�?����h���]xHP����m-*ε�!���v�$�&�Ƶ�eM�G�#B�g$6�Q&�6�ݣp�R��Jζ��e��فus�|�E���n�8= t��t�K�Z��NtV��u{��sQ
���I��n�5'�����+]ǚ���(�&ΥR�4Y|�I�ȍ�س�>s:�iy��y���a��lu�J�<�f;��[�+��
�R"��F�b��	r�Cvd.�J�w�ׁ�����zv��`'��ůs�z6�/8MY�.q���8թ�2T�ʩ�71R���7�RTN
뽬 \�lwYWǑr�as[tq֑2q:j2��H�'	��8�K�VBK�c��S���V�ڸ ��h�ɘ�sY�>
��G �C:yQі��_�\i_��x����f�R{,Yy9��u����*���>ԩU�_I7 |R�Ce]!�V�{�sg.��w�WT���
����FRr�u��L�1���(��P�l,'�,��O�r'ٌES-��)>��p�yEY]�Ϯ��nL���:���Ax:%�]�19��"�o37;b�����VO̭Z�j�h5:�<�?��t�!�#vj�E|鲈�w��<ֶ��*EV�+��`�R�Jf���S�6K�yR�RR6�]�k z��ǰ�U��\�I�� �j�5��Մa�`�{EIe���9���CR�d���}s9=�l�*1X�n����QpZ�r��8D{Ŏ%���"�E�@>��G+���N(���P4�Ј�kj���:���PR��2��%ޔݖ�l#���J����;[��p��
���bm`�mh�9g�oYƲjkY��Z�V���}�� ���:w��ʛ!�>��аs(v:ʜ��B �@�T,�B���,T�P�
�5(ѣB�T�puD4G���,Z1����{t���\�#����I�}����6.F]�5v�u(�A1N�.�BW>b�C�3E-4���+��WV�;��Ôs.�C�ľ���L)�L'?t,p��[������k=�B�#΂��}ݪP�@��]_�����l�(vLM���D�YQ���yYp�g����td|5��o#�"u��ݦ��c6���y���tvIԙ����'��r��e+��ĎbH�r��Z�M��Z	���S\AD���e ���r�E\x^����ܟ��4��_st��p���ݼ;t�[�)�o����w6=u��Dg�Jz�hZKd�U�1rb$����T�sk��G ^.�*웾u@��l�����)�CX+��u^L9պ
����J��TE%ΕЎ�}�5��\P:Aq��e4�¤���&�-�.(P�SU�MN��,#2���R��NEvat�=�^�h�(u[���5#��F��-dW�,�]'V�c��,j됩��KB�*M���5�ifn�Y|�J�wR�}�U޾���2��}:��R��X	Pb�"9T���h\�v�`�B��'��y�mf��fU���9��®�N��K��q��f8��7#�wvރ�0�cA�;xOa͸�G$�佸�Vs)Hx�M����/�hVV��߂�������*���Z)h�$�29c.Vcy��1ó������F�=���xa�;95����
z����������xzxz{�T4y�1Uf]�Qf!{��4SE3 ���tzzzy�RUUQ$H{U�4UQEQUUV�UGOOOOOf�������̊�����0(99s0�*�y�SDfE'>Û�E%SIe�DV��&@dQEU�dQT{aEDDDP�Q��Uue��D9�'y�0UTݲ�N�VY	Tyo��h��((�(�"**�1��&"����#$""�y1A�c���0�D��9%PTs0�"��*����`�"�(!���9>f�c��&�� ��AB�*�[R��
�ud����_ �n�]�g���<g��~6�R�����ۼG0p]�X�ǫ�a`��g���Ҩ�a��F�����a�p]H�JZ�.�E����؜�ܮ�����y�.ɻ72v�T���7�9zAy9�MEᦋx���T;[�u1A��=�O�=�*x�~�sVA���62�8�VܶlS�+�'OsQ=�O���,�7����W�1x:5���8��q��M>af�.�׳��r��{�"�l1S��͋5��>��Y8J+ю@گQ�^J>R��ՒZK���}ڹ�y=\7?��_�3)=��vK�p�|�l�^��5~�����=�j{����"��]�{��_\�������8��|"�Z�t>��~��:�v���;���nv������/z�&�q���>�0��	����'O��'�߸y�9�v��wY�2SrS>����t�w����:��~�}��o�/7��M������lM��F���յz�GL�?!��]�������5�Aw�w�3p9 ��*׸��������.�q�]u�
�F7rN�A��]!���I����������ڝq�W�Sj���\ؖ*Q&�bY2:�Z`����J������^p{$ɛ~� ��?�K��pR�4�og���o��C
�sg���������=�n�UW�z��߳����S�K3�קJ��������ÿaG^��O����3�g���ˇ��F��&��{�ߧs�����B�����'�����S�	�U׽�]h�H�75������]ܙ9��j{����H,�N<�'{��zE���x�bZ�H��]{�Oʆ�F{_���כ5z���{ې�5SޕR�/�O	j������������6ܺ��unA�Agj��'*�ž$������ٍ�yK��z龠)A�_S�3��BWe�7 �v�	��bl��~�k�x/k�S�E�H�W��W���3�g�3ư���K��Qy���]%�Wꩥ�ۺ���5�o�kd
7>���/a�I��W�*�w���b[��W�Q/�v���J�%���JV�osU�-�,:ݲ����9:��,l���暄�:��g�~�}��S�x�k�רm?�Aǅ��|3(�V��Gm�����!��S�9�F�g����K�A��9B�@uxd74�s���A쬬�=͏U��>�����s�4^z��:E�كN_*�:����N��f�yK��>��2�S���lr��.z{�N��37�u:�+���=��A�z�W�ؘ�*��Ӑ��}��W�T���s����&����yr�ô�쌽;��}��v�_�Ў���v�[�zH�7@?/�]u��k�6�p��o7���r8��C����!S�9�g7�R ���~�U+�]�^��z���T���H35��?g���٬�ˉW�2"�����K�t�I�U7ڨI��Q:@�ꓯ��L�v�ʖ��3b��f��<9=�6n�F��v٦�	�]?������ڿ{j�C/oT�:Z��;��p�/������/�.�f�R����o���}���q_���m�^����@&��vS�c�j�"��;����;�����r��^ǩ��u���q��n�[�|�T���4�ɘ���������,at��^��6<�x�!?����Ń� ��U������N��z�3��w�㄰:�X�^�BqY�c4����jlg�}BX���%����/������n���.Ff���^�6�:^��3T_8�k�/}�h�=Cn-�޵�i����x�	/$�''kNLٷx,vC]�n�u����W�ހ���LK`�����|���7Ct��Y�����9s"ͼU���M�D�=�//�����~M�[��M��ݟk�9~$�Y�5U~ݰp�rՍ~m6_t����0���5�����>a��M���s½g���Ș���v>z�өm���-a�<���v�.�)�Y��/0O(k�7v=~�����{�}�V\t�gڪ�����N�r_>񩖉i�]�j����tMu�Oq��^�{u��.��=���\^�Oh��sSx��y��"�tݎ'q����u��zy��Nʩ����L~���f�����g� ��Q��}��o[�5�h]�o���m{�G���Wu�^���(�:r�{������$�8�w�:�k+(SSu�3I�f��bݬ��3!�`�sf�͙*�:�-֬}J��Jj����l�щ)���B�(#;�������Vj�Q�aN�[�ںO�5e��C\�O;6��;�'Pѹ4�	�՚�_�p{�`ʳ�Ƕ�m6�'}p�h��ݰel���#N����u�GD_�[9��ӷ�^�x#^�(���)`�ݮ�Uu�6����NpU�FXP��[;��>�-�V����(�~>]����q>|o~�@�jg0��&e�k���� �m��.N���O�iO��^��Վ��Z���.��Ԛ�t���1d���yQVNH�FN� �c��/�ޏ}P�Y]t��;ݝH��תլU7�9�^)�ث���nb�d�M����N^g�k�9�h�|T��<�\��,�����}>�Y����z�>�|�������z�@�.(�|���+����o=�}����j�~�D*�O�|G=��:;�x������wV�e�M��>�ձ�i��_ ��=�:;�滈l�5��D��x��s\�E�L3��xn���?w�O��`���l��gW)<g~[
�+o�z�,��0nq���7(�U�{�r����A���M�8׈4��Pp��8��sn!�-H�8�%kV��M�f�;݇gvqJ n\�>��7������`�"�1d��2u�9�U4��������ݺ�f��x���㻒8�ڂ�,<T"�5�}3�Ms�zÜ���i,��^�}%��s���w�y�Cgeq�Q�:�.?/O_O�-u������kfc#Շ����G��/�b����:C�e�ۓ�Ӷ*"�{�s�T5��#�B#L����;��q�{���{ѐ朓2����L��<Y�쪟������t�gg����f게��^_���S��%�r�}ׯr#�z�����b@|���,�A�$A��Sv%��/A�f��Ӥ{��mQ��B�q�/�dʇ(�9� ����ǰp]�)���'���^�["�}t��A�1H6����/��j�%���;����Fn�<�����m�o�׻<�@�zG_��vo#]��,�^�>�Ӧ�w��uw�u���Hj� ���\{��ެ��1p}�'���D�q�#�F�%r�̭��s[g-�kL�7b�܌3;VtW��~���9��ީ0-}��惝[X*�.U$�yU}}}���i�8�kO7 q
�1������|��]'-����4ܲ��9'u����������?�el��3w6����U����^�����_�֪���*S%�c��sy���v:�}��ˎ��H�=	�^۠��9�u���o���I0⍁�o;A����t7g�a��<�W�#��90y�>�A��t�cσ�j�t5��m;���<{	�׎9`�o�lѼ���ݷ�&�n� ��o��~�A��.���}G[I��a��׎N]^�{�sU��Q����ٵ��b��<��e�L�=O���i��/C���=ʆ�.\�cv��흫���tBWB(Cu]W~sj�2_�����2�Ϸuº _]f����oEM�;�!��j��W ����8J�U��F31$�֞т�n����|I�x�j�p�Ʀ�&6�R�������������٣�,����a��Le�法Ǐ�����ӛFs�'��1z�n@z�2�:X�^4��9{�u��,;>W�,��U2�/{���~�Ì�^r�=婘}�]��T��M(y�e����RR�y������舷=FJG,��Ou"��e6���).��giv��e�v�V��+�L��&v�ٔqr�E�Q%u�R/wtz/j3j�HNH�NE5���t˨�~��<�$�����엒���	7�Q�훂e�^M�^�֚��_]wyT���/vuk8-���R|��
l��k��H����T(���b'rÕ뿽Ž󕦜��7�{�K�^򙋒{[8lNm?W�J��E�3�[Y�yO���ډS}�T�B�]���9�zmwyMc�/���������Bt��*�<\咔�qx����n,���{��^��^}FNQx4�ώ[<l��i,=��#���E��-o�o��_n�|7�>���'hY��f�(�Xi����O�bF;4r��Dq��j�����J��)���f��������Ö��t^QÕ�����˘.�����������g�iZ��ɻ�jr��	�g����d�\��T{v��uK��g���vW����Z�����ww٦�����)R�Y�Z" l{o9�[�R��d��4`o���!x�3��ٜ���g�ʢx��q�P�T�YC�)D)��p�'m���ÇG�)$�Ss`����/��t�j�eu��'+�����V+�0Gk:S��.�*���=�9r����7��ݞk�j{�'�ad_5Y���oy�{�6���d��b]����cw�Y[7�{�?uB����N��G�gw���==�!�/�(����Or����L̯s}��O!�w��>%_N�r�=��o��5^
���R/ط�z����{.�����;Q��70�s��7�q�ߩ~��#�z���Z�s�*�����r��域�od�ȵ�"u�9��L�g�JY�BWN���Z'��i����^�4.�1�}Ѩ�o	��b;�@���]��d�w5�"o��M?i�t:(�����n����^�g�P�:+��A�N��C2=���al���ۯ]Y�fC����g��4[�ӕ���ףCg�Z�+�+*|�&`�LNz=��f�:�GEY;'�l픪�KQ��PgX��o)��V���N[o�C�+��YH]��`��;1��&W7lV�U{7��t*tʞ.�f���O�W[F�J���N��w��}aR��u;�m��tZ�i�,[EI��B��F�X�u�N�(�����s�xdJ���:��=���
fM���F�Qyz�f6��VO�{��鈙j�w�_>�I�A�0K駙�w��'�?E��,�%�����o+��(wXUN�x5^�o��D�Q�6�_�	�w�U�a[���ww�V���Wz��'�J�����5�^��3dC��~k�{}27��k�tO\޼��`��u9�q��g�z��©�X�x9έ[}��^�{ٱo�
�D�<̀�m=L���n��K/i,��]k�5�K�~����5�~w�X��׽�|��������i7�1�s�Bc"��Pk�^��.��w�J��t�m��I2���fRCD��B/���0j9�`��WE'����#k;�"�$o���."����O�DS���A�KӮ�E�j���ny&3��z�RNw�-�֏Ng��L�sJM�9��1��&'Bs�`QHs~kxH�����-HN��&:������WI��d���ɩ�U��G2�e�����b�]���������/+��ąR\����M˃����9�ur�Y�Q�4*��Hf��_��qZ�;��׽���1��h�ݘQ�|LrnR�e�zL���p&�4�nR%��bbܶ�;x�p��y"p=�����M�k@=u�+�9���o�.${N�	w�E�oNśԡ�8u+U%ܕ\��\4���	���n�ԥ���M3��NX�Y�98�[9�`֬f�=*�mZ氊Yk�!I)�wb���t�kNTr�f0�aڀh��]2Uӹ������x�y@7�m�o)�l��l���5b����oM�Y��œ���;�i������VŲ��n��ַ2]�(����%��W����(�4���7S�KjĪ#K`�͡j�Z�XW�h���2:��K���.���s���3���`m��n�j�V�n��w���*�V�=�;bx�0���v,-Sv���L;'X![�t�	��Y��u�sm�!<�L��İ¤�Yc]l�)�u�)�����i��.���<B�T��t��E܇-��;Pתw.�w�]�*��O>����2�|�[Y`#�\�R2�$F��JT��I�m�����	���h�w4G�<ɶ�uw�bћ�4�
|�`:v��-��Ve	��pc� ��M��®�e*ں�Uנ��Tg����R�s��WGճ,j�lO6�Y�oZ�U7K�ρLc����SAkz`7H�j*sC��k�`<��p;�Z�m�E�ݭ
4j4:�+vkO7�c �ٝ�۩�F�)f�2ƛH���י�UY�:[��)���u3%Y�u"�E�l.,*�ἀ��ךf��Eg���
�[��{�fC7����D��J+��I��������]�=9x���G$�jZ�Wq�6p�m�r�˂�p폗e�q�iDeS�M�CF$���&5��{�+6Jy�
u�y�`�Ko����7\�)&��ո�eQ�жG�ucI2������G%����u��y�)_c�xv!�*��6�愩�^d=kr�hW�f�MH�D7"}gy��nQ]���`y����r��j�ܙmd��&��b873Y"&h�K�=�Ғ.�.Ҙp��wt.�<��}h'�M��uD���9�ݾ�E�]�U�k%ә8L�X�:]mւ��+�۵�=y(��;�1��tht�T�WY����%m�M�P2�%��O5�ŋAz1p�� ]c�X�s��}J]\c����K�X���^�aNђ�%�&�[�*�)�7+��)ɞ�yÒt���j^�0�]m������9�������vAJp����2�+�5�Z�"c.�S�C)7x���3��.9���7%�ή������ ��-�e3-ASTU1SQ��1�0Ç���|=�j�/,�("/s��s���9����A�Cu.S0TD�Ϗ��O�ؽ��r��
�&�h����,�i�3)*jf�d���8i�����߄EydIAspxE����)*�
(������Po2�k/��N~?�O�����'*&�*�` �"`�fQDs�, ��s30p�g�3Y��Y�VFD�Ufu�")���#�e4�3	��#3*���j�0�*�,���,�
�eTS��*��	��)��b����M�br�"
��**�H��*�����0LSW'��r=�EQI�� �(��r"r\
���+�ĉ"
o3$����0��
�� ��*�&%�9e�W��U�`�Ī��?
��/�P~��gg��96��T�w�_=;t �h����R�$����|��ڊ��pr��|��N�k������ ��4�{�ՎY���H��L�n&q=�u����xO%(!OR#:yM�5lz�ѝ���η��;+���Ȗ����)�K�_Ec�gݻA۸�i/ ��-?y�:�-��)��s����SQ���M�Y����Q�Q(y�CMQ�����HZ�7�>��ɘk��N�EJ���Y�4��3.�\�z&u��%t�;�{w�Oy�KT\�/�l:�%5��Y<GUbc���p�ٜXL�uf���<3��E?j���&�r��.��ug.�5]���WwJ�a����fL�}�}�N��2j���d݋&[h%�Z�~x������.ǭ��'�����O�or���R@�Ɣ;[�#$s�����S�~8�Smx��p.ʜ�֡�ʫ�au�	<�i�'�䓺��}w�^��v��hA�Z�a!�I.9�������5P������\�{�S@l�W�n�����(�<��h�O�.9���9��ojWX"���(��R��oe�O� ���=o���:��
��!��]t�Q�������U���6L#?5>�h�q�]!�#Y�S4������p�ͼ|����f����X��e[��ǜ�tЦ��yՐ�ʻ�I�Ϭ��FfR\��w������_GkDL�}W=g-�մ��P"��nSV�Tǜ��amT�o�t�u2W:z+ym�,�)$���Y%n���yݱ]񜓻5:F0����12G7���L��r��U��@�����)�U�c/�޺����B؏��4�,�<`��ŦڹмƸԯ{�n~*��z�&J�`����1���y�-;��qk2g���ꛛ���#����vI��V�4+6}sS��6���?������t����r��|��*Y��:��\^��z�~P5�C�4S��	��jU^�֪�޸�	�(pU�=~b����/��U0��%����Ϳ�,�������1��\g�e3e����>#BML��F�t��	3�U��ԃ��x��~��|>� #���1��\�K��sp���]��j�ߪ��%PV�Ng��/�j�⽕%N���>�)Оv�#��.�2A���[����Z����;�])�����i�J��r��TG�TH��yfEМ������JZ} �K���}[�~��,j�q���_��He/a:����1�S����P�N�e|�z�/ح
��);�%{��`Z�@o;�6�J׼tk�b��W"syV����/���1�w��Ч��pe�=8��9��53���N���r��ˁA݁��I��7ƯzG���ٚ����^6e�wT�7n��J�B�P�N��W�3�$�Y��L�2�Β���/R�'��1�:b�X�ůD�XF�A�S(�5�r�^��L �/P@P�U]*59��j�ٳ>�>Й�_���Ca'FLkuGd�ml�L��Z�O��9B��U�����Ⱦ��������N����!������X?�J�E���E���1	>:�4��x��.������ i�.�,��#����1ŕ�"\�]Y ���Ѻ����i�KqD;�!�5�v�g?$�Ly�x��i�P��xUe�E,��}�P�6Ľ��3h�Sv���E^@u�h�&a1N|�����ʹ
��?4;��T��%�5���el(<CT����ں�kQC�v�}Y����"�v2⅛U�,$d�9�|�S�Q�tJ�M`	�?�{�>��ʼ]~��wM��J_[!ܹe������@��b��U(q��P^�W���ZK�3�z���d.���j�����!��1�D 1�`͞�0~��Ƨ7QL�A���q+ln T������Z�pD*�9Wb��#A��idLcC��������?5���\�1cByW593z�q���:�u����7�f�6��\+��z�+��* ����=D&�;8^��'��V���i��(�\�^��i��4�u��A�T쾀�or��C*�V3/N�BS�J��me�ȃ�)�l�*��qY)���%c7L�i~g��ѴNj��"3JG���x�mV%��#�=u��-V��a��q�g>۳^����ո�t�H����D��`����ˋf��Rj����yD����DH�8\J�k̽��c+������^��ok	̇h����Fx�I�?X��0%���p/�掟�RLo|	b��Ȥ�ӷ���(Q�u�f�5}�&&�F���=f�P�mBD�Ր�����������"%]�Y��xۻf'�c,��l�����"[�щ]���Tb�V�b����Ȱr�'5k�ï2�D�
t9��]�қj�L�^P
ǁ���*���2}��ٍ��fL�i�y� q��ψ.U��Ux,�xy��}/A�����Eϝz��σ��?!�(�T�Z�M���9`�,;tK��<�l�&��s��۪�V0�
�Ɂ^��W��k�ۻe	��s��&�6�nq�i�m�R�25�cz�=��酄�SݞJ���/R�9*rZ��[L�E��9�V��$PXr��d;s!6#�d�-�Ɣ��iM��0:�NY-��k�Bpa��9��oRl����ݜ(
���z�Dk�T������Z�W�l�⧓�~�:�W��ݯ���o�+�]��+�yB��0�Hj'�4q�m�eޢ3�6�^�J�͒���ɍ���D�1����V��)6��77N�V1?1��c|����[���56�8 q,Q]t6֖���f����q��?a}֒���Ř�Y.�>�����}���J(��k�}�s��>�t�^����[��4t;�cD�{���LD&ޱS-��-��`&U�	ƹ�p�3dK�����M�����u�����ʭ��s���x�_��X֘��#��ͨ/��'h'Z�^�������Z2���� U����L0nc>���כa���)�(h��퓵$�6g߿Q������2߯��}��=�S�z ��P}����t�4!I�B�ʊ�;�>���wzF�'��|sXM�L�mj��~=#�&�ދ�gaqz�]���+k`P�k�[g'��܃\SCH��M^�TP�f�5�����Cgm��v%�n�-"ĥ6�=qxm���w�������P���~��&|8 "��o���}�,�_�]ˑ��"3�^��ַ*:�m2�d�8��C�[�;0,���E�n.39Y+�Tɺ�V*���N/u��0��ז^�an~�st#-���@�lxIIf׮K*�s�u��l[�W���<U��}��k+Gn]O�=(�l��݆�DJ3 ��$��x!�Bxbؒ�oS���ֵ��!�r)�lg�_�>>������_�>�� Ä�D�N��S�!H��&i�{|�>Bm��e���ӛԸ�m`\;��Q�ؠ�%�\��'��9�r%)Vi]�xv��{s��iY85�{���Y�ʖ��.�I1�8i���V#�D�ч
����0�0�'*H���~�6�~�9�v���>h����u�Ĝ{���y��G�i��	l*.޹E�K�;˔����i��s��/sy��|d%��۸l �E�ku��4tI�����Z~9���Z�a�ol�W��wwE�����iu�n�l{.�8�a:���d�u�{�׼��4&*pLEͽ��}z�C���x,����ʆ@��#���W�g�}C������C���0���P]��d�OM2��� ��슅^|�WX6&wp��Y��P��_��<�-�c���Es�mEj��3v�5�GC� �M%�$d�p9�E���wvو���Q�$Q��33�=4ͧ7L��m��΅l_=�UqT�m��y�:�Y�S����	Y��?�u��~K k¼4Rک�c��T��"�Y�_9ha����<�q��u�3��aF�5ygKy�)UZ�^�A}�ȅ�8���l��6{z�E�6��6�9N� 9�MR�����倗�#nG�.�L�cQ��\*�VA�[���C!�\ b��{��zw�O���h�|�!�C%���f�w�3YH�����w!��#�;RG�=��-�˟�SU�<���V2�����MF�^�6���Z���`�m��z��Չs�8���S���p=�wb39Z�T�5��\���5-k�3z�Vq�T���9�F���L�`vr�����wɴb�gi��1J���W�B��Pp��x;xPr�j)���kԻ�4˶��y+�+�N�Zl�%��E'�֪��>Tm��TY[vx�[�!zU��q|�B-�BWP�#��:�!꠾=v��Ҍ��G�ߌ��WF<1��������8,���UW��(zB�9O��P�8���w����]�ff��O�U�/�h�=��HK���h0��op���X�P�J):��P��8�[|�%��k��<Ŧ܅v��K��D>J�(�?|����'��}Йs�(��x�����Ɣ��^V*j��2�C�8��-�@^C�u�oGiƪ�>�x߰�T�d/>߃m�d1��	��ɳ�����m����ٙClw�k1V��Lڬ����}C�A_�T�Ծ��'������`�_���ٝNq<S.~�	={���L�LW?6[���e3�����jX�+�u���G*OovL*�GT��[֘Y�LSڊ�]ctsm+\P�����a� ��^�����EvN����lP��_���.�ɇF�k�6YN�s��`8%o"A�<�F����nLd���1pdg+�[L�3�H��K�(��<����.��Ц7�Z��gd7�����Xksej7J����S�+oy�]i��j�⌕��uYBj�8)�ns=#ǃ�b|�S���9��]�N�ң$������c�z��_g�i�����!�*a�a�F�M�a�Ć�|�5ù~h���n=ї�pf*e �j9�?s�����e�p�\:�Uܤq�N��y@?:N�����r��<G���s~��S��,+�d⡶T�ȅy����u\�!�Q���$'�`_[�(=t�Q]�F��**:/�[�����í�k[/����z��YV�r����j�p���|{�TZ5�UJ�8�6&�@f����>������Y�ε�7��tw��J�c��5W5�����0����*��T�?N�Gҵ~+Ο|�z=���8�z�w��5�+��S�d3V��1�����K@�BSlyM4'�t��U��]]����׷�]����F�0@C�(5�/�����ږ��{�9NCf�BD��η���p���s����] �,iߵ8�X����f�B�mX2�_%T���(Jh�6&�iO�
�3Nm��o�;Ѯ�O���
בT3���]�;�[7��q��t>�T���i�t�ƌ��'�1�^h��뾺L��zi��b�om�*J��͕�8O�.��*�� T;��U���ֶl,����e�o6�uo]ɳu��j���~I�/�vw#�ב� ��,�[^3<�&�d�QV�A������W-rյ��|o��b�uח[J�d�Mug�f�	�cK5+yF���/�Թ�U��+�k���n98h`
/[�g=�n�S��{S9�w�QU�޳9�s��#�&K�������!짃J��.j��W�:&�wD&Y�*�E�iU�o2m����`U�:��р6��mޘ�7v�����;����!\�k��{����s�<L	��Qn䦇��������g�4��GS�
��Bp���O����B�dЃ�� ���wE�����K㫛Ó?7IR����9va�D��)���9���L3��*g�t�"�P����e>��nެ'(EqU�}�Pi�]ф��H���N;�Oe5�`�ˠ�1�Rv�h�m��3Px\�T���ޘ�ܽTZ��P�h8����(��$�O/���-�aӖ�r��ʀ���������2����+"�G�㺞:&�tSQ��mQ0����j�k �M$�GAnʵ^f��kW�v%�71�P����`=��wţ�y�/t�s�&�o7�:�=k�tm����=vϠ2#+Ɯ��l#�:���F��T���-���U�K�;ut$�����;��cZG���3�Ҷ����%(!P�`�j���v���d<-�yN�,}ܘ�0�'e5z\b1C��ݰ�>��L�~c �����N�s|i�.�����e��3H���9X8�!2+��=綦��Uη�������J�ҷ��}��A�%���btN�~(��<��:ўX��u씴:ȷ��gwJp{��n5�>���.�>�fd���퓛�]FL��s>����gy���G�o�S�B� ġ�l�D��z���w��׿��<��
j��^]��;�`k/`I���.�{%dp̻�>���EU��;ߍ��O�Z�vM��t
�e�M\��9U1����B��tqTZ��8�t������K4t\ժ��cl�u�5���=�3�O6	T��ߕ\�e�[N�VżD�ӛ�����|��,uʗ��[I�h�W|����|����,|�A�H�ɕ��M�d�V꜇��pˢC�ۯTWs>��"���e.�)��v��	���Z<zފN����\Cf���� f�����5)C5<k�iɛ�\+�O(l���1n���.�C ��U���8��4��Qi�熪�;SrjUUB��nkq�e�r^�c�a�\$���j㙠���;YՔZ���k1l/�Z̙�7��u��\h.u�$wu,�a�[�Fz|����Pࡱ�*}ȇ/L{b˜��ɞ��T�uG'V���61����l��ýya�>u�	+��2�^5]鳼����b6���D5��t;.E5�0�]4s�%�������γ<�;�s3/w�E��3�࢘yV+�g�~�s�>;7��z��-D'b�dRfr�Eh��ӱU�(�ЃvM�*eh��QK��&��Q�2�Ӯ�lu�s�A�ls2b*wG�%���n]-n�O�R� ��0�"�5u��a�Q�;��'(�d��WZ�
�E�}"U'�9�����qЫ�Ӿn�km��}�ojj��Ü�MLT2u��J���n��������w%��v�M[��Gy��S���PJ��K?�(ba]%��[4ܼ8˃��ɹ��E�m�o��] ٔFޞ�0���9\�`H�����w;n,��]I[��ղ�J<���3������B�hE��@��=-�X�G1]Y���i�1�a���D�7�&/1�2�1$m��y%m���4q�μ����TL�N����$�&먘��4~�q�֝�tF#���{�NOVT�r(�v�� �մ����3/�P�)G)�kI����d�lۼ�)v�&�Mղ�B�(CQ�9ݨ�^����t6�^f<hl�m>���Z�]�B�j�=\��Eg��=w`��b��+뜍$y}:j��TT����'yn�iqˬKV-�krX��u

�:������F�y��)t�e����n�q6��C���[���os��!�YҔr��6�"���M�}�`���	�&�J�a���S聑��Ӭk����"�t�!�8Û����S0�q�oD��4b�[���Һ����R�����8ti�����8Fi�0�â8AiàÇ�tpç�՝���X+�/�]IVi���I򭱋]����$~��[��l�/��R�w�0�R��f����b5�����{ki�&�x�t�, e,�B�~9�t��0�m��B�=ag�zf��t>�q#�e�)��-ٺ�T��-�(9�WP���n�K2�k��F�K^
�x���.C��JuthR��3K������*|Pfp��
!k������+A��x�$A�k�;[�Ѩn��]e�&,]�g���w�����kkK�o=r%���k��ޚAL���ym��R7yIō������xZ7s3��t����!�-����x�qo����$�����Y��ɓS��ge�n������Z��r���e��%`�A1��N�+P��\���	�Z��eIٓ�s�b�c\���)آ�cu���:j8Vf�j����܉�JZ�ɓ�]BLeٷ��]��Z"^��s��J��܆F]�u���{o��gZu���t!Q�k5��x�g��jQ�܉��$�)�u��ۄc�GX;�b��|GkR��E3W#+
�����^L;xFGɈ��B�2��:�c����D��P�����&�|�H�=�tEa�ed�4�R�Tk2�"�٨�����يq닷hK����K?ZnTW�:&;Kf�J���(�_	un6���.��v9���c�ޣ[51��M:���ou�}�3(q�j��X[F�'��e��o�QGsI�j�ݙ��ؠ��D2R��Xe����9��ϳy�ó��4MMRSFYF�DQAMDTQʋ,��ʙ������O�^TW3��f=ɄDE�E��RA��S�15��8G��OON����s��-f)�?q��(s3�&�F~���fD�����ã�����vd`P�QF�˽2b����*�&����*
&�
��2cH��gǧǝ��rJJ;�(
is�9U4�Es0��Y�CD��)WX�IRIDنu�ye�B�e�A	1DA��DUws�P[�E���
��*h

�
�*:�H�Y%QIK}�L��rr���"�9����eTAE--!�D�{�(;���k� ��2���hh�(���Og"��S�L@Y���\̨������3��D�^��C�T�������g1*�q9��*�\S��Ub̭N���X/V��R�i�%�����̎mԀ>�{��������:�s�
��$���� hA)������_�������і�^aB�I���<�^�l�.�)�j��{g�pv���'� ��}�pc"��`�@��Qz����4:ؙ��s�Գ�FPU�7|��&-����m�'�Wz:���h^���s�d�р�he�p�a��~��{c�1��qvnLD`�n1u'm����Z��fl��&��}L��Π;>��܇LU��=$��W����}�XoR[��]���k��0��®SzhO��}4��|DO��#�qm���$%VS��f�]2d/>�D�,����L�� }q��h�:�~�!i�S�ʯ�v���Z������[O:�wH�3P�/aP�yJ�õ��6����n�C?Dp��j�m. ���nU�^��ߺ��.�&�Pi��)���+^�P�z��O��r'k�c
jx'v��������h��[��*�ύ��������9�����v]���<&���	�=�QI����5��Dzb[0U��{z�A�
��zr���C���޽6ӍS8�,��S�Z���'�9}�Zvاs��9o�^�2
zT>�^����3��뭩`�IJU�K��9�ې��H�X����{.̷ζ���Z�׉6�^+���y\^��T��1ҲP���/1�z�Q�8��p+��]���m�ǎb;̹�I[�]�\q�{�0$�j�����B@J�B�B��xy���������v=�T���묻��=�+e�c븦^�F/�R�'� ��,����&�Xv�z�!�.�v]�)Մ�M^]�O�i,���̘���n�#��3�~7��%?w��y���ʓf�EIdp:4[��B��
��ﾡou���m��.�ݸ��<��`�����s��mw/I��6��XH�dq�����v�jB� ι���Ov�vt�4�M���%�X&Se�{��6.��P�moR���	W!AW�w���vE�[��3�+��?��L�<�sicy��1����l�����q�V�Y|��3Q S��Y[�8��cy�=/�mjc�`�Y�����d<��L$@}k깦I�e.�5�x�y=�:o����1���k�1�I�-EG�=)�Do�DiyR���W���|W~��Nca:w�������{7�����~,�K>��UI���^]er`������j僕=������yw&�)�E��~�)�j�Nd[=�S�9�x܌��7����B}������N^���
��\��}���^��I�pf��to���Ӻ�ώU���ZGrx���EG[�wj����{O}����ut�+q{&�y9�Z�5e�X�N[G��:V�J�G��Ͳ�k��<�K�so/f��u""����tys~���]���A_�(9� �@<���x  �2��/S:~{�!!����E5=����R:���a�`M7P�$Iw�G�w=�ǽ������uτ-9�ȫD�Ϩ�2���0\dz㚥]U��cu��s`�fM�����t���5��el޵��V=�C�ɩ�.���A�.��@���.�z���sU�J�5�ˮ�6n����7�=�Q�q,n�����K2��ݧ��[��|D
�:��=8j���O���_U���nQaC�,�����ۨ,��DT���1�����5{O���gG!g�#�MTa�}A~��tZ�Oq�<�t��$�I�QUm���s��$ͱ�� O{�WϦ>��Y���� �>�O�89n�	�ɐ��Qp�T�tE'氺9�Y���Z��D��DY}�g[�Y	Q[eU�֒'�(�F����x/�F�U-"�S��Y%�E{��O���ϝ��os�����hz�̯AT�?PwN�3�phLs	wM��4�wg]�%q(�:hn5Ë�D��'�-Cv�����A����r����Ɔn�~.Z8�>��ɠ}�(<f/���oە�%\����:]�1�/���6�Ƿ�-���AB�N�������a���\#�>*�����^b�S�:W�m��=u��Ow�]YbˡO�R+�;h����j-[*���ǩӆ&fVwmU~z�l���w�=ၽ�=�R!T�Db@!���*��'W�kC}U[_���.��uj�?�S�oD�dw�����*Ш��>�:�-9O���^��k{mo:�kr���c�F�
�Չ����3�Ǳ���O��ȲǨ|�oZ���B�mo4
ߩn���z,҃t&ã������V�!����`q��w=Ø��:D8��cs���ݜ�F�Ph`�D;o3�cz����9%�K�*7]�On�v�;�S��`s"[FrZu�;�N �4N�[��k�C���FW�������1�7�O��ڂޏnk��`k2F>��u�c}����r�q9���E�y�Q�_���Hzq�3ۗ���0��QT����j�|S?�|^����k�n�h�u5�;Z�y�0�6x����'�JfOI\�b�a�\DO����ס�C�"�0T%��v�9�m��K��b�.j|:��*ֱ�2j�ɶ�Kn�g��I�<E�����W��&�q+��+o��l�^��vk���f�z
�����]k����@��Nc��s��%����ν���e�]�^�9`4y���R�m���ӏ�#�
O8�+_�TZy����\�z3����J��Wn	߄���w���:��ܱ	x\�\�ܧ#8�,�8���p���Z&+��5�w�:u�ڪR����4�\畏v_<{ύ��5�6��9�9 �j�8��KvR�e�M>����q�8�e9J��w����:����"�IP>�\!A��� ��w�����w�Z�F��27nq�s��$��O��'��_L����u��n0���$L��2:�"���*�b���U"��iT	oO��3���< # AϾ��}N���Θ�3i�w�j޹E���F/�:5��;`ؘ�ᵆ5[ ץ��h��P��iq.��<��[S��*�<�4f�
𶱆��)��F,Ng�-�+;D��tʕz㾫��?�엩�gX=�/产�y�h]��Ra�1O3���g�t*�:�,�rפ�f����|��Z��mxQ�c	��!�y�T��a�Ǥ��dv��\�#"�U쎓�iC��얍��
�[���^&,4s�`���vl�}�v����	��d{�r�D����dKכn��U�Z���x�@ɘMJ��>/9BW�*ZQ�V~E�Y�~t�VK67��i6᝱S0�a�^��h��6�}%�����0�a����ޚ�C�q���"!F�؆θl��*�u������R�n��@���mn,�|Tly���+�}}���~T���ʇI|�?
�/�>���)�>G�'���]r��*V�s���^�8v ����r��/��:5�t1�]�n������/8l�j�eĎ�\g._�z�0{�LYs9����M[~\j������܍��qt����R�F���٭h9�����9�y��T6D?�!����0d �(�(�J!H��4�%'��ϼ�}���>�l\m����-��p>��UB�82���҃m�|鍕��"]w���t�^\w��wS��z���e�}_Q�\Jݺ�[s�[�xP�%+_9�eE���ie
�Ӈ�i,3ט��ΉAP}��Q�DG�[�P�N��s˽O���L#�Jln�L��ˆݭ;!?45�m���n�$���)�q[�*^;��x��i�ơ�q6噽���Y��M��Ŧ~���#syAD��O��+���F��r1��h�V����z���;�o��a�V�QYo�l���F�3E�I��2��	�UC}�~y�yu>�b�{N��2d�6�C�=�`����n�p�L9��� )�cO�	�֔����i0�MJb�����~�m��i���ߕ����q��yۑU\���Z��<Am�. �����o<�|�EV�.m�ŚS�9#%��2��wUs��Qiq�`=�=����O�̭���f�,c�b5��fsb�}ӜhW*g�P�=�%�2��07�Уƽ�lW�����W�(����&cS��S���,<�=���F�u�v�9�Y˚�Ҳ��d����eӀ{���{֩V_�J[�s^���/{"�Z�׮֣�2ݜ�t���;��r�ġer�U���rŴ]qJeB$���=���5��yv�c�����k+���I]On�=+wd&�to��u�?��7�MUL.��`F��x~ox��T�U�G!�0�L%Th�B�����}���~���݂�-���{�UM�^��^�v�]PҿQ�:.���5GE����}�NG0aO]kLUpX���Z���0�1�NL�\��7�+�SCӕ�-�}�J���'ͫ�dmD��ӳzr�K�%��XM����Z�t������4�����i�UE��0���&�l~�ԝw�{��wc^}>�������ƥ9�����n�.���5��8��3�VL��A� �1g����_�+?W�=?$���]#�@�{7��ӛ�M-W�XÕ~�ޔgm�V�8��WT����ZF�>��+�����1|�*_�ȴk�M(8��H0 FM���j@=Y���^�TЁ���\jD���yCTC��|i�����ڄ8�}��T��{D�yK�
i�7�(��sa��b;�C��i������{亻����~��*�P�p�W�X���{8ƌ�2�K�!��i�<���s�U2�:��yfV0�T^L
�h��5���I�;�4�S�'�|�0���PHu�]w�Q/��,˒酥R����E�R�:�J��A��C�J_�1�/l���֐
>�w�y3E
��zyD��w�U� O���m�c��kn�o��kK�z40]Z 7���}�{�Y�V�\�Ðu�c�K�����Uk�J��)>��������_sI�:�)_Ud:��t͑���T�@�g}}w��>���{"P �TrA\!" �H� I��:�Ww*k��8���mBK��O-�2hL���6���Ғ����7/�S����Q�s�M���0}��>9F@��x�"!>�zz_�dK�%���0�ɒ�
U�]螁`pݦ�=�1�Y�8��~O�ױ��/D�^G���Z�wsn��3^�7~-��ҽK��t��=��;�G=�b��C��i�(��sO����3�;{R��CL�G�<S��my��B(����r�}c�*)��9����aN��
9��O���UkQ-��h2�������e��Hx	&�!ګ����F��y㟋��U_r��)�c�o�9�#Ŀ�q�h~m�4�1ԑ���b�Y]��	��z �nt9�|/���r�����Ϣ˿]CF�~Jn��Jz���7}��"��F���_�!}��+�|u�/*���@��^ݔGw�U�*'�������7��{x��e�׼�(/3eØ�����:'�P�qA}U��L����qK8{�y��4Ё�W*��v��d��9=;i�G"��5.�y��t	w���Mm�¬m��Gt�c��) >�ş�$�ome����;���A��vvmA?^���U�O�)i˽<���L�(�K�[]B��*�q[N�����/ne�{��g�ܶ4!sz3*bX�ϧuu&��=�3�$�O�o���f�A���~����w���!�!"X��DC�UQ�ó����.6�Z�e�߅ͰS�&k���,�k�Jf�U?}��3�ƅn|�$��o�#�}G����vu�<�z����9>\ԅZ�V��B��ɢsΙ�-�mK'�S��Ƹ.lK����+X�}�ר'U����5��N�r`�k��8��Rt_���hiqB۫]K���*7�����t�Q��oC�]y�{�ӽ��{�;v���Q�'aI�:$��Ug9B���F���w�WϳJ��R�]Fi�1닗8��>�����j㙠_O3��`���K�®2�6;�ou�6�{|����Z��MІ��/�4F84%�sЗ!y�4S5�fsl���.�\�i�,��H�3�C��K����?F��(��!U�!�矫��*�Y�)Y�خҥ�K�K;uԉO|�Ke�G.SI{�FK-��}h<���cݴ����]�(h�1����c�Wjz`�l"�/%�{�/��q�U�U��7h���6=���@O�<{�hO���.m�r�Hs���0�K UC��]f�<��hx���4ŧ���c:����h8�X)��)l��U��#4�8�ֽ4,�ӵ�b�s�X�қ;�(\lV�3i���=��R߽/�������{�M��Qvd�۶ޞKZ��r�wa6D��'-��13&^�D�Y�An�ȧ��}�}Y��u�63�ﾪ�
���Ģ�J����` �f �M\�����ߥMk?�~>�����F�xnQ�md{���X��0Mi�ub� 6,�s3��wC���3e�&Ũs˾���8v��R1T����E��KE���f�L�ܽ��������x�L��#({��/����B��g<�R�k���sKR���[���K���y��7p�d�qa:f�%��%S뢝�mQs���o/U���ս��(���U�U������L:���n�J����=6׹H��]9�ev��⒯4ŷli�ٲ�������|�v����n��`ؔ�|�A�<�J(��`�z���̶��zѝ:��kEA?v�(���t�`���G�&O�/|�S��	�����s
X�e���tfv,cn�#6����J����Yr±�SE�����֨r�āo�?3^*E)�]���3ܤ��D)�@y���%>\o��Yw#w�V��k����
����&'��D�1����HkˀC(3�6�o��
u`�o��9�,�m#t7v�n�\?3��C��l�=ɖ��0]��r�;��Դ�RwU���V��s-SR��T.�{�ոp-w�ʼ�V���'�.Y��ݰʬL��bVD�8�+�Y�#	K�;��Yl[gR�i�X*��V�)�6�֬��$tn�VG��A�
�Lg�1��"]�,PD��gY�*X��1� 㻽���km�x�y:&j���2f��+���N�-Yբ�*�k�-�N����4U7���N��(���g@��aT+n�\}�I5RWZ����9XP�Jr��ݼ�e��5�R�=�1vT�)�I���4�9
���-+l5bv�u
	K\�>kV�}#�N�K�î��L �b^p������StH�I+�C�l�}V�������Ρ�Y�u]�6,��LPõh��T^��ٜ�ʂ�I�*T)�X�v�:�*]�÷�u
\5;J^�e��fe���˚�OaȞ�
�-��
l-�r�[���@ۺ��K���˘;ʷ\o-N���q�:!Ј��)���\{��rì��]nEd.l*�r�_;�R��/��	��l��u�)p������#�赹��+�me��y��\��um�4rv=yb#�S�jج޻�eK�q]a]�p�L��ՇU�$G��E��Zι�6��,Pi�<���p��;��]��R�w��j�[We��E���_Y�2Я3�IB��o�g=k=cV7D�{��a��Q��=zV`��Û��|w?�+�[�	v.�|ڗ�y
l:��X��5�[�5u+�Q��U���VVR�_��{)�8��a-�dz���}0Z��p]5C{!��g^.PȬ�W)-'b�Ä�:�
�R]aܳ��ԨT�������;�P�M�E(�����1�u%�8o;f�n�u+Yk�T�l�>q^R�A�\�f��vB����� ��a�#o��A�a��٬"#\g(���vtn�\Q��+뚅̽�u���)G�Z�
�A��sz��*t�ئ(�ͺu��]�� �za�D*��iY*���c�����%Z|jV��C�ϰ-6�Q�'�&Va��F�H�iT互�5�X+sk�䔜�Q�����<ܮ���Qc�\��;��j���q^Ċ����w;�����Y%�粻�}�zҭ�øժR+��'P6Lm޸e_;��ʈ:Û�+�nl�#n��FrJ:�f�9;wi��fn�T���*����S[ȕ^Á��aec˾��_�AyS����%�J��/,�WH�9l�� �^��:W:�A�p;Cq�+��8y�ԙOi�"���ɻX�����]h���ܷTϵ���Kov2��4*q�m^͈��WT�-�iթ7���spjLٲ����ň�s{�w�Ck�Mj�y�^��H�C��<�"۫�}nN�ڎ�LB�y�C(�s��c�����t��O�M�pY��{?���(~� �d�;��#-̪)� h员e QH�|F�~><=<��Zj�c�¡�r���CMMQFFDfHFc�Q�b|F||x|y��U--e�����C�HD4Q����������~;<+�>�E�$�	�`Rldu���a�T�PP�U4��<><=<O**�$��2h�9�U4��E�@P��T�M4m�񆈚�=# �J��S��%%C��-T���d�ɐ%4@U%4��e@��y~�h��(k�0���"�1j���)��S(&�K�@�bih�*2,̃!�ihz�/GY��w�g^�s�̂Nk���Z��ԋ�\>Ȇh���'^\<�nH�ES�wm\�4�����ù&�$��("��4�ח���}*'��\ �A"EW$R�i�>�=�?������;���K���<��,�}��3	�t���"�nSUwc�b���jT����\#�~��'þe|:5^�+��U5�,ҞaA.�n5{˞P�s5`4�u���丹?��
 J<$�%�h�@'8*=�/�ػ�C�xy�@�xP���k�����+�����2�
��B�a�E�Uo�t~[�Sk~>���V&)�CocT���l�l����yb���H��е�t�����cA{��q׌�<?��x� &P���&Y�:��m��s(l+&�Xפ��bb�Ɓ�1���pXe?G�<�4=+��.���=�k�/vַ`�wON!
zQz����m��q�ks�4���,�\[6%TZ�VU���Z�_���D��_N�r��6ɕ3��G�bЬ�H�+�ƻk�3%�F���`��^%�`Uno�&��%�d��ɬY��ܥ� ��F=�>�1��/
h�T��Z�c��v@��;���~��'��w^�>�"����Ȝ�i��$�;	������8ׂ��=��8��R�����y�ݪReM��:�7���:�E�����^�u<A�c1p�q�ƶ�2Q�;�x��;Q�d�)1�K(.�/�P�����nV�q�ha�U�]
�O�����<��a�H�w�VJ�u��f�X*�w:�s��κ��P{��� �B Fb"(�/<��翻�]�jo�s�����&�0"��yCTY�D����=�@��3$�/�W�b�f�T��\u�Y�=�;
i��2}�4}9}�O§W�o��7��Oк�R#� ��_z��0�����Ơ��>�)ےh����a�ze2��UL��SmԳ+QQm�����dӛlW,FB8�9�|S�<=�;��u�C�Wy�yg\,V�=���In�J��W2�/kkg�Fe�]�bf5�s�1Mr�[Pw��BR�S�+���0@�d<��H���7����}ve��N���꨹~2�-l�M����@�y��n��3�:#�4��ǝ����;~��Ic�[Gd�S�!���2�u	=�:����ۛA0�e�:��kۆ�O�ϩ<������]z�\�Э�����P��j������C',����m��������hF/�W�?7���DO�?VE��ѽ4���YNxŷeZ�3T�U�\[%�ц�UR�&�y�-��\���f��{�V
�C>-�L�2�������*���d�s����7�>A�<�l���!�2}7< �{o�C묥L�ǣ�YKavؤO5�uw���A�z�O��N��̢���y*�B�e5F���N��A�V^�,FF17ϊ��X����u�L�e*6�V��6U�*l�{;P鞋SqZ�����*��xt<����|>�N�����y��|�� ��X��X�=�"AB��O~녯��O뛻�'���ڻؗ��������mz��V.5���iw]�jvX�O�j �w!�A�-@�Phowv�a@b^/�xc5��Jx��J핁�)�fuR�L۬�4p�ݤ�_�&�&���;���m|s�9�h�D����(:F��5�!�9��3N�V�^���lQ��hN�_(f��#˭�<���'���w�iai�Ie��u�}�V�c���?*t&��w�l�p�z�C'�*K6�%�+�j�K?rĭ���zq���WOBeN����4��`�sR:���\�5�d�)D�l��U6ߒ�ֺ&��V��o0
M��e���X�������w��6܌��N�t��H͐z2$�����R~��v����G���~�R�1�˫"���-������m"J�m��o3@����8�a;�0pg���5�.��W���/��~��mk	bj����{a�SO��a��x\s1�yMa�
V���Ģ�� K��آ�eE�I�s�P<�-��%]i���2j#�a>���PV�EZ��-m76�C�� �'9oN��jv�Z@viy��L�kn��l��3E�ڀ��|��_K;؊TN�X/8���Q�Elg+#��W:�	/y�c���l�#H�)��%0iR�@��w5�}s߾�{��o��]}���_�#���H	��
~�}����������w{�!����p��&�E<{�����}�(�`Lwxg��Q�1
��ږC�V�d����z���u"y��"��|d��9r�K�`����	�"���ݙ�6���1�:�����K�F	:N��z�~��a\T��O3�������o�^L���2̮��P���Ol{�x
F�@�,WC���s)�	1x��o��G�h��1}��PӼ��J܊}&�+�x]xC� f�3���A.����O�,����p˸j�Rڰ��&�	d��,ny��;��&f���"9��%�M�d|h��w���<���5����2W�b������3�����}U�e�x˵���SW�E�'�yw�N	okuoc3)�6jeF��HDdS"bا�*?�+#5s���O�@������p#6��B֛�S\�2�/���j�����.2:�
���2�8�����C(y�*f	�ܨSed���/p�S���egq管*!��Sn�ӕ���JETg�@�~��ya���{Ѓ(}���~�ڱTʴ>K0ơN3���N�5�0i�f��6���u*�iU�`-��6]�֪�N��J-0�n*Y�WE��R,:{�yEO�b�b3�vS8��e�`��ؚ[�J!�p'�AufA���v�Pi��8
�y�N�˾�7������9���w�_��
DL�J
d�P�?u�������ξ�w�﯄�V����a->Yr���λ��m��q�!��5R�yݩ��2�$��6&/��7��Y��\��)?b���u�깆y˨4[z=����)�a
ť��{u�`�]���u��L�����k)?g��.8�V:����[qn}w��S箐a���ӽ��T^�K�۵�h�j�Ri�t�N�<���J}��G,l��B���5�5��7�3���V����O��1O�\��z�<��`>�I�+�Ԧ)��\_��j�%:�|�<��p�ݩyڅ}�k�^Z.���BX>~˯���r��;]��{<�P�j���e��랆96{���[Wߏ�𬯝�,@� W �}hUK%�.Ͼ>���skk�ڴ6u�����������	�dw8�JK�P��9�k�J��
����E��^�'����%wA�TУU&o0�oq]��AۋO��~�cET��X���(w�CJ�I��x�lTse#
�y4�e�`�=2UsM��WS��b��q�kz ��x3��	�5�!���Gc^���sFN��Y[KO�A�,�;xu��
������q�Ѵr�TE���9�Q#8^��ΈcI9yr�LrF�k�A��Ԡ��+kN�n���wO�6��[�&H !h;�gS�yW�i��]�v�e�7Ҟ��Y�5oY�UU(UJ�$Hd� !���>��f����s*�&|́�u�oTf��pq����r\[7%T[���<�֦�W���Y��:x��P��|��[��y%>�ͮ7ٗ�^����^16"���s�#�

&�vle�ȫ�d)�2WV��C�*�c��^��UV�3���|�8����Cɼ��/��A�]�^�|���?��v��9	��	�\8|�u:�<5�9OmB2�	q�Wc�yI�����O_<Q��MH_���"A��	��W*a��K�?g�.�Y(8l��V/�E�a>k�g��l-&^'�A���e�p���6���,��ئ���N7��U���6]qD��_�nXK��p�X�|U����5^:�����u�k[ �tIa^ޙL��e�uE6�̬`Vv-�f�u!Ꮯ}n9'ز�2^��]�1�BF�>�=nC_t�Ru���%�*���y��u�R�B�z�sNWZ-Kڥk����|jŴ�h�g*��xBn�d�d�yƐ��fnǜk��V`��v�N_j��\��G6�R���80�h�+C?�����F����Mg+5�=��*Tӡk��C���8\w\�)�sq��'�����g]ؤ^@�+X/V�cH��5V�}�A���5+*�P�ҕ�	��[�Ÿ��d,�.�u&m��M��:����l�
ղva�hk�OC['>�������-W����{�?q�Ӯ�����(�	�	� �� <�<0aUN��)uB�7�{Jס	U����=*�`'��_]�eԣ@��/�n
��|�t�F�#�r�s�r��+l�ɖ�t���)T0�0�������ç-�Z��h�ͽ/Cf�ۛ���d���ڃ�r]	y�MR�hkw���,����_����h�ጱGqFM��Ѹ���wv��
 s1Q��_x�G�u��*��	G��2Wy}>���e<k��F�����j���3>�:����;k��c���!F�����b��+Y���6J��R��ܪ3n�q��&h�A���b���f��(-"VIj��¢��3m��,��V�-�ދ4gt��z�Ӷ�ؑiO�m8z3U	���Y���{熙Q�vzZ�ܲ�#��Y���a}±t��^eT��T�T��^��cH]o!��'�}[�:���"�e��ԃ�Q� !,������x��7�g�J���0��J�̞�������⋈���lvo�޷D�?��Ԝ>$�?U���ֲ���09<����5D�{΄2��Ĳm��H5��]y��>�F�Ɂr=.�/��'�>�����$������n{r�AJ�̦\���>gN�Gc|Ub�@E�
�Lk)N�-]�y�J̼Ǐ�c�"h��IY;^=�n�jD�A:�G�� �ۓ�_ֶ��v;J������I�`DcaJP)s��:��QK��3���H�D��\�W#*#�ݮ��/H<�m�oE'\�SMX�&�".���C��6Wk�0%�X9<�}b�:\��zr��������䝚(l����퉳��љ��k\"��r�s�DϹ��OI���W�n�Z�a�@����v=�A�`�)��?N���]�[j�c�2�����ʔ�;N��p��TR������^X��B���1./��0��{���qj�t	��_<4��xlk���yD1&�s��}��ߟ[4yc�L�w|a������ ��nB�ޱ_Q�u�����O���B��0�n�4��$�e�c�[��n؆{i��}��-�6s�Vq������>���
�˼P\~�چ�q7��W����-F����x�٨ٰ�6�i�S�g��<����?�!aU�l�;.C��Mz��;�2{*+�7�;��H�Yŝ������T1��:DeJ��%�3��E*��]�#(���r����2p˰T����5�xoC��b�c��3�C��e;׉��(��q@ŉ���.�tl�%W�i�hwau_NX���_3�Na.�uk���;P�����E��s��}~J6^19٩d��w��٪7^Lw�-�T��f��PAf�V����E�<�X�.�a�l2��Dcy�Fe���&!}�r��:枬�:Tu�CPr9�p�.0��[I?���~B�0��o,��"qJ��=���f�2ݯH�3�v~�^,�׸��J�-F�S�yw�hp�؃7�"�>R����/-i��yS��:<�n��5��<�ݸ���\ˍ��|����7*�yG��6a�XP.ry��-��Na���~a��ա��1ۘ5qv�;ݯ܅5$g!�w���]���\*E;٨/��m��S	5:�Φ4w�0z�c�J���i���+��,��E����ʵ�2ۇ�Ψv]M�L���,�_��|vZ�qh�l49yYI9_fm(lPbu���.{����+lgb��>�""�$~�U���E��
�k������pB�T�8C]3@��d��5�c�U&�	�+Р5���ho+���c�07��(0�r��B�^�����z�HA�Y��7]Q/��ͧX��"�?���v�l�c)�ZQgS��sU��$�oe����\A(��}BC��Ǘ�!�2�I5)�8఩\�;�B"�&�ֻ=�������zg����a 3��pv��)��w������:�����ʞ\�l�����u1��6/�q��_��awv� �������.'�U��n���9������sz[�n�N�ԭ�dm]%I�fVb�c2�@�L�9waђ�1Ә�Ot6�֐��[w�ڲݧ�aA�������NML�E���fm��|><��`�0����f���&ԓ<Ɏ�T����ȱ�a�[g�2
�M /��Ъ��Ul�v}����י�T�O1\�<wp��#�&�8��>��1���/�RXHX�/�C��oK��T��@:��|mq{�q@J�(�յO�F�S������[�q8�?��/P}?_~m�������o�g����ۢ�s����.0ኜW��0p����1n�;��[��q\c�ܙ�x3�(L1麉���tMj���(3t:�۔��Oޗj}aa��������0�w���;U=t�ԼG��^w��z�U|��w�����a�L?D�j��:M��ƥS���i�N�
n����}��J᡺]�ƅ��]Z�ԽŤ>�6��w��+�:~���b�H��*�N+����>�v�{����L޷�V7�}�(�P�L��@�]7����O�L;a��l��{j�m��9�i����`�[��[4�Κ���r�&��ʒ��av�RV}�*���p?�M���y�LK퇆����s^�����,��<��6��	q,�_��Gb��Uu
!mmĺ _���*���U��w����
���_
�M�
�,M 
������:\���v.[�r�<�$;g��q���le���sGV���Z���l3�Wo�]B���8w#�)��4|��
�/si(L"m��{ZGٽ��깩S��o#8���ig.=��{k��W�9q|L]��Ap�!�]N�]뾷��F�.��a��F٧�9���8���B�Ktv��:G-�+�o����K�f�����V�d�kQ�ėv~����J8&@�l�>�im
��C�>G:d�k�rҫ3rt&=9a�/-_=��3�Gw�.��F\�d3�NpGi׹h3����e��[��u���X@c:c��A��QrL'f�>8�7ս�c�Uy��`��.L�C�I�b=�q�	�Oku%Bԡ/wmR�z�{}��u$��uu����o`[��p��*=�����T��վ<f���%:�1+ )���epHx� �L���e\�Mv�Ll�p�[�CF��W�<1{�:�EJ�F���j�l��l�B�R\ze"z�r%ڕ��eB�oj@�����n!��5Ƕ<���E)W�/;.S���I����/%NGa���[��0��j�v�m�s���Tk�:e�8^��%z�T����uu�H��ێ�Q��.ܓ��q��EQ�t�:@e�|���V��W�5M.k;�Q��m�f,�1�A��t8Mdܺ��&=}pS�٨X��t>8.`886�\gw+u$e����L�JT*\ѣ�B�cK�.T�C�*T���K�.P$�%K�1N�?0���{�ɞ8��Q�`�ͱlL�zvr�j�Zq��/���$��uË��'H��@�=&R4c,G[}7ve&y��'df[�͠��3��vlRu���wh6�@��wR��ӭ�vU������	��J��53�'�5����G���g���љ�d�o�T<���ٶ���ĭ(@��]ݑ?w3�E��7j
��t� z�6 ��t��yg&��t���(�" ��k��uБM��m;^�|��1
�x8%��+0�3]em�w�)���;�������U`��x��J�.��P�nZU�k��s�q�ؗ��{��[�C곧u�t^,��c��G�r�U��R����{u�!U�dd��$�'��M����I*s�Eb�{^�J��9��^����î�V���nJ΍v.u��η91T=sF��BVuN�Y1��*˺a�m��aື�,ǡ5.�u�r1:��[	�`��N�&ԥg�8k:zh�Fw�]����j�kB�ՠ�������������b��Ni��(�Ҿ�kaݻ]Y��[�0D`:O	�`�Mu�鯪�kS-Z��V�e��.�X�)ۏ4�]��q�#x�Rq5�n�j9ǖ�O1��;�p`�U|�K%v�XʂX�3g7hN���x��B����RŬB���ۉ����pN���S�gQ��D�&�ξ�u�6�I�H�oowS-�7�%+R�N\�)�|wi��9�_m�d>G��UM-!KHQ����T%4�Q�����������bR�����*X� ɤ�)Z��xF����yE%-P%�d!AXF������HЕTS��B}~�E?B��� PD�)F�Ǉ����?@��%--_`d�%D�QE4�U�*X�����$�$�#�0)��i�h�(hj��biy	䜩
��L��q;�=��6��*��ʨ�W�!{�6��P��4�s�rS�J(vJV�[��G�r�wrz��n`Y�A�R��d���G?yγ���:><�J]8���\,q��&V�&GY��޳û9�3U94�r�l�9��5ϺIۖ��ד6�	��E��_���(��(�*�J:4�g���~J+��*'G${�P���͠o��XHޙL�%T˜��6�d�lo!���ndG-��'�¾�z�e�"^�%4i�vʘ	�\�F�0k��"�{w���mg�Լ�f&W���jۨ~�����uHЅQ0*^���>���E�!���L1�~a�ssu�)j��Ņ�F��y��AtsjP���T":m3ǌ�B}jz_��t�pw��:;<�cO(i��o/]��q
�OA�w>���Zk��B����3^ղJ7�_��J��b����T�`�"[6�L�O�M���*���\�y(�屐���k�m����X�\귦)��U�[�+새`d��<��^��5z^[Zcw�����~��Wߊ���C_{���.����SWo�قT�3:v�vm�fC���t_Zy�zO1�#Z��M���#ۏWX�b��.�V�MR9�!�Mzs�Y�5�>�Ba�`2��D>a�Raz�g�P�f7�|�ڇs,]��v�?r� E��<���[G��璔�@�H�m����d�qeD�7{a�����
����,���(�?_�,VWv�_��E��a�swW��<
LF�ո=�I�{��h��زe�uE3{�%��@���5�vt���:ق�{o��:����Q�4�OV�L����#��s������޾�����������H�f 3y�����rf��h<���H�9�6|KH�!)������<��M�0o�`;���_����oQ�d�iצ�[��|Z/2�[t�v�(��b�cO�[�y�=sӾ�}ڍNr���֜�B5ן`SLljz��*��`�{TW�2x����[�*%���a7��3"��TF�Q+\j��^OM�e�P����)��`��7zw$u�M��K&ٮ�����,��(�~}Z��C����l�P��_Q0��ث]]��"q͖�A��;�MȞrU_;�����cn�(��~�"���8��|lW7�쮚=����ĕ.�^���vTb�7.L.��x훍�vɵ}ή�:L�{J-99������	��mE��m��'SO��Y�,p�6d��xR�v���j~Cc���{��rTZ�����)>nU�_@�
�[Ol�9i���X+̉tr�1�V��q���KЗ�-l�k�]�9N5 M�.�'�r1b:5�#�S$enLby�c��Oo!n�:`Y���^=	yO��D��(�/��s�	��$d�V4�Ʀ��5ƪ9�Ӏ�u=cŸŶ�����Ĥ�1���e u�e<˃VV��\���J��n��;V��\u��S-_.]{m�l�oC��۔�f����5O�E��82����|�l�p\ܹ��"��V�W�0�@V0���ys,��,+��������
Xa�a��TK_�ϻ���~�u���?���\��>C���
����2���sU��"�ݥZaٷ@���{�/�\��\�g�tUsH;l����1�0��zg)���K���zO�GT6s��E������lslb�yA�N��lBΑ_��i���|v�E
�(o!ϟ��;_Z�N�uX1U��P]���%#4����]�<oО^\+��4�r���w��D�~W?��)��p�_��#�z�����CΣ����K�	���>U	��Z��X2r�]���]̟t��;�����|(���8���UY�7d�����c�-�i�Ʀ5-w �T����>{G�����9�/�y4^�F���_�E�TQW1Y����z����!�鉡Uo�v^b���5��'��z�S����l��������8��*˨�mASG�1�'��|�7J��.1m��5�1E��K)�շƵ�2뇇Ψv\1���W����Di[&���!��5F.��5�}�I��s�\��S��a�𽴫u�ުۖ�L�"���a#��i���oΈ�mk���)Vn���:N�1�+����TE��V���m�#L�c%X�JjYƊp���-T3���%�L)+͕ԟb�l�^ݬ�DF@J݋��ڑ��׳�9�~hF�t(�~)Z�u�����Eͩ|���h�ٙ����wAdco�<��37އ�gɚ���&؎�m�I�S����`�{̹��˞�-'<(�{�9���A�T�=z_�~��CYpͺ���S��)�?bS�"����K���
���5���Xh�����U��.\9�����.yCw=�'�0l�L	�L~:�N�?�Ø�.X��}����B\���?4;�}���DF7`�xM��1�#y���+缹>:�OO�U3+'� ��|�o�Ia>����~�}�Y�;F�����ɓJ�0�K���I��oP�^��4)a5�S�q�נ�;��PXH!s�S��vŜp��X3Mۿ��a��Ų&w�:��3��TS�E�C��cp1R_"�~g������ϥ�7¢�zy��ݐ�������Hq���>��ĲN�Q�irf��q����\+��6�s�{���(*���b��7_!4��3�ȍ#�*PS��Ļ'��#�B�?x���^&}��A�W7wTi���z�CY�5X��b����Ƀ��/ڪ�y�o�5)�~�ޑ�~�fX5U���x��U����NPw[wv�N�e�f��Rʜ9O2�&:���Ŝ�3tP()*%b}�r��u��z�9[4�u2@������WUn���2:)cs���=�K��L^�| {k�b�\�͚���f�̊k��)
��4��X�=�V���}_�y������Yj��]n���!��i$%6��r�hO]0��D��l���
��ME����xD!sI8z�xKÛ^���T��\�oCH*eC��9K�!���u'���lKd����ubo�R����w3��v<0����7�2��9	MjBmIv֣]d_-�9����>�͙��=�f��+ld3b�}bZc��
��6t)��w)d�c�.�1V7��Y��d Oi���ΤN�ܙ��ȾH���:7e�5��y�W�T5ʴ��5�nw�� ��/�lP���7�/r��������[%���|�G�����9MR�.E�)�kV�˩lyU�4�p�X��5:�|f�|q�����������mB
�mj����e�62�Gr�]����/�3�W�>�Nk���E氺9�����r�y��[L�������Cc2&l�8��;�;R�&�6�ԅ��0�G(E*�=��]v:����ۛK󻡪���7�[��E�+��S��+�,"ȗ�`�鶽���~��tZ��PԜk���[N�A���˶ǳ9�Ա������5� �<�%trag���ϧs�ڽ�?	�Ch����:�E2���&d@��ȵ��%����2;`䜗j�a�g�r��@����q����y�'
wW��Р-Y�ܲ��������⊣�ăZ���_W�_��	��U�e�C}��!����^�/<�K�kH��m}���:A`:���X.��E���X�rc������.�F77�%Z�:5���G�g�Ҿ�HJ�O�#[���uo����X�ǌ���P������d<6�(,&pߤ]_�Һ�-�]�x���ǲ�VL�~��t��K�x�%(!O�jDgW��Ahi�KQ>u�;)6bqqMyx�����g�75[ިg�0��V~��2��_]�"���0��)��v��%�����EU��?f�,d���UKP��N�@�A��3lH�Pz��������G����W�!��W������\"�뫟M׮m�bQ>��,�J�͏�+�lC�s�y6M�����'�~B��+I9��ZeY����d
k�@����	��ܝN6�B��N�5�[^�jՖI<�kɹ��Nֵީ�xk`ڣ!�����f�P@��
E�g>��}�z�¢��[sn9�ih�~�CTR~�[7�Nc݂�e�6���Aw��T;{ݒ����87�loDn]~������[�.�Oga�%��
���iܻ͌��������r� H�v�v��7{��j�,X�`��겍g�f��"�n0V�5�\�w)��Z[]�V����Ai�t��x)G�te>��H��j�T�X0M��]���-��z�T?~��xJ}m2Q�a�'�_D�Z�TZ~9�T/���+D���3ڿd�`�i�=Q>c��1����Y�����M�K�z�3E��v�⨵�QaDR|��!0�y��hr��'g:�],���9m!��DB\G�1����ɗi8z��r����]�m��5�D�Z.��e�0�p��j�IT
���]z2����x����~�q�^9r�S�ON)�&���F��:���}�����~��79q'?��tǅE��1���]ޕt�KZ�O�Px�4n��a�:y�=,��]#\��lκ�í,\����«�3W�L���<�
_�j�g'VC�9��`c\a]"�^��"MN�x��v�ݛ!�yݴ�G�\��ɥg��U2��ez}�9P��\���cn�zy�P)�^.��r���o���'_�����^{������X�ݦm�7�羞�LTx����P��"��(�����=�S�
�,��TU=,�Γ~z)�����*?��[c?7s��������EP�����ۂH�����Ė�Z��:�'�9�z�$�z�4(�Kʕ��I�Gx,��0���nJ�]�|�fT�;��8�k�w{�ծ����U��N���HҶ���/qڕ�(2����%Ԧ�ը��J��觪��vkgV8��|�Λ}C����5��T�̫�}�y�� ��;'�/�~O�"��~uu9%=K�8���>8n���:+t',۲�[f6�㘤4á�r�xN"_��tG�_�~��&�^T]oo/n;�b6��޾!�[fZ�9;���2�6������P��ʵ�)�-�Q�">�A`���	��������CfߣKU��{ dbyv��<&Ʈ�L��b�O׋(^�*�\]��jM�;j\ed�c�w0^GF��F+oVdc�8�[�h�8������2��%~�.9����Y�Cg�-�Q�C^�諧cmwwp�_��Ĳ{�
�ǆ!�nH!��`3@��F��`�V��6˟�^ʬ8��
��s��z�_e����C������1��r˞������H�ph?Luq�Z��:x���� ܚ���e��N��9�J���j~���D�3��,��r5��a|��^e�fg2�кz�j�^&L8�F�k��G�7�����-��v����C��F��%l���ߵ<���ݎ�ߥ��[�Š�J�al�:��qh�0X���l8�<uL��-�u����%��wbA�\f��<��{�\���~�W8�)��E����!�ﱐ�<�E���B��+N\
���Q�F��Jڳ��W�#����5��j�f��w�ϕ�S8�yM����3��&_��aO�ҫs���9�/�z������_�a���00X��iF��U"|�X3|��	���u�>��M��qX�I|���jf[[8�4iS\�=�ep�f��i`�(<��Hyc�����1�YxX[WV��TcS�F��^(���A��[���U=�����P�mZd3:y��>�<�/��H���=���t@:�͉F�R��oWq��A@~��U�:ޓ�W�uA�&�JK���I��x���?|oH�!|O=�ϟ�B����ͽ�I���ͻ렢86"�,`IV0�=x̳�����"Z/�XHm*qwR�ݑz�̆��t��0��wv����L��A���$N.����u$tö�x���,cF�`Ѧ��Bӽ�����:�	��%��J�����Jh�6jWU�lu��'qeD=S�)E7Q۷ܵߙ{b�Ƽ�A���S��cЦ�r�O��SL��V7��0RmŅF�+'r�d��S���D��8O�ٳ<�Mm>���t��kd�%���i8��Ws͞w�Ĵ(ݎ��X��Ps���^��j���;T��}l��W��j���yEf���|������}?::~�u�\�{�q�
��X���Ui�^�9/q�ݓG&�8�ڜ�)����$��^f��/M�B���L6�,��{�Y-뵭Џ�>�tY�˭����|�� �yW���6�h$�y�PY��n	"���Sx+K�S�߇�R�Rf��%Sk���5Θ`W�E������/aعA����0;��F��؆�)��G�K�����!:=���s�>��R�O��UyF�@\�m�R��X�����x�d.U��[nN�>�w,�-ޛ��ձ,�ײ[�ļ��*�:�x%�`u#����(�f-r���v*%z��^��kӘ��Й�8U/����ޜ��;�)-MCp�p�X��~nYР��vi��BJ�x�/��tCBv�b��hhzC���{��t�0�U@�3B�>�񊾙�kڽO�\�%Z���rgl�e@��2"�?>m�^�۟�='���ʤ��|�;*��Tj�-cuw=�g��t��55�&������}��A`�`d�^�bh,�!z[$��C,mM/��M8Ʒ�7�;��hp|�/�/�a���v���͐(-ޗ��˼)o=~��=�qKC��͝�!��vq�v��ωi|����5P���}e��7��*=���*r������@ݔϟ�������I��N�^*Hm�>ql����ۙ�.�R�K1�؃��k���mI����T+i�y��P����,}�\�,w�&൚�J���Q���[ոr�w^r�%�kP5�9�ƣ��Q����{��*V��r[����yf�2������ٷ'	ثR=��u��%f���bQ�D����j��͹�ʵ�J��Y �;r��}e�3���L'-B,p�.�0�Y"��7x���!1�L�+��k��آޝ\�+���-���N`�s�BB�1�y�k��0)��t o1R� 5vP2��OP�Y�&uF����g�N1j�76�&z��T�}�����l:Z���V$��Ɛ�|��u�Fg	������-ƗWo#�׶�6Y���J-�Zr��b���B��[c:p����7F�M��U�=±�P4��n�'d�۝�r�(xl�i������;�	�4:O�5*��J�l�9ř8-�qG�-Ghev%�݅x��N�oWwTg��/�ȪZ�H�[/L͠��J6�Y��)pd=�)me\z��v)�fz'ͷ���6KNR}���Fu��3��y;[��cc�ʸ��oa��b �s/f�X$Nq��w5N�8��u�9�upУ'w�=O�+�m֚����"�e�}}I8�G��Ex�t]��j�����a��|f�Z�զ�T��캐>ۀ��+ř�1A�������U���,k˻ZB���\$�gaIiWv�:�ְ%`���܌�I��t4�� �)^㔪�VVUӡF�*��q*���=�'@��@%�C��^�9M&]��}X�O_lL�	5�/�1�88F�`׉n�!��,�ee���:������ɴ>�g�����U�[v���d`��&����)������is#�{�󎸪{���in��1���e�ͳ}����}a�Y����a�������nIy^���tC�-��ۮFv(��i��u�7sVZLڛ�r�G9w~P@oE����!���V�-�{kS��GVwfΘ�U)��I�w��TP*-���q霞�U�QK	[�MQ<�7��_e���G
�����Hm6ǂ��S��K)�;6�ݨ��P�;lM�k������w��ǷCgg&���{	W�j�<��6�;��wF'�Y3U+u��9����})�I�XO;�2j��j���h��^�;3�(�B�e�y��sZ�T�r��yX%��^�c-�w�+�U�zV�V͆����C��b�"���Z�,$;x��&�ҩˇv�*���B�/��W#�������M�d��Rd��rgv�����Q�"1%VV.S8��ޭ.>'v��gKˡt���x��i�f]�N����q�O�^�5���.u���������N8��'����a���k׭�i�z�;���bZpi���5��'�p�CiTP��d6��E'&��
G' �t�O�Ǉǀ�@{9rC�<���L��
�ʁ�Y��JH����~=?�@�6+,F�)rO�yd�$BdrS�#�O����S�L�7�<��� �r��\����N����Ǉǉ��SAM	�� QG%=�2���>�(��C!;���C�rZ� rC�	T!w�d<�M��l"D�	B�#�1((� �Ga�-<��r^IB��E(Ё��R��p���3�{���d.��!�J�{�S�@U
%.C�� u&@4)�;'���}� hJUu�\������JrJ�а��s4eJ�poW]8�@ѷ6��ND��]z�������o�T��o=�~���>����T�������b_�Uó%*����'��3'�5����^b�;U�g'jO���"y���Ї�yr�]FH��q���*����~��bv�!ϱ]M�,���;��s 1�-�誐����$�Ի��E	�:��O��?�Jk�"�ʾs2���;_�⚢��^��ڴ5z7��]'�QI��)�\Un�b�l���s�X�TS�5�b�^nj&⎁H��Ѣ��hNݯ���ΰ�p�s�Q{(���j�m�jq��x�=zK?��_1'�����P��c]딹���>�GCk�u��4_O3������QI�>��֖�����j����{��(K��h�q�/��.CsH��M]��y�錺.��ǆy��7K�C-�����v&4��jCI�
�;�G�5��x��Cw<4'�¤N��)�|d����yyb�9��=դ�Ӥ��[���_`P���f~I%Ї��w�e��ǫN�'��l��}�X������>��bT�m�`�yfϢ��:�L��pv�׍�ȇ���>>�>�]j��t�5����_V=xI{Q)��us
�&����6�����"��Bb�Y�����]wru��e��\]����jL�A9������S�
r�(U��l��*�	i]�sV�r���@����o�~a���壱"#�>��c���������vY�"�Ҧ��b�9z�.���ݛ#�4`M���5Nj��eݓ���$9�5��3��s5�8�w ��@́e�z�f�����<퀀F	��?��gx�}�%�hi���TB���[�,Ud�cv�#�3u��aw�2큮���d�>�n���gֺZ��"�1�d�Ҩ��=2�|�7��O�WT&��Q���b�*{`�,��H;�{�v.�fA��H=u]����ٖ��g�f���6���J�F�#(ON'��q-T����S�LS�=�ک��b�~����z�c�EC��xm�|r����b�]�oq����v���l�©�3{Lc��Wy��u�42��S���H��ʵ�5}��/�UDG�?�1oa.V�B�����j޴��A��z��O���#�Sc_t&\��)?^,�`m�R����]��^a[�v�ț�x|3���ŝ�SF7�nq��	�,�Jq�P��놱�	>�JF�����b��4��4;��~�3] RY[/C]�4��1|z�2���5�۪��钝JI�;�ՕՐ1t�a%����%�1q�CsPvEѢ�	s��o��ImLc�Ѣ�65��'e��j��5�khѣB�}���EuO<�0%�͐��i�D`���!Ψi����W?4ڇS�r�js��.�(ZK:���m�y���������$3%xy5������>\k�W�lu�b�"G?5sע#�2��.Cw=xc�y�������/&�*z��i�i������E��!�z�>+�?��_.���aKO̯��L�\���?וVk���g(�Y��*��qVmW0����c<�k��x�F�@]P�І���g����B��n%��_V������[>2q�T;J��n�:����q���Z�5���0m�mb�e%���٨�D�bg���^�3\ߪ)��;�����cJ2�����nW�A�%��Y�b�]	��SZ��N�ʖ�t��oHx�����	��}k�����;�J�]㡜�B�;���ڄ���kZ5פ����=��;�k�tdDlap2]��	�X�n�S�j�c�{�2*[3��rψq�Y��	U�hu�if}sB#� 6"T�q�S��0�nA�rW$5����1�;�6>8Bz-�rv.C��6�%�)M�i���L>���m����.���J��[��q^�5���U�ͪlk閽6��$NP]Y��@��0�}����ܾ��O�r�J%S$bm�mU_�j���������r\��~��L�5�ng�nn̺�ZZ�b�z]1-��w{.H�(�T\�4����m;��n!'Nl~��RGu�Ʀ][�����b��c�SL��D���Q��۷ѻ���0 )Z�#tq'l6��ڔ�.L�S4�����Bl� �R&��֑]�8�+���g�ll(�I�ܴ��F65y����
���M�>-ݒ��9C'���oYP�*��02��z���Ǐ�~_W�]]Ԟ��:�Fcз�qMmCF
g�.�� �[go�$&c8Vx%��ࣿW)��r����ك��w���1ا��U/��&��[#'這s��!�����od`�v^Ŷ.s}�":.{]y�Jr�ҩ-ݞJ���Σ���h��ѿ~7��~�����>5�!�M�H�ƾ�8�����.�1*�|
"��_�G6���� ��t���.�aU,fC�C�T㭾�}
"8a�S�����Ԗ�|KЊ��Oa��Ԏ�����{8�x䲞-�v����X��\pC^8T��wM�1�z����J���s�n�`L�����rqZg��o֡�\�.�8fӡ�hk�&Q���<l\?����9�'�>2�Z�d���bk9α֎�����WNU!���D� ����d_�;C!^2����hX���j��ڥDnd>��*��v[��\�m�|�#'Z�t6sں s	��=�k�����De���q�ȣ��kT�	����)�Ց�1�_Цp�-��Wn�8F���^�C%h�2wb�K�i7ך�_A�h��1��(���	�v5-:�N�����n�� �G�ͼ�m!�U�K|���3�Ǳ@�H��S^�r��|�37��ݛ5��`6,w����7���tw-�'�wC��@i��#Z�"˼�t�[QzO	�����:�H��P������{��{�U�4eF��
�fl]�A�t�i���`���|��8z�O�z�;j��^[���Z󧹗^�e.�|M������ֶ�.Y�M��Oޖ`"J�P�,�;"w��G|����{ћ89�����uU��w�S��usl:F%5�p�'�C��c�=VO!�e��`Y��v~�kB�yZI�ߌ�G0���:���W��y��uO���p��/�ST���ھUݚ�������ɶ�ʦ%d�V�S�����F;�X7�$l��=2ǌ��L%d�R�{��J�l����z):���O�H��N#��YcS�>ݡ��?���{�8���V�)w�^����61�$>�,�+^ҋNN��j���7.�_tb�����fM�a{�t`�^Ϡ���k�}2i�J�_�@EE�����]����2pe}$�:,��$9`��z�6�s]��8��kܹV`�J�`t���b��Y;Pͺ(�Puõ>�޵s0Z���ӥ7tf��	��}�N�NS���Y��]D'���0�.��&d=9ȏ�v�~mnœn�u�p���+y���n�gq ~�2#	zL����l���͆�#\UK��rSs&�U�S��8�	�E�����34v��-S�<�w!˖����~�������ζA�/�B@yO��H�p/�	c�c�f��Ӣ]EЪ�ӽ7ήf��I{�FK-��})�5���v#CG�G0�B���Ð��p��2�"s�ҩ����8Ȥ�m0ovl�izY���4�^c��(1U�ø^jt���A��o����u_?2���Q�%��}�ē�a]"�z�a�#(J��%�;�Ѧ0q�������%��&d-���S���^�Z3i_�����?I�OD��v��b�GM��Zdʥ2^=����ͷ�qp7�h�y�A��n����R��F�z��c:��^0���/؎=�C��{h�^�n��0�ƣM��0�wdS�{/�m,l�ߎVQ��b�O�ֽ~`	�~"�u��Uv��p��mz�c2U0�hͻ�6��C�:�fFAO�^�ŷn
k
Jsd��M�_Cs����z����A�ܠ�]9��f�������1����5q�O���[l|19�k���;�����zlt�j������o�>�畇=x4�b��9}�Q~�c&Z�c	��y����Z��*�]0ݠc^��)Ueu*VUСB���v!�[��-�.�����h�j��!<�ٗ���.ʄg>7���J�k��\�E9�)�v�(�&�k���_�"��DXr�-}W<�Q�P�����\�0�L�{�΄C׭E)�m���y��r�aMU��(�莟���gy� �����������'����~���bm\��!��	�=��m?g�m�*�\_nuPv:+�q�~�$�X���!�7�Я��ܳ)�[��:y�tL���O��l�x���-�6[76��`��\�(�F�}w�n(P�)z�:f�N�|�E�Ѻ�����)�Rn͉x�Cwe�)<Sw?aS�n���d�~`2��?&��q��������/�WW�Q��huh:�5�+�jS��.!Ѭ������?��K8�R���{�g�H���<���`�6���y�Y�"��чiO0��dY�� ���~vx&�m-������6��;��Ϻ�a}�.��}N�����b�qT���ި/Adw8�JK	�ֹ}|�0��dg
���ڧέ��֘s��@B�4>�.LƗ<)��l7��VH��^�Z�k�\j�V�z/�Y��ۑ��m����h�,���U*���CW���U�>����z�O�_Ւ�V�=1p�;'@�e��0v9!Em�󔭡̇71���QǕ=[Bn�|��Aԗ��F����zX�e ���32�VmZ]�N[�Y�u���{6[չ%���n�]̒v��If��kY�=�����崲���k�Է�ef+��P�^6J0�YW�[�4Z1���b�����@gj��ʹ�vk�>0RJ������P��n*�"��h�YjyT�Z���<�`d�K�hu�tK>�w��l2"}*p��˾sŴ>�k��|�z[î�����"���)ߞ�bm�	i%)�A������(o�������:�VI�D���t�(s����E���f7v�k�0�T C*�!+�[sՐ��r��y��C1Y��L罆�� �,e�9�S�q�UM]�U6��8�M-HM��Ьx�y:��k#ƅ��ͦ%����Rʈ~iwư�ml�E3��zN
��W�j�SmC�K'��-�D����ࣲ.y�k�Jq���Ь��m��Sס�
�X�}g�"?�*���U{5V���ӑ��p.����1L�;�*��s��ۖ\�*/&!��p͍~�r�&e����VY��f"�5���8�<�@����t9�:aA*���H��Y'_��f���>h�f��|��c��L{��g���1��/f%A���⁊U���͗����T+}m���c3�������u�+�5�&��Ʋ���6k-U�Ȟ����D�!���i�#�U�:��dL:s���;l�QFw4���s�yP�Ԙ�`�3y1N�0o���E�η�[�o4���R��}X2OxJ�UɾW/O"jo-u�Q�ܧR3�3H.�;��6��{��k���T+�X����""1��v_�dK)�T[�8��8����	u��Gs��i.�N#��?E��/����`�㤔9VӪ�kҙ\)�$�o]L��Ϋ-��R�jN1�+�&�@�d�(k������p�saA�i:�.�S(1�
5�*��?�8Ǜ�mO�[<��b�lE��x�4{�/�x������%{�����iV������z]����0ʂʇz�Y��cW�ۡ�sP�N>g��׎t��4���[�H��S|��SV~�}��[i+�����OC��V�LL�n�x�U�(x%�F�y���)�$F���c�j�#]���T��;f�1^l�c�z�d�0�Q���G��6�r��پ%�XEM��=-�����U�Q"�����8J��_����i�X�O��^eT��4�
�]�|�,\����a�M<C��Ϩt[�����v��"�К�uй��D���-�4ۖ[ZY|#���&�3z�P=<ͧ������!N�gń��0���?�����MWx�S���7^�뤒�R� �ߒ�����u^�5$�h��.�=UZ�l�)uľ��/�'�n�_�9���/e�׵�5t~�*	��l�X{y[sK�W i4��9 ;o6�=kj10ިm��%�ctՊ=�(�e��w,�:n~BD�*�vG�bw���-�|0 ��뤚%\�����3��MV�Y6�^I��<�u��NC�H�C�&M�t=n�_��]�@2v�[�����ډwjY4^쎯蓎����6�����8����E�Cϯ!�Ѝ�0r��<�2�����1�^^ގw֯Ot�m�������W屡+�NW@��4��JL��vo��r�d�=�+%�F=�M�%�O�d�B㙣0��ڽ�Ib�(���6��S����罊�\��v!����Ĝ�a ��h�pk���;��A����?l�XF5>��l���WNK!)��nf���㔞<Q�͝�Gl���w�3�i��ϒ��Юwygl��4�dɾ��d+	���t؝.�c���4S�P��wm����sO��,*���m6�7e�#�_�[�t*�^D4.��Ra��y��yf��?yp�m�~"|)��E�_]�<o�p���7��r��ֲ�r뜵Nz��I���0�lc�e����AgH��5Z�	���k�[�]fc٪�fS�Y�ᝈwf����A��j��>�V;�����G����[�:�7ސ��*�O2��V%��h�;�GE�̖��[�~J��٩��s������&qt���[u�B�j��1(fZ�$D�5@��h,Մ�ɵ� ,��`�`��b����	���4܂�4��I��;O����h�����=u�HE�n��Y��N��]�s��LGeФ����ĺCHe�5Ù�{%�b����&q�����n�}�":�{o=�Z�dN�W)N�1�J%3]pfc.㼣U����&�1�l�7WA�}]S�%�EN���Zޭ�����4�VLWQS�;�c ��Dş��7&�T�uN[�f%{3xs����L����1v�k0H*����FN��)Aǩi9ծ����y���k/��R���r�7o��P�c:�鏺�<�9ɲ�gVv�U&a�k,ùQ}w����ܮGe�r-;�o�X��E,�/2.�lEH3Y������\��ָ�Ka��W��r^�ᬨA[�E�����tdj��խb�&W:�w�:�5%����_�[��h!�pD�n���Q-u7jX��9 -�*~F�n�XltX��]�V)c�X15,����-za�\:�+*�,�m��s[�Lu�x&`[�fz~n�����7�e{���3%d���FّENs��6
b�?֊T�>�Kz��e��j	1��S����[Ϝ8�!S6")*5�x*�����;+�����j�+�_7�}N��W2M#�eȵl��7�I��U��\=8G����[uo>|�)s�ebδ���]��\��w�gÄ|hvC:�#�M0�t##�N�vvtp��$@��E �(`���|r��ƚB�3�kW�l�u��2^�B�噮5�p�܂�/c�E�5t�[���\���^�vԤ�_�;��E1%� v٫`f5�l�c�f�[W�@|�4]�@�s'_:���0���^YƏd��`g,�>e<9�V����Vl;��M.�������g@������)�t�ŕfΞ�V�JEvS��nts�����I#�*�[,h���R(�]�n�Xū��qs��_j��0;t�����фm񂲲ŶoKIN9dQ��U��c����t�(/^�̼4;�]FLS�P(yLQy��ˎ��e������7���������z�FG�>t���vF�u��
��R�d>IR������¸�V�@o��0�cP��MF�h�c1";�:�;w���Q�{H�e�wG:��z��YWT/���9īt;Tj��C�բ6�Ȳ�ܶy\ӎ��z����J������N:J���0��v�[��u��Z�� bh���� ^��`�7o���W.�:�s�Ja2��N����E�,��R�t'��c:�WV	�z�֍�ƺ�k�K��۽H�X����"���^�2�u�H�ȪU�T43��q0�POj^qM��W�݃:�ȁo7�^�6���*�_�����4��Vk�.NN�p�{��){I��_�\��*�XB��b������P
ڝ�̮��t�m>M��]9]p3v(�6a�]i��+,4d4g(\�2)r{���2ró��~<?y�AM/P�\����_��*G`��0�������'����H����Wd�̡)��0������|�
OdR�2\��&M(rS$"0����������V���^u�L��!2ZG�$9%9((w!��"�$�
v�Д�#!2(�?@�cԉȥ�
#3�
rD�!+%��L� ����	�rL�}����9(d䏲�#�>�B��M���B��2 �,�h�Z�rG L��\� �_>;�]YF�WQ�B�睓^j�dR�����s/L��c�>#�x��nlG�][��%�k���ê�m\���&~^� Fm�M�be����'�O󥓾�U+���D*Z��t��n��Ʒg��gs�X6LT�|]Ӷ���Ӟ��4�˰4�7%��SBz�},�5�8���К��H��b����7�3�طVS��2 �&m;/+���1���F3HJ����u���:�f_����7}��&���-UN1�ۀgٕ�r��2��P�*�"[(.��y�xiP���סjXv�YG$Fp�0��قO�jB]��U�|,��N���e^�3e�ȝ�U�)�jډv�w�E�ӱONϒ���S�����Q?��ި�Ox�Z5�D<&ƯwBd^ǱE'�W"�*�ւ�2�m)�$I��+��{]�S,��B���h�=ϿP`��jk&���χ���g�wX+y�@���^���סٙClt����C�<0�0�|z�!�VH!�Y��{�̰�hub�=���c�<G'�O�\�J}�H卿I�Ɋ�?6[��5æ\�.C��[ye��
���ӻǯTC���ݮa�帹y��#_[�R��{�*^����U�B[��[�_�gu�]}�DK+����)�yb�9�G0=���ݕ˿yQ���aʹ��x=���x�Tv��N���om;Zhݽk0c���/��{+V
&(�xx^��i����,}�kb�}��v�)��9r4D����#���a��ƺ�S����#�1�� ~�q������~�M"�����^�h\dÃf�X�pQ�e�=�s�N���}vt�9/�Y0�W�E�sf��@�|lDSL�4C�s���}ƅgJm������RXT,P#Y�tE[��{�m	��0l�6$8���39���}Nj��H��-�M��I|���u��h��E�3����PUT�k{hO��7x���y�g�S
��ˡsL��ʹ����WIȯA��[ɯ7�ip�J0Y�>
���~�SC�h��Di_���"F���S������4�zg���f��;ƛ�%I�N�9��xY�Z3HJ�5�huC�Y���l6�Ԙ�1��5�ݳr$F])�
k'����mqy����~.��3$7Y�$��4��i�=t�렇k�{L��<��� uve��3�'߃�(�%�;�_R(l�op���^��A���]Y���ɂ:KI����փ���?W��6;�DX�|sO9��]շ �CSW	��Rk���:�0'�K~$�|g>���֑T3�$x2p�����t7���i������ߞg�`��5"{�F"B�1����E�kw�=3��u�u'��\�Wh��Ϸ����M�`�D���`鯤)��;���^��5�����Ь�*_v�3Z���E�^���i�ݼ���M�Al�N ��V��.�����ue+t�w����-�����Y�/~�GJ�	������,AT�����ר�P�[͓�"w)����i��1d��0���%2�?b�mK2��x�����A([�a���C>?w_�%ydؽ(��hK]��4^쇑�s߃�It�ҩM"��r�1S�2ʯ�U_w�i	4�
�4b2ǝ	�a0�ke��/;�=r�\W�)��b)>5���h+_��n8�X�j�v�h�{8�;f��,��4%�K�X���n2�Jy�7���"��W'�Q͉�5=d9��U=�D��@>����B�X>�^��\)���2F�P!�Vr7��
�Z�1�"�';�jP�P���v3РBƩv���" W�<�]!��xh�Mޗ���D��<�0��C^7t+���p�lKg�
���BT��#*A�����\�~D��d��A�*u�V��ԥ���qЌ���^1�y}�N_U�\��wD	����@V4�����|����dߠ�&˫���r�ܽ�GK#Z��;�="��f���JU׷��-�ﮱdG
'w�1,����W|�lae�%�@�XX�7}�5��s��[ƹf����Xu�������X��a�B���9�0�Vm,\b���h/e�R=�"�����v8��ar�ի�����PK�����$���G��J<���>�������;���������K��UFk��Jx��J���E�P��ҝ�z�Mޤ����_~�F��N�TJ��A�~_��Y9^朼�ƽ�.�˪fB��w@�R��������1�؊�a��\K���:5]W��T��6����}�_��
��W����YJ�g}-{�Z���o�9���Z�����Q� �;�wkf]tEȦ��sJB(`���KWB5�{j��Z��2cJ%�e��M�d��f��P�����~��9�����>U3=3�ɨ�2	�eݕ
�a�	����ބ�&1��;
�m�����S��%�6��OW}+�wO�����	�����h��_�8��*���7�^�Ii�I�^�6[�wkuQ����ɿDvǣFƳy��'�;z�튎f���[�W5�@)G`����-�m4���=<��y�H�TNPۓ�!���;Cc�N��\����u;�2�\�� '*�u+��V�J�\�ǒ��[+��P�]�<ό1����\�&�o�ND���͜I]p�Mፙ���G^�2nU��*�_]7���Zٌn��_2�&
	��$����TҬ�h�!%����J��*ʵ�����a�8��r�_pǗ����a�)A`��6�����ym�.�R��³����?�+�����qW�j�nh}��Ӣ����-qȨ�W_��M��="���=G.S�$d����!zJd" A���+{�ZE��՘��`��4[�:����H	��y��,���3�>9l����"�%�54�Nچ��]4ek2�t�xr���I������4+��N7 b�e�/���Y��c�E�q_0Y���́�wf��a�[���5��4����Ꞽ�Tƃ���g�|��tƼ=w-sB�8/"!?36&p��;FE�А��3[t�qW�����e���X_����Ns��#CHJ�5(�hO^�}4���`D(���-�?
ݱӛʫ��#�/.�ږ�r��NY��%����S��ty�D�y�k08L�����d?�s:֟s?�zj&|���wʡ�gBeA(A��H������3�Fm�O�a���ĳl���h�r�쬈��>eR*�6�
�R�wSl+�,z��!�=��m����XSTf���%�6ʾ�Y;����3?H��P82�|]&L�^����tJkk�˞�(��Y��a�YN��q����;�L����4�v���]��*����'vi�n3��,��^�*�B.��K��ٖc�h��i���o8���������L»a�o,�ʓ��׼���<y)�XzV��h;�1�'i�N蘻IǡP���
���_r�I�h{z���1�߳v������4[z=���3��r���}����i�3pe�>v�ؙ�����}ȡ\=��Y�(r��z��)����/�ީ���d��+���v��9x�����{~�)쨦\��{8
G,m�&s&(s�����8������ौ&��pncjCa|mj���	�M���O��.���j/�K:��~�C߻�A��6,����^�<st8��}Sоt�7�8�C����Q�����'�~�'>��2��LrN��+���ꘂ�4LtT{��M��v�j-���Tw>2�3��M$7.���V���s�U��
����B�Q�u�������jz��|#oo�����;�HO��H��~e��S�Cq�����x���*�;ʋ�����
O�Ƶ�t�M�Yv�ݘ�n���Y�+�1��sF<&�4&�X0�<÷<>#c�9�
%�`|�gDj9܇���tX�*%8��i���H��� 4<�D�C��2��'�`�2��c�����*�1ԡ��<�W�STvvq2����W)w�:�-H�h%hhu(�-�Z/�Q����К練�e�΢�]��K#뵱��L4����@![�e�F�m�l\��ёA�-�P���TF��J����~>�5��t�Q(���q^�����@�Ɇ�������%�`I�����B~H�wg���p�nf�g.];�Ѭ&��^��9��#'*�jvz7��B�Ѳe<Zō��[ȝ�$�h�_u�)�FWLc�w��ގ���JԦE�	�o1�Z��+��˅tMA^=�y��FJ��щ���s���.�����u99�8ñ��{7A�Q����+2�ر�<(-MBy���{ӳ���&b3�\Nr�}�#�9Wt���q����>b�V�7��C_�h%q/�Ljy�n�SWxB��z�g��di6�&2M�lKÚǡ���ȓ�՗��o&u���,������\KGRKc٬Y�z�Ԛ�lն�h�֭�0Sǻ�e�Ӳێ����83_�g��n|�u�b��9?Mq�;���?x�{�Ys?U�ީ�6j�a����'v�����{ʏ������Q��P־��p/E�^����ҥ�'��RE�G{�"���=�l��(^x3 P�_���#{��]�-=���,PJ~��ӝv�O��û2�vҏ^�l)�����\��6���˷غ��J/9�p���E5�N�K�Ġ�r̖��I_f=��?�=��쭡�wvC�v]��ԟ���_+n�6�f���v�o�U�6x�4{��� 6�%��`�S�:��3%JDʃd:�߻��z$�t/M1y(��P��j���٘C�m��
���}8� ]jS �y�P�hG<�o��y�>ɳl���ub�5D���h���C�s�*��g�n�w�k����& ��|[~�X�6��PX�j�k���6)�!�� �ʬ��ڔa�B��[���˖#/A��Jݠi���R��u>|��7U{"7��6,b�����i�]ϳzUxv�|R)E��u<��:Ż�TՆ���=�������Sf2�y\�}@����^+&m[��j�ɉ�b���ښ����}]���#��&}��f�����[�2r�����elNE�M"���2�a��0l�Y�)Ch��zՎ���u��)����^q���)�y>+q�������W���7%����܆��@�d��N��euKmuF$6�C��HR��g<"��tUlWY�4��t�#����/J]��sJ��`�w/A��%��͎��z�+%�Gg��o�7�O����G-w6Vz#��m��U5ȅ~O"�(�f6b��ЖQG�����6<zfxa��ӣ���ut���#Oxwd^���6/����m�)&4[u9�����|=�����(W���:�����?��������"�t>�l�fM}P�J�9��U�r7�/��Ί����r\����2���=�)O�L�/6��-]q|n6*7U�%��WJ;���@X��7���_�X�g9rw�gf�u�'#�������|���t�̫˺]�56v�b�M^��ǖ��]��r��;^l�Q���di�c�+Y��"�i�YX,���>ަ���(���灉Å}"�ˤ:����<5~�]UڱkO}~M4�����6K@s|0ǜe�d���>��B���sλe�w֌M�CB�[~s�>�Z}��$��r�R:L�3�1Y�L ���Jw65�Օmd�k,�5�����0h�]N���r^@^np;gW	�"Ǘ��yO[|��-|h�)���NԧPM�}����7�	��s�N���@�ۭ�6�BC�h�m��ٔ�Tr�n|�lJ��k�2Pu�s}_^��&�ݺ՗x�v�Smq#d��P\ޗV56�}��2�z�m(�Z"/�NowL�η#�j�ٝ���X��(�6yt� ����0'.Z��vc5Ewg^��dG�^j�@��bvq%�3�O4�jo,w�)ϫ�2�uqq���=��>߿Op0e�U���-RP.;u�n�����sRhfe%��������>7�I�v3h���^�WnH�E����D��v�!�-�u�s{�c��r\W�v���w��cr���6L%�љ��e����"�T�8Ӝc.z�q=��>J��Wu�[H޹���n�^���>�Α6��QӼ�J�dYqH�{w��ia<������=�f�_P�*co4���D��=��t#�67����<����WrK��sh��!wF�jnwR�Z+0�z��ebgO���]S���)<���?T�֧+,T�J��w7p�G���W.���i��(w�5��_��BU�]��a+��Q����O2D͗˨ї�V�v����d�z�=�&H���Ҟx(���C��y����U������qsJ��%�eLڹ<�{�, ���%l�e�[�T'3E]���D�P�p���*Va�����v�N¥�t
��2N��^�5�Y��Ofd�na��}unR�p�Cm��u";�xǧ[_ne�&�ϕ8e�tFU��F�fRʑ[��������\t�1�,J����zY4�wj
�YOmsm��ڕ�0j�]1Y[�����a����Ly�㣊8��2��w@�\Nn���T���j"�'Ii.vM��(1����cZLv��YT���� �1m�W��-c`�#�E��:
�J�����A}�;�1�']+^;���Ҧ��j"�h��j�E����4�M�I�ƍ�QRZ.:�&fd�����$����d�\to���\��wW����A:Q.�8$t}�n��R[ w�\3$X�:�Frro:�@�Z�A�Hs�1݉ݱ*�	O�q��c.v=�L(���c&��tLX)���3���%E���˭��hɲ�����ѹH 9Ҙ����	C�NmS�T�Δq�'tPGhu�g.>�y�p�ivh�Z��MVlW�t�,4�`f[B��>�NQ֋��͜1���J�����|#y���M���=@p`�0G6�=G&�NQd�GɺOh³x����Ϟq��S�@�-�O+L�S!�
�%]���R��2�-7�ی�*�]@F0�Τ�<{�v�I�cǩVj"�+y�m��/��t>&�����y����m"_!ғGn.ʺʾAV̛jTw���VHIkB��M;xX\�+y���y��kn���%8j��Ӊ|��owZc.��"O������hت�]L]:�ӳ]�d$%\�g���ѝ�{�:lW��T�AWy�چ���]�ǣ�w��X"'��td�Mkf���&`8���'�Q^�.�	��f�h��M���R�[Zn�M��06P����z.%Ќ����t�,�h�ոE�V�K_-
]��:�[[2k�'v�|�c���O3�Х�vo@\��7�����~;hP�j�!h{Oni�0�%����ж��.��H�y�Q��]���_P�E��|�T�۵�p9hT��V��oh���x��66���l�5�u���ܣmŴ!=�i-H��Dn�5�ٛk%E������:9#ҥ��B�'w�K}Ͳ3v[��A!�m�ni��s��u���*p�ʺ[]���5,�cN��0G}����zŊ�5n�[|��RЬԪ9SR{��*�t��}S��R۝��ۭiN���\�	�[
���t��yʯ��`��[iQ���nLW��v����bܰ�1�-��_5>��c����L������P�9��H�y��}����G>�: ��:%��2r �,�����2��0���<<><Q=��J��@�"�e��<�����������r�B���������Hd4���������}����ې�(B��q��FAF�;{r����"8ti�����y��C��˗S�l)Lf!�g%� ��2
2�Br�>��(��<����HS�<� �d\����y.JlGP�Ð� P1&T�y!�I��J�N�r�ZZWe�(L`9iFCԇP+�d��#JP�!ɤJA�J
G	z��N^I�'Ю�Tvxxg^����{�QQm˹��n�7[K(�ۻ�ft�˧4TZpN��ޘPA��4�bd&ԡuz�t~W� �����
�AK�Z�m��W��-��6<���h9�o���`��I���K�_~��:����ۼ�5�c�syZ���M�`v+<��J}�$�)�	y@��y;�����~ۑ��hv�D�_�k�bӥ��@w�]���A�f��i�����멂.��ĩ<���N����u>{��uM����Iŵ�΋1/��%̚\�U<�Y�´`�ɽm�9��ۜ	k䨴V�P��$��X�ڜ�/�l3�51�<Y�י��3I� �Ý�����0c�v��Õ� ��;G�)��?�c�@w���#�H�6�T4�c���7�U�6�j��nκ���Q��T��F�(߃��g�]y�nB:�E=�M��V���y[��|��!M�F�h+2�[�P[U�޾���T�v߲ҍ���9��U�$������r��F�Rv�����y)��|�Lk�:m- WFwF��UL�.�n)wXk=�Ҧk{�ឫ�0o��aGO���un_v���ݔ��5Ў)�1����S��Ex+�*��R�+�`]$�B��5\���)��#&�YqI9�ޏ���w�)�%�N+�o�=\��:n��h� %dtT�4�[�*�3!��	t�)����κ��R2��g�*Zm*٥x����;!�w��N��wt�U��3�<���֨��֑�q��֢���əV4{cU�n&͵�G[�ә��$gS�qF<� G�)�zWp��s�D	������\��3nM~�g9�*���������LBީ�����\�Ƿ����*��J��ww���g�@�r��򶖹�6F�93q�k����{�@ſ�J{������s_�OS�3�ũ�w�c�ٛz�[u��D���z=�s�~ڬ�+�~2G�$�~��o^�����G�"v0^=d)2WV���z���C�����X���ݛ����1�n9S�V��3EAX+��l�#�C���p���Dr*�a�ّ������u2mT�=�yk�>��_%�7�� q�8��v�FK_<z���U9vq�����cȫ��%[�ԕ@�Η��^�����s�J���K4�B���/�]�N�(����bWA�̎�JiUu
�Tj�WE�/Lj�oj�U仸�ӣX��q�V��I'�	��ɯ3+���Q��M��](ݫK��qb�*ao�H�7ܡ�8�u0�c��	�C�0��@��sA	p�����>$��:~��V쌲������������GiwS/����W�oV��]�ڴrC=�(���@F�㐞_���z��cY��^JJ:��}�sj�Sƞ$aK��RmJԪ/+O���`�xw�,l�ys ��cR�V�ױ��aݷ�J[�H~�Yz��d���Zq��n
F1\��%�����w�6�V۲���\�M�J���wW<%���"��Q�x��)S�=�yח��u�oO1 �P�T��}^B����>��޶�T���͵tp�ϙ��kYy[��@%?6?R�����Ȃ4��{���32K��ɼ�Ͻ�Z��z�hq�U���ݹ>H�-�d�gLA0����N_V�o�s���Z��]7��_�딒��ڑ]���57Q�{�O��_�>k*c��F:�t��+��s�y�Z<�9�]�����Ӱ���[I(R�����.In��,)��D <��]r��)���sb�>��=�f�Lg���)Sd{��yevg���E/k\�R�N��'��](K�ѕ��Z�|U�t�o�z2�"�]&���F9�^�>��9njЅd�]Q�/��`��yӥK��v_w��W��{�P��rvq>�u�Vf���,��9��ڭ�C\t[��_�^_� �L:����]"���m��Bbj�V�Hv�ƽ��Ξ��>ݕ~�d9Fz��q��;���	4�����"��z�h�֝=��w5sG�d�)��}�4O�uC�uТ�:���{�a?I(�v�Q9�Q�#�Wrrm�Č���8���jgW����s�C��VZϚ�<�|�SW5W}��ܗ�F�p�ҧ)v;j+-��n����[�O��#����+y�ҕ��˥�6ե��,�)������x�j؞�ݹ�ր�w��Cj�[r�!��l�}�Z�i� ר���KL��*v�feu�{�ش�JWU��@+��Q�W��C]�ڸ��kDkS�e���k�]�OjN�-Y����z
�	r�clһ�U4�.���n�M|���@�`�\k�[��K'&�X��)�T!�In�c�횙��;�2"k�C��3yL�����J{|�>ݵj^j[N��WWYK�HQ�Z��\x����R��Ҋ�N,����7I�ݹYӒD�kIѦS�PT�<�*��}���	���Փ��~�^�emo����~�*�2����
�d����q�ޚ�M-�^.��q2_3h��!����j��v�n�T	����V�[�#���˸����0����e�����vC8�; .ސ.�*�6Q�y��%�b�ԠF�!�q�U�\r���H#j@CC���7gH��d���ޣ88����=�,��#N�[���Ewj��F֦����j�>y���;+��A�۷p�;L�l�z�8����"փ�t܌��}Ŵqk�&��܇����nf����n,�oiƳ�{w�er�A%�@�:`?il=����-6���U����)7��Q��+ ��K�s���FZpc�Q�Z�Ea���tk9�0ss8s�\�S<s������X��݌�GH/�=Tr��B�&-鲥(�	��[l{���J�f����^}��ƶ���9*SA���0�]������}&J�l�.�٩0m�nu�ԡ�`�0���G36ܭз�8�wJ���ӣ���8�xu7�]2�������ڌ^k��i���0��R��&���}�yX�Ѯ�Y(η�vDds�������`���xJ�QB�*ȯ��Χhާ�}��Y�Lx="��~sd�9x�V�UJ̾�3&����hS+в��e��c��{�݂YI�2�v�w^�?6�C�:�w ���mm�*�+w�PZ+�f-�7g,�ʶ�����ܮ�{�����grg��t%Ԕ�j/�ݪ	^<��,�T�ʁs7M�)X��ׅ�e��-;C88����׎J��-�J�ٮԠ^�4ƈ���|A7q:��{�:M�d����>��2ovG
�rx�D�K�m#�IgP�^m�w�0�_�߄
h3Ky�@�;�j��l�n�kkyWT��/f�T˖Pْ�Π3?�va��"!oz�q��q�i�����3��{J�XI��_�?�����ʢ��L|=��{���2��U���Eb����{�|��7����(�Z��͸J��0ҳ��	��[`�.��$��� �t��]���y��Qa:w�Λ��W��.�NS`�Y#��[�\��}P<�� �$6�w3�>�9Y�{��S���L�p˘%1y�X�19���	�%v.m�!W�7#�p��N%K�Sޫ�qJ_`������S�}�0�
09r�uq��������>��U��<�UT������u{1l�Lp�5���[����3!�|���Ɣ�#"ݛ�M��z��3O>�gp��h��~��!�zu�:��g��C9|�B���V;��u(NE���n(�f��Gz{���b�Z�R������/|�%�ݏF�l(�/���ɴ$��>^Ϗ�����	y�+J��e>��3�,�>k��c�9�^`�%9�wM�k�?�}I����()�璋[N�u���k0��aި͸�+���e珞���U�,���y��
�R���)��:ռ���xfLf���w<������:���^��U���ڃ���'X�Ý��/ݝ�z`�>\��G;�^	c�[��M5ߠ��%_6.�g]��D��a�����d��fo<���"N�z�0�ę��������_�5fQ��~�-w�Dq��KyՃ��-h5��D���N��:�̑x�`��m�LGy������0QȦp0�J#�uʵ���5��d�}�*�<aO��)hYWա�u}��L5�Z��)۔�f��䷰���ޕ+�>s���s
�p���_��
�(	S�yk �n"�+>m�����ܰ�G��[옰�Hg����n�Mc�7���	׾#��恷�}�+�������$m��[d�u���q�~f�z��9�϶��&3z�lV�U��^}F�����w��-��ab���.��n}���~�3s����9H�K�F;E^��(�mn�{�����a�]V�T��Iɺ}��-L���<�n��hd�~�>�ֲ_�O=d�&�ӿ[3�"J/�ѶM7O{Ly�8m�6(�]5|�+6j�OjT�WZ�������g'�u�v'�؍A� ��<0��d�$Ke���n�g���GJ*Q/���C�d�?�xT��}��v���EW�{C� �Y_l��".��&ʬ���y�-�"�Kg�IV!d�i� ���m��ɶ��n���]t.�a��'=9H�T��N_ǿ��4����t{�}b$�o����,�e�O��!h��Uҩ~���TeIݵu&9�n'ה�Ǵ�G�j�ԓC�m�MV4+�-��:�U���\IkR�{�f��g~�M���Y�]\f��,\f��W)�&�sȪ�]؀���z�ZJ�����4\5�� 1U/f�:`UKz��J�[�	�3B��&��=��먩>&������<�n�@eg���\��c�H񚴅�ӌ���ޮ��"�׊WW�^O�����u>��]�ڹ��Ғd�7*�mX�h:��}����9@qI�f�܎V�5m���m�ɸ���о��{�=i�A��E�M�)���P]���݉\J7~���ݓ]�Y휹�S��a���3@�#Gt�ˊ�_�;�O��U���ջBhZ�LL��`[;��va '��W�E����s�joP�0.94֓�-�ʖ2�M��Qy�A�)�1q��ᮈ~�"׼��fj�	�>ÿ.�=�z�T5C�����5���cI��׻n �Ŗ+[�I�YA�t>s.���r��h���S����סA�t8��e���wFNϕ�?~�R�2�PJ��jN�B�L0L�)�/�r�����^�(i�J�v9�΅l�0<���q�s+<,4�B��:�q�e �1nC3xz��\�{g�`tzJ��Z
�*���m3��^�����mb�0����grf&�F�K]���/��b�h���r��F�|��>�<�"ǆ��4���bΓ:k��x�k�jk�|��m`�d�ny��y�Ӎ�68.6�T0qUNn\h�ʒ����	�aa���]:�^�z,�r�<�-��L���StS(���2�Ov��ʮl�6�t����{���'�J�f���.�\�D���Yu�2�%0����i�~���>~��U9l3�>��B��?t��]�8}17��&�rfVvMw�	Kh$�={��#��:|���G�;)I��3~+��뼮��CzP�A?����6�@)b��1T��^�b#SX�Ӵ/<�<>�m�V8�,3�{��Kx$iV�^W6��Yyo/��̷�]j9�O��H�t�H�,��B�v3�gg�k?%�RީQC/&n��UWW���;<1Y�z�����ئn
�ժ/��y# �������" �ܟg;[�2gZ��}�ݶ)������{:�P���sl�
h*e�	<��5���V�ĕX��i��'eq
��ڣ0j���X'!��$�ݬy�݅�s�)86��RȂ�a���|�r�ų-���'7� +��Z64:�K^����;� �m���_\���ξ��r�n�ꜜ|�D�7� w�N.��W:�S��ɡ[ X�i1��i�O%��eqɉ�B�d�+x�%C�x+D�cG����(o,���͌��¸���f���Cqf���Z�J��}�ɧ9�w�t�|v��$�<��XkVT�W"�.��9�pm���R��w�S{Znv�yP�x	dN�1�1�ց�P#ʖ�]�D�D�3�V����̬�t�a�^��Ԗ�����/P\�Q]
�^@�Ṉ��G��Y���Y�d%:�w���ȸ�@Eю:�S�v�PJ�)εY[�u����A�Ʒ��ֲjX��Y'���t���쁋�_�]en)׼���97�t�֤�899��k��m>m��� 5�%IQ5��D�Mn����ap�zr�k-FwD��}%�Ȧn4�q'9�\�JO��sT�JWV(�z�73Az�T��0vJ�� �N�70R�)�f�D]�7��`\�G��>�D����u�ۓ���fI�'˛�}���v�4v�

vcr~{�[��:j��%�k�zC[
�T��9v]dP<�D$�ZNG��gGʒ��ʦwu��)QV�TN�g�K�vP����4�VR����Á���N�tvG�F��R�B�
U��V����x�L���v����D쮱d�DΩ�YQ3�Mp}�"9+q������f��X��~6')V.J}�Z���yR��a���	q�4_T�!��m���`�C�H.�4h��+	b�J
�wD�y��U�s��]��\F���d���Yʲ7��l�b/���yL��X���M5)��c�t�h{��dG�x��1_9i��"��;:̳q
��Y�[ko9J���.�Y�un:Z�[��ufQAԻ�T �$H���5�۝\������g�m�y�^gn�p��L��1Hc��gn���P��xѺġV�Zxl����.l�:P|y:�����@�K*�
���-���X��y�*������鴇�)��E����R&��Ѻ���e�\���H0+����! �-i�u0�ە�qMwr�������Fcz�Uǜ�J= KMk�Z��%w�u��s���mn��!�ή�J�,A�ì5�v���i;������� �ũT���+9��If��ˮ�[�k�3÷�=�H��+N%��+z,�ʌ�)h+��:y��$Vs2����Fo^̻���ccs��؄����M��8el���w
�YeS؉�z���w[�Ĳ����0��6�i�nID:�[r��1� �!�'4+ܡ���-KHw9+�˒=A�+0,��� ��Æ���|x�'��BPJR����R��=' j�#�:===<�:�$�h�\��� �@��h���2�(��ON��OO=��:��L�JP��cH#M:===<c����40�P�rʄ�^�U����s�2L� ���<�{�;��H���W$ؠr@��#	� r rJ�M��Ҟȹ#JdR!Ȭ��"�����\�Z((���K���<��s�3�dU4ą&A�2"���QU!�%�	� (b��c�4<�V�C�IJg0�\���%2�����`za�G<�O����H�+X�:v ��yKx��!0�?&��¥w6��Ţ��V:z��:�9\��v����RT��ݻ�툷� N40�v<8�b���i4e/��iJ�D"�O�i�í�#��9��J'N�K]^��Sioj�zr	n��Vuf���� nrٟ�թ!�^q�n8�|D�V�X��y�J �g�n ��Ɩ���lF�<���UI���u+�<�^�H��Qo��v8��o��z��Z��+!�s�C�W �se��x���]SG���s�v�|!�vכ�fX�� ޿��������ؚ�ZH�5uIl7H����F@�����Űݼw���2�L`Wp��q��r\	l���=<�H�l�z�d2g��1CI��<b�xP��l�.9��Ub-@�JK˩�lL�/�!&êkzT;�}ټ�ڸ�F=y�S[ɠ$A���,v���&s���n�2r6Hۭ�y]g;mZ��bn��l��#o��:��Oq��W[=�iu\�Vl5�eoY���)tq�i�Uj�V��;�5l�k����-|�2�r{�5�\�
��%���\82�/j��DΖ��˹Q��3�������g �;��εHk�w�����*�����Ώ���`mc�>���)�o]m���^���꺝P�jF�r)���`섭���[~���XQ� �ש��wYx�Ǥ5�UM��+�]��W�v	��{����N�'��.��[D�QQq�2�H-�2���_G�Vg���;G�G;�m��*7{���������mr��v��)���� ��!�l�!c����`}�]�v�$�'�K%ufFvB��x.�h��'`��Ue8��41O�
��6����%�Z|�G!�;
�V�; �~�tw2�_@��Sr3�|S�\d8��Uve	w��	��1�)���٨�u��Ж��3=�1@����[b�P�\���rE[�w��$R��y����GC�Gv�q����͇������J�y��E��n��鷓a1�ݽչ��������2}�1�G4`W�W�(4b[�'ja�r6��]���ֈX��aV�}�	��<j{oz��y$�{@��x�=���bz�{�7c)��Iü�%��_���v�%�;��EE9�3Tʊ|�{c}a�p��v��:��Ū�V-J��unF��V�Wm�5�q3]}�&ruk��F�uSDC�0f�f��LuqxZ@������/MCg��|rĜ2^C�0�C6@��6d0R�-A�I�c7���d��ءY��R;��P�Z����*��-�1O�
�\�vvԛ�s�x��"&���˰�3y���f���l�T�^���Ugh��'N�_cmC� ݲ�֣�iL'��՞�k=�߽Rc*�1��絙F#*mm���:m���܀�R��5W��Z��O߿j�=Gt�Z�@��'�[����jw�q���/U�~��Ey�!nϫpй��sa��6���~�_˪ԥB��Wu^����xˤ5�m]GC6��j����­T�%�8��ms��Y%"o
����U�5m&d��m���ˆe�n�rݝ��n�!��4�Q��?IT2�o�&�R9���q�%�^�o5��tw�����	���P�{j8�j�m�H�ia<��ᙲ�K3ղɐD��yѕ������Z�x?go�8�s�|�'_j�Y���.9�Ԏj���v��	��&C�R�k]Ʌ��w����2�w���ָ'���9=ڝ7IZ�3FY�e^"x����=�q&c���x|�ڻ�x�V�����oR�� 6�H��$F���{7}f���Gtçȼ��m�44�^��t�wo&RO�w�� �]V>S,��}�܎���͹Z�<�<�>�����&����|�L`}U);*�pW�>�7�'��8����^ �F@|�)�~�YEk]!�9;���^��>	k�n���n���{�rc���/:vd@7�r`>��������A�W�~�/����wϟ���{�O�����۔��jDfDX��j��_vm��h��h��Y��l6��⚻����Y`���,��}�o3x�IkQ~�Z%ցR8��zfng��+�VG�A�PK� ��j�O���fl\t^�0��E2֒���n�]yy>,D��B�.z��q�RKb�� 7Ly���n뉹���4�}��lաF2�QݝUh+�Y�\�{V4�o=SNdV�EsZ�B������>�X�9L������Ma�V�|�
�1��ĝ�p'8��IE��5zŌ��.�Z��Q�B�
I
ɥ�{���7��k׮�b�8i�n[�4�kMd�R�h��'_u��7�Y�(�u�r�; ZU��7�+6�J�\��4��Խ3)a���US0�b���BJ�ڇ�LGΥYQ}:�ew ���8�]FZ�w4�p��^�ˡ�vlvF�l�j�2�m֫��؎4;�.Jҋ�g���%���nWI����v�Ǘ�n��,��n���؎׵��g�t�����ϔ;��{������ڋ�ٟ�>�$���M��f��ZaF
���Vv�.��8�x�u-	vρK:�"�_Pgh32�"�]�t�S�K���Ύރ�Sg���\��f�����ၷc̰�9۔��]�������0b��\
����$#ܱ�m-r16jP�"vj.���G�n�FݎߟyO�v�uWrYA�k��c�g�8��5\�Wu=h�;t��A�hb�Ƅ�ͥ/�d7v��8�޸���P�r�N\�9��Sl�i�̬�7Xe���pǹ��7eU�ھA{ͯkڞ��F,x����9{҂F�
���mfY��#��H�|��&"y��^d�t�ܥ��Ck+�_Y4M��r�B��6%�����04�Q�-�y)n�/��_�Y��aͫ�|����]p�b�#:��y���Cmn*�q|_g��L�����!��a���1��p�c�GΚ�M��M0���3v��7���dl���PZ��R�:��}����@k爕�����",N]<]hNx��9r|2��(�1#t����٤+J��T�xb�&6*	i�΍!��̾��>lU>�վ�������^�7-�h���*:B�uF������Q�%T'�~n4����E�t��oٶ��������
�.k;��v��;[��c����vL�۾���ِ<ơ�4� tkzLy� X.����s�hg�|�#|�4�TV>z�`b�i��k�5A'��Ƣ)���ߴ��bO����^�#�fo��Ups'|��
k�;�$΃%�X�3w��d
Ӽ`�}��mE��6�)ȕ׏Ԁ�݌��)N64l�V�m:$��۽k�|�ʮ�m��3-�F�I����䀑�̽l�B�i��m�H�c�p��Ye�ݑ�%I�f�n��`L���cc�Y�R�d�ҧl$�*ݳR�׵U�M��e��(�m��m�7��� �����OrO7h��T\����>�,ȍa��V��j�Kx�k+0^�flS��a�-�Z9�8�{��s��|�3��ȥ�u���T��ft�\d\lV�Y�L�g�n�$V�t}hv���̘���f}��52���Xpۛ0w��97�wȬ�
��AY���f��<Fus�ܮ�+�4�_�6��+�Gb9	�s2���z9��m�l޼�޺�@�YC�:�R�dLdi�ᷘb��n�σ$p�P:�m�uv蝓��-LL�n�Gv���h���X���UÝHA�����֭�o��#��(�]�������62�9S�W1��,���љ��۩�mǈ�S|�`^��k���I�ŨSI����&� v���y��u\H<i�S���?��=���G����1�IA�QR��m[��;��(Q�Ֆ4���y�l3缆*����bv��2��~�(oL�,m��e���jo�X�������Y���/������'�J�+n�;آF���K'��K&��/��)�� 	���n���a�j�cZ��*�5^U.����7���<���S���dY5��WX6�:��p��RȇR��2	��s7�Ox�����({�y�l��J�o�}^�/מ���iU�=���9�W��Z�mv�vDC+̼��]bX�͟��m�F����gb�>�n�W��M�b��)]��᛻�cgS�3}Q
��<�s-L\�v�'b�z��;Q^6�UW���<W���n�w��m���Ef��Ȑ2�=C�:�R��}��Q4���,������Y��굟L��#��i�v�ܩw������Z�| ]�̀ɟ�F��k�)>5q�O$
�Q��A�a�$2�v�w+������M�- ��;Wx�GY�}��+dR���ڰ0���xgG���qj�h���t���D�=gj����""�b:<������(��!=ї��	����݆��O���,e���fo).�ns�r���h���cL�m<i"虨}�ކ��a��AS��20H/m*J���D�:ĪϮ���Yb���'=�su���ic+=�ȈF�H�J�l��5�u�}G�o69������� +q�F��E�ӫjVP�T*�e����q�M�m��]I�byՕ�Lʼ����3�<jVB#�b�W3�3{�)yQ���_[�5�"��,��\c�� ��QL
X�<��u��ogC�5���x��bʛ�77\�
{9-u3��*R�9&���b4�yS�v�!�2CY3�Kk�6l�&��Ln5�6�:�l�莦ܸsx��)��\-�hiyC=�S��W/�[+���gݷ�Ծ���Z_�.������m �3�j/yo�kW��ˆ������>kʟ:��**/�i��܂�JU�_Z[��m�ӵ6��e��������; 5TT�>��i,�;�y��Q�&2�Ep�x83y�m�'�
�Z��|/���ᦙ�Khd�[�<�����>�,�GGKg�v�B8Ԥ
Vx❏J���̚50�KΝ�?��Z��69�@������Ucp��n��y�D�H�s�A/ �z�5���K���;J�^���:s(K6c�zcmP��+5��u��Πx3f�gv�/pj�*9�/���G�v��,4��M�,�-��3)���D��;{p1[wE�Z���+U��kӧ��%f�s����1#�X�F���y7�Y�]ٛ�fS�Zim�K��]�9Wf)5��	���8���ζ�!����-,}w�5���Xcnl�5?;��{���%1:�B�o~S������O���`1NO�>���[K_;91a�k�sI��FS�1Βz56Kp@�lh}�"'ө\��{ުЖY���D��툕�B��'���u�ʎ֖�����&~���#lȹP~z$��>;�-S��$S-g��B��`w^g��`a�B1'z�)���S;G��xMa׎�u��e�$#>�c��:C�l3��t}5ʩ��תrf^V�yY����}N�����8��8��*Ryu;�C�C>�y���v[���bLwO`��dP�Vk�я^dč�M%�B��V��]3D�ro�*���I��=�.x�aU�z��
��*v��8�R!(�m��ӌ�جŵ�l`��_u��_Y���lΗ)���ĖU�\@�cTT8���=+r���5<ʡ�� ��!���h7��-oz���H��G����_�ɺK����%�.'��u'�ʝ�geJAà�vő��]�)+#L���3��s�n�̓o�kz56b�-)�{��쭬}v�a���������)��Q[؍&�^��q`<5���pLf�Ns,���R�0_`|���V�U���f�I�J�۬��_]�(lˣ�FL�$��q�!����M����6��Su2�O^�5�;�Lp-�W� �����[��Y�O���j�6�U�CY��57;t�\n�k&1�L�,�^�X��I��ޭZs>�^(�Y��q�}�z���/�f
�]9nf�W�KX��O�fv�
��gp��-�*ˉp�bt_��	O��ٌa��ocN��#��h`�]���j�a����*�[�1�v�C]�iP�o����ҮkD��<����X^Uη�V�Z�=��t���'Y�d_k��v[�:9��J�=#o��]�iтNy�U�Χ!ְU��)�f�1�
0JNɂn8]-f��V��µ�L��ѡZ�)isF`Ok��,FlP��� �*Ԣ�y�d�m�y�I��w͵1����Ƿ+i}���.4{A�Pɡ�c��ŌN�N]Rm;��+o`Br)��/�5��]vI65��'��	Wb�mG��5ԋ�.�q�w}V�Z�vr[�^�Chђ�h��Jģau��J�n���Ϲ�0�c���8�IE����o/�T�b���C�]C�p��}�)�[]�,G�"�j%���v+�`[�w,�bS�WN�e5�ԩQ����5���z�>G�'��.�:�;z��|*�V��,S̓ [w�;�ʛ�Q�F[��X�����q2�=w2G��WL�푥ɳ|��u���]:v���B�T���fY7u 9IW1d�С@���RTc���V���]�S3���\u�9��4Nt�*B�����WqM �./#������v�fK��K3%��(1nV[�G����E���T��� T�+5�Ť�ͳS$���u��%��Ԡ�aQ�-u,�Uh��	�\��o%�r��|e鍭�����s�(�u����o1��n.���S%����ᖋz���`�˗��zL�i��ܷ�nٮ� �U,b{���+����=�*t�ݶoW˃Z\�_`3�֞�1nWpw�XUm�mpz6��T��u5�}�8���p�xd�X�7*����l�mF�⮗�7�x']���9L槜�\@����L^#���(hSm4��%l)�oU�YO�J���ޑ����A)�>�.v��摹
 �flEv�����F�]\݁�Nm�~u��';r�w�Pk;g��q���TwPf� �'ia'��@��XH�W��kc嵜3���^����vtΛ�H$���u{1䔭v��W:N��{�b��>k(�,�̮�ٙ���N_sRl�h�6܆n�W�w���w�ݽ��}���y��0�x:C�P1SEPf/�>�T�.@���`AAAQi�������{#KHS�ٙ����Dr���9d�Fzzzzzx�)T@R�˒P��ӖC��)(�=�"�`�"8i��������d�4F@���cU�<� و����������2$i(�H�2X�(rL����"�!¦���_�	;��(��� y-4e�OQ�9Dđdd��bTT��	�cوs((B�����&<�¤*���
*����0��s��DMD�0�0L��
�����ɕ� (�(�R��[li������� ����2��H�!�"��������z�3}�1Ǻ�\����s�{�DB�x��{y����f%�taǳ��b��Bl��I{�&=��> ��	�r4s��?~fa]�f�jQus?���ڳ�z���*����e����\�M�����"�y�ٌ�u�������g2��z�C�R�)oW�VI�[C���Ʒ\�$�Pqub�AC�u�Wc�QCr@�
���0Kk����<�ԯeu��(���fy�M��X�W)�5���#����m����o۞�Ŕ6�}B�ݘ��7@��k����ȇ]"���jU^�&(�45�/1�P��_y���`�MS��r�4�_���;��_����I��O�5��h=V�5�M�Kލ�ۋݺ�jl�f���hp��P��KZ2��c�ÿ)��_'�3X_�ϯx�_��q�l�M��8�6�#�E���7�zj��Mqܒ�l�Z�^��ǉ�떎�<��#m
��sr]��1��>�九�ȑ�6��9�5X�H����y�Ay�M�� ���/\��v����`-�4.�K��TD�hսO�Y�'׆�q�m��/;�)�tV.c.�k^D��e����8''feb�i�upw)vT^=����:���
"�)bZCg��u������щغ8�g�)�^��������?
��N<�9WF� a��>�Zzŋ�r�{w��3y�G"��8�F��;��`�����$jmL�^k0ʯD�U��ϰ�='��Y�h@�Ux;U��;�=PE����+�[���a��s����jc��v�xn�RkA�;�)iܑo�'��F��a�U��lw���*�vܹG-�5%1�Xҫ�:���c}薢7.=W;��RJ�J�|�c'*BWuVg!V�Le2�]�~��]q�kr\;e�C�R���m��Q҆*٥v�֩���<�Fh�.�{�N���c)Mn1�+r�W��h�g+��Nsݛ��$�gY���-�Ք��^���q�Aϡ�T�K&8.�i�@���y��]���[g�D�mp��{S�?{�w�"��Bi?"�q����ٌht��vyC�����2Z��s�"es�J�wO���:�+O��X�]R���˙�}짤A��=#��N�b\�U�B:�:�:�*���P�d���ʀA+׽����1!WQ���y�VU*4�P�QLw�e��/����S�X�F�u�ov�ۻ:%TX^��b&V�9���>�>t��͹�r�a���Eed�Ȱ�Pqy��|h�GD�8�z�J�ܪ����X�$�������'�N�=�,��/I�NB}3d��LC61Q����]��S�{�BI��k=��Z_L�p�W�݁��>W�Aj)Dm��������f��'����wa�m_U���J?��23���R��5���Ly�˅f�vީ��wN�br�%9�<M�ON5ٺ�:��'�h�@z��|��ȼB�",�������6���Q�k�1-�_�z�A4�G*u>�ms��ڻ�B*b��0�ʅS��Q�|��˘����x1%)���2<S�{M:�6[���]��k�y����&��ݳ=}�^MϡmS�X¦Ei	䔻��_|^�4;��\���R&N���-�'7�R�5=ʞ��l��r
�=D���HĠ��H������w���Q�Ur��>RT�ob8�t��Y�*LאD��p�d���۩0�j@����j酵yQ
Ƃ|t���y�uF��}Os.��<U���/�ԋV�{A��+��g�����K��i՜��IZͨ\�������9R���h�<%���s�Jt�F�:�ec�2��{��{�:�!�����=�S�h᭣t�+�1��S��KT��~:���2����;P�tI||������q�
�T����]$�ܠzꏾFW�|������nӚ����ts�5��֬%�R��!=:�^]>d�1��a��|b�PjN���2�W)�|6_��$���3z���n��۫i,>�i�����ʫ1;����+Tȭ\�eAKt�u9�ѕ�7�������ֆ�
b�E=s�b5(��>�����o��踭-M��s��o_GO��jh��~�m�s�>0c*��;|
MF-�^�gC�E�7����]j�foz����2��d@Y�ކ�gހz��ߌ��u�{�g��>dt·��^[kv'C4�_��߾��!Gع�a�לm�i�-b>J�C��w%�T�!�N��y[�b�c��Vk��e�����g�t�����a�VuWN�Q*}���j��/��%�sk^�T��Z#�T�Шc��r�W3í���{4vr����`H��H��s�5VZF��GGvT�M��Nڛ�zfx�g�]V�]u,�w<�d�-�5˾c<�Ҏ�y�7�A\.H����V�ӗ"�>1�f�w��5���$�^�;��}L��O���5�3���Hc]eR�1���j�a�uV�:m��M��K:�P*�=u]I�5<N$���&eS`���y�}�i�[�k]X��em��J]�L�����n���u��;[���`#"�v�t6������;B̝�*��VeW�Ǐe�(�a���Qkc��F��F��ls��blG�s�Yi�����[U>�y^og���2�D�*�}�纠����;�A�\3
��i)X	���l%��h��JLg����oC6�����+2�C���!� ����:�O��q��j�g�6�+0���r�ة�p	t�!�nCP�Ρ.�D.2.6<+Wy_�z�"��ys�P�������v��N=o�<56N�0��]�r�v�艈߇V0���Q�vH��qr��ҹk���rok�IG)Υ�l&d���F˫go�G&(�m�\oeZZ��]̺ޚ�ҫ��%�ds�Y��*U��n&u�1r�1�"9	ά�j��+��z�x����􎁏�w�2c!�ޱ�~(�؉�gUu�.KV�v�#�q��w�>��M�جB���1y6�3�oZ�՛]>~Z{Uz��ee���4�n��4ˌޓ�FP�%n�}[���!��5�)%��6t�7v��7�G�bX���%OI�;��ΰ��pا�3��bY�O�]�a�����G�	�����$�&�mm�5�Uw���C�{Ϊ2�6���Z>�����qwm3y�W+���T��OW��o������t�C�{��wS�T�l�d=��]6.��P�-6����Lҩ���׶x����޼/CH�J�yv;@F�CY�� �T�=�����@2 ��h���;����ȤrA57C*���DzY�շEP=���۱8NhH�j�Y��+4��ԥj����8ꁉ�|`Ѩ�EI����	��Z�*���8v��"՛}���K,�61V��,��M;�x+�M�W�un.�w�w�c�pQ#�2ޚOB��i���J�h+s5���p�s�9�m�v�aufͽ�A�]NNx2��
*�R���y�zd�AIw���3:��z.��2�����+y�.�s��%#���u�"=h`G u(\�w�Ió.jݨ+$���H?�3:_z7o��u�M[*Xy���#E_�j<�r�ͿO��W�z�S<����t��d�yt��ͨ7q�4�P��Ў�ZqD��
�2�g\�Od�$֣i�m-��ml.v���g�e��y��0��s]ּ��s��H�ƀ H�ȝ�|��B���YX|��l�,�[I��}��'�v����랝f��+�]�7~)<	V� ���H���۫n~�Ym��Xo�"M��CQ�͘�����Q\�>��?K\�;'�ߦ��;�����]���a�6�q��.SV���F��-��q��o4��ٹ��Ɍ�
���#�C���H�g��\+8,_G�V�a����wh��ms�O|}[���N���h�/!�]��?`E�az+�I5��C���pxE�'�m�h�;��2��S��� Z�w_�k �}]_I��yY��Q�(|�r����E-��z��;�˷�vs���:���%�K�R��B��ޓ ������z�9�4�i�q����R]C�{zr�كER6�:u�|�\
�B̬�-\��VT��;v�/^��G�d�9m�_��ަW���j��Bˋ���ĔQHlN�ki��:mԋ��h�Ӻ.��#��ƽ۬�<�[f�v��j����	W9[�x�'۷�����s���}�|c���Gqh} r�u���iA��<��Vħ�gjΜ���y	�Wj�!��>��(�&}�s4��l�.&��gfú�ݛ�k�OU��&�%v���eS@b���k��W�ه�_���`�Gpnõ�U�Kz�*���Gutq��{b�`��p	jΡ>��͚\�[�D�g`�@�	���+�49��}�ŋ��g\d?G�}�j.�~���v /�Po����C�"4�z��
[ӹ��\�ev�pJ��JO(岴�S�q���}��Cv�_s�+z�6*�Uz�d����ʹu�w�TҶ���q�Y�}Y��+����-������y_��������BX���P���`��
ֵ�g���\b�w�s�z��C��{i3"��6�=#9WR���1����y^���Լ4���$��l� �+c66,3rt��#7���չus��`/d�kX�y��:�%��w�IK����.uc��Gv^����i���MM��1]�}�u�/o���N\�{�<����Z�n.�=Pc�3��a�}���]�#��o-mC��l�+s_���k�]G��e��޿�/�x��1=<��sB<�wP7�x�NOS5����}��:q�[��-A)\��*#Co4f��v�8k�f����W�1/�}"&�fv�d��t�>(���tw�];z�ٛ���a�6� `΀��_)N�Oo�-u��^R|��}Y�/��x��~�u"H�{m�4���u��b�C��קL\JB�׶��-�oQ���2H��Up���ī��VL�ջǵ2�����i���/lp���*8������@��W�g
2MYU�̪*����q�z���]5�L��[{I绷1�mD�[�g�wO��.����rR���Y��DҨ���"�B����k7��_0��%�rV.�?:8��s9O���;�a�96Z[��j��3��O.b��Z�:�o�ZJ[yzUIw�Fgb�5�A��p�J'��oD�����-��ٳCEZ�5����x���*k���3��'J��O�=M]������[(H[�7
��K�ͤ�e���X���U7�Y/Ci�.��f�mD���,���F�
܃?>�eK��ie�9Y�]Mޭ���d��P�twPt�x�l,�u��:�:����ԩ_^��g��y�g��Nl���nS��w���6�oLAE;��U%��Cu�Jʚ�ѧ��Y���a��ڗm}'�`O��~�篡x��i��n}�]l0�U��4�(9�J���-s^��vI������$��k����3�{%U�ɺm�B�[އ["�J��13zj[)�q�@p_Lʻ�xw��_�P�3��ᆜ4�Q쾟@J
��Z3�u����&���T�.x���,�>ː��S���x�fbo�wm����LSJQ :}[��I�sn��W{�꧶��Z��f��7��k{������6Ei�{�F� ������*Ѵ71H���s �E	UBP��  A@�0T ��@7{ �P	D�A\ �� %	 ��@ !�E ��@ ! ��@  	T
	P �% ��  $P	D ��@  P�� ���@ $P	P ��@ $@P ��@  JA �� ��@ $PPAHD����	D��� �	+
! ���p��4H$��	�@J��S�G1L� !�Q��ޱ�D����( ���((1�}s��G�~~�/������ُC�(����|>ߣ�d#|?
�돋s�^H El�������<Q_�~�0b����O�S��D<��_2�.Y~� W�n����ӷ�25"
p~�He��{_��U�x�"75�TDDE��fA�E�`Yd�`�bE�!ZA�A�	FFY`X XdX�f���a�bE�A��Q�E�H	IQ����` YXXF`Y	��A�Fd�fDa��h�b� (EB�P��	W%@�@)D`
Q@b (� �D�@" � ���)D�T()@�)""&D"	�
	�d�bE�$�F X`�`��iP(�S��
)�!�hJ @(�y�QO�O���N[G�(�6������n���� QM�� �ս��׍ˁ>V�G`�9#�d3|� QZ��ȟ���a� Q]r E}o�{N�J����XD@{�U���H
���.�����q��/5��W:��G�^�� ��������m� Q^�׸6�]�G�������|㽀�w���P@ƞ�����РR)H �*P�B��PB�* �
� �#J*P@ ����@- 4�@4((�P�@-"�*PM
4"�)H�"4��)@*4"�J 4�P�"��R�B�H� 4�ҫJ��@� % 4 ңH�*�-"�� PJ�"���J�� � 4 �@� 4 ЀRR@(4"Д�P@�H	B 4�� P� R�B�"� ңH-* �-(4 ��P�@-4��#@�* 4 �#@� 4��+B!J� �"4��#B	H�@ 4R�H!J%(4�РP)@�@�H � ������"R�RR�P�@(
�(��R�УJ� �  �#@�-*4*P�BB4
	B�J�(��� RB
4 �(҃J�H
P(P �"*�((��4�� 
4��+@�4�РP%���B�"� �#H�B�J*�"���J*�� ҃IB� ��+B�HP�@��@P�4-444�4!@P��44�)BR�����!KKKCCKM@�!@RД�%+@����-HP�C@R����%4�KKBP4��!CJR�Д�@R�)M	H%*��ЀR�B'��E?��S��шN���{���r{��t?�ZG�06˄ W`��*��~{�}��������>$(�
���0tO� ��xX�v�^���p��(+$�k3y5V�CQ��B ��������1��  ����( ���( ֢�T (�ln�T��T��RB�X�
q�	U*$DT��BJ�H�TF��Ef�R���٭�%�T띕L�$�qͭ6kM�h�����v��,6�m�e����w坵v���M���\B��0q�v���]5��t�wtq�t��k���Gms��I��uu���a�:�RAb��6�Wmth��cjB���`vW5�f�M����X��ͳm���ڻw6j�픰.K��Kf��S;s�]7b�j���n�mi��E	�*��K��m��F��̭�n]�;@��v � �P%6�c` t 	 	 w �t;0v u� f�[��Q;  X � V� u�@2 4l v�: ����K@�:�eTe�I�U��J��k5jj�     "�2J�(�      S�0��I=@ 12i��i��&�&	��0`��E=�5**�@  @   9�&L�0�&&��!�0# � 	RF�M4a&M��ja��Q���y�?W�������c�I���DW��`��3����8�X3 ���܆@3C �k0`���;0�@f�3 ������������a�ŸX�,� ��dX`f�4�3`�<Y��a h,��`�(��~U�/L�?�����P f4~r� ��������_��S�& [���?��?��!c�(b�;zP4]X�a��o�zq�U���0\xZ�tr��ڱ��O�Ө5S�������f|%�Y��Ni³��8��d�3p"�[�[)1�F�'2��J9x��Y�l�d��SC�mm�:L�zoD��NeR��i|F	c,��W���vfݧaʛV)'��G~���,8k��]��	����)U�@��{,\��V^�u�mPvCm���xt��\�y�Z�1�oE@�����7.�+0\6�J�P�/(嚗w@]�Y7�.��J��R�]��$BX��۫ô͛ߵ�ZSV����6s�ʦw6��H��r�*]i���Pǹ
�Ԉ��-Tu��f�"�l�-2��⩁H��������!=�2�m7o^0䱰�wRSq�Sw�jѮH�n�Z����t�� {o@�71�Xc-�&�´a$Q��kq݊P��;�w�LSڐ����<v;BY��L��׈�ѩӒ�CdnhB�d�]�X#�V@�ǂ�1���K`ͷf^n��1�NM߶�3@m4�ô���v��.�'iS8�+lӖo4R�n9��p���U��`B�Kv�)�ctFA[R;+F@]O��E��dÂ��	�X��J���nT2�m��~^���Ul,��r�L �u��le�l��\��A��*�F�R�6;���A�SE�Y��2��Cv^��2���wp^ږ�� �3*-ʍ���w*2�>�;�d�e%+lJ�\WVmK��q��܉"�9@V�z������ӹA�X��t&(���FVA�v��J�P: 5���scN�7��k%��$�u*¬6�ѭ��ݩ��,��Z��[&�У�.��Ԉ��ޫ�G ��!�,]i��n���ŷ�(S��od�@%�G76	��	i
�!	�y��_d��W%�^�QRP���T��F$�3���J7Cw{i[ýw��i탏h�:�o5R��j�1�;u���1��9��Y��h�fV]���܍8܎L'�m�5��^U�
4+�T-cͬe+���բk9"X�lڼ�H�^lw3Pģ,ۖ�Z��X�G��r�t�ӌ�B��Af��ۺRe6U��n@n�7$�ǊZ�/U�6An��pk� ����������˵�=ȣe��k�>�j����ҳpS�wQ�Ԕ�l���he������ViT�6������;(Qt�2�Wo���(�Ń�װV5�R-]#���S��M"ә���S&L{NXu�^����m�ݱ`^ѹ��m��
0�?�+~V��Ѷ�<H �z��Ѕj-��{Q7K�˭�܎�t&X���h�7wyxn��en]�l��ʴZ8-d,,^<�tZwV�3u̦�bk�i�~���YA���y�x�^k[B����U�u��
a����x�i���F��l�Yp(2�l�u��X_��ϖ٨e�J�z
1�X�h�TΜ^�OP�eZ��st���rTE�UY�g(�D��4�C�<�V���>�[Β�|���X(h���]iu�|K�˔%T�#�Ľ��&�?����qĕn�Mzk�F��j���Rx�J��U��«�rU��-��wf��WY����^����&"1͙���.G�×Zt�,]5Dݶصh]��Ǭ�Ԗ\/5+E6��@*kI��2�e�ܶ�60Ya�b�!���7����peZۇDtD�v4�y��l4˻�m�xкP����:k ����[�,G3&23N��s|�$�Bނ�G1��Gg`�ib��`mm���C1�Ňe*�f
d�����L=�B�L�lM)Z��rX ZKu��hs)�
���+�{Zl�s�`�G�n��hm�djAB�X��F��v+]�e(E�u�S2��kin�b���fmQnlAkfV���2�r͵N&f�$t�Z�h�{��f����p�ܲ�$�R��tn�Y��v��eF֝��A��G3��Q�H�w}�q���͋`KT�/p�*��rU�2�������c�W��u����(!�����ХV�Zv�컻-�t���&Q�r��.�e�'B��l���hGn�	�[��Y���֣Uz��n���*۾-�T�c�w3�)1#)+���7*<����T�5V]B�%D1��k�9f����=i��-]���=�	{��݋s@��V ��ۥ�j9����X�I>�S�omj���1۱�3�7���5��L-Pl`��Q�5�[�l�a�Ie��P�����aA��J�f���|���i���H}�j́Kk1�Me]�"'�p��0Ì������
VR�rT�(m�ʹ�^䆑g���da�u2�Yf�4*n�N�D�۱�Ӕhr���
�r��+i����)��ʵR��3 hީwF	�&)d��9������˼�R�5�Ό�+$3t�Zum�֏�ؘ�Yf���5���51 $6�-, �+	�ႉ��ͬ�������7BU%Z��ت���r��(�Y���H��+�T8!c����n�Ue�ۣ{�q]����?��A$~G�~ c�$|%�I �M�|W�[N��XzO�s��'uNٷ�#8�I/�B葊R��'�(.��m�'�wG��h�.zo��)����F�өA��<��j�o��j����+(�u�W>�ʕ��d֌�=��6ڻ��s���V��Jd^�W,������yg�jf��MY�"�1b�{&����C5=}��N��H�e�\���ۻ�a�B�֩1��g*��a�T�ʝd�3'6���s	��<�ޑ	c��h!��1�=�mD�t!PYm��)�((�1��5v��ڈ����t��ط:zp�Z��2v��	�a!�u�"�¥)u�YhGJ{n��� ۲m��ЗEqj��1��q�s)$�`PoGZ�����Z�m^^����5��gs�b�xvV;+*2�]��*��H��Xݸ7�·^�Ҳ���ԙ�ν�&65)k�)>�3�M]1Fo|��ݭs��ӷ�zgn�lt�G�+���RhTfj�9����۩n�Ҥ����������r�N�Gz���z���gK8`���X�z@g�(�"O$���wHr��7|w�25�0b):]\a ��F鷨n]y�Χ��V{4h �+pݪ��b�Z�*Ƿ� ��c��o�ӻm�x-�ժ��Vږ��֩:oe��B��L��V�85۝��V�v���8���QD��b[�	��}�ǦI}a]�wl�t�ǎW]���X�`��Y3�G]R�pS��x{��=�e\���[����s1ٙ6��>�l�%�r�N�˘�<��^�+I=v�;��'F+w��E��tTb��^�Wd��(�(L��oùK�sdwJ�*��PN�7��(bw��'�oN�%�\��J���cM��G�gA t�2t��E,	��B�J�括2�J�:y��h�õ;l�;��8��{\�]qT��YG����k�_J��!n��Mݚ�MAb��U�څ:��u��nЇ����P��ldVl(oa��iމ���;�jeR�xn��������}��v��PCW	WZ�Z�V���{�X*ӝS4�©e��]��|h�y�.��"��2�,��2��yRsۇ�(݌f++�k7�I3r�i!ګ1������j-U�g����1J��Waz��|����Y����m��5��u���۝��{ʳy�P,e�0+@o�`(D��#����6GK����]k�W���X�X�R�3�G}cmDeQsܢ�K�W^�=$�-��z��su
�V�u�\ɕ�r֕W�'	�,�޽��pR=Ͱ���p�t��7hQ�x��!֓%�)}���[m�jYgEXfWMǡ�Y�X���i�Xv��]iyd�e���cU�X�t9m��T�(J�ժ|n�N�t3�y7�B=sv���C&,1�v��j�V���I&�{�nN�-tť��nJ��;���j�[+��m�%a:ղ���U�wz�tu���+tm�O9��p-�;әVJ��j�#jNVp^T�5���1����5��$�G�&�R��C]�1���f�N��2�i��g�]��j�E6]�t������T��t�u��:
�޴����Z��T+��ʋ����b�hh��Y�`�wS(Exh��d�V���.�X�wv'��F�$�[�=KǴ7@�À	F��h��a���ܫB�3n��R���I�̾땺C��
2�"�:�@�Ʈ��wg!���M�^S�4Ū=t3�ٓ#�Ǩ��u��p���"�4'��N�����@�ۼo���p��6Z��k���B��g��"���@뫴]�rԾ�nnu�uYt�je�'�]܊V�F�8.�g��T��Z�Wq�4��!�N�	�(U�9W�)]����Z���[:�r���L�@���B�wqV0u���=��j��8��Ǫevc��D�ٌ��u�x�c�{�**K�t�',�qo:&u���b���5�n�`��h���4j>W����h�f�-;m^�V����Ci��������my�� ]N�o��zb�l^��5�ɱLn�0�����j��iV����$��&���A�m-�[�^'W&t�$YḶ�;noE.�ލ�9F�3Oh�Ν�����a����Ï�o6��Qm������7�j����)L­�S���[�h�ԼR���X��]�I1�Eɜ��4���8X�j���N��
V,�^s��eۋ.e"��۵w�p�IzF9y��jY-_*��]_a5k�ImA/�T{�
z�-]�fg*f��HLqzz�9�.�{	�l����0I�!Gj���%��$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�I%��$���b�y$�JoHTy7��T�$�M��1Ǳ�eg &A6F�Y*P��d�X�d�Fr�ij{�p�&v����qSC�h�����\�ӗ��Wu��	�K:�� �ٵӹ*�z-��K�	[+w����IS�8���zVgj�ݥԮ�\#1�[�AV]��F�>�Vݍ��*ok�[�eMʕ(�����7�:��³.T���α���t�3�^��+gT�La�y��W��k��)[b���0
p5��l��=�"u����~c���o�� ��Ɔ"e�� �fa�f�a������~����>>�Ork�d'�:��.g�;1`��N�K��F���I�ܨ��Nu=o�����eI��Q�x񔍽<�R��p9w����I"]��9��j;����,c걒�9!ႍ Nb�M����x5"�;+.���fSS����mnP[��ޙS%�F�@�všg
.�U���)ۉgmX׳j�F���� ������T��d�aо�M�Q-�n�nR�Զ�RQR��"�9��F�)�ø�y��x�3b�1.��G/�m�:��z�7r�Y���F �������;{���U��\��Y�h^��Ĕ�i��RY�Z��i3�{-e�����!�h���t�hYI��B�x���ǐ�F3v��I-
�0��3w���F���0:uYF�T�Nt:�:���.���ٗʹoU��k9�v�����wr�����[cw��'ji�{ 8^����B���
�^+OWF�{v�ΰ�c�8ᵑ�,�0��{�֔8շѩ�գjQ�����%�R?�\������5ea�Y�F���bm�t�l|��6�#������:ؑT-�Q�IɈ����7�.��wȷx�Y*�8�b��s4��w-�&��cz'ID?�k�eB$2qUn_U�bӯ^u���� �.���n��tƑ�B0�y�@tu#|!�}a��eŦ��pS�
J��˺�������5����i���2R���ݻ �7�&;��iҵ�w)ۙ�'f��ek!α���b�n�ɫw�d�-J��a���R��fuZEaxm%G�[�s�!ζc��7��h{g6Nރ+ɦ]���|��L�05��C�)�WXo��o���|U��SҌ*�<�ٹ���&2��7�/�Qn��XV��k������8�/�q��^n3uf�:r�^S�n�ތ�:qi7�V����N����.��4�{F�hiS�9��ڇVh����jR-��IM��t�&��AXw[f+�(Ju4�컽�Xc��V�㳛g�$��@��x��:&����9��aP'bH�j������K#�!�>V�#T�ʇ:�ַw�R�f0�L����gл��{���X4�Բn�a��1v��@h\�+�˕�{��[�I��z�� %�5q����jX�hR�ꦩ>�����̈́8����Z������J�֢�P�)�̹V;�Ճ��uܬ�=Wr��W4���ib�+��,N�p[���M]����O��.�A��U�tu��v4������5��Vahi�M1j�c���\�

x�N=�/��͔0]`m�mr&��Lf�8n�A|gB2�Hem띕�5XU�OC����m�]�ij�&q2�����}��!ѓ��P(F�X����J�|����=c"rCV9��r���T��VkU+*�9+ �����lMk�hI-�{�ar�����gX�%�qU��*��T�Kp���N�OF�KU���/�:4	�w�pjF�J����Xx�I%g�#;���]��//���ܛ��F���㎰U³����L�����ř�f�/`��%��	07\AA�)X�Y��������,��(�k�߷2+Dt">c���S��հP���$N<��2�s�M�n������y�J�N+�ą�ٸޥ&W��m��c��g��U�R�o��[ڎ֪NYY��e���Viz��s)5B����x�9l�[���wY5t:�vhb��j
�Ӌ��cʆn�Ҩ�kmw,'�&z>Ԯ�zZ��G�K�.�����ݧ�����}��K���i�a�����H���l(4W.�;���̻b䶌<�����b΁��˻�x*����i�M<��J;c6�Zn�,�Ϋ��4uȗ���A����6D�5|��l�n F}�0�v��Vꃍh�kw��Z�ޣ�<;h�T�+�)Fr�.�w.l?r��gT۵����ک
��hL���؉�=F�WP��M(�|!�pcݻ����o-C��;�6"^��D��W��l7sg����,\7^��ʓSAƕ�v/��mJr=ܮn���i`q�Q��'�M�N�Wy�/�;6r�Q��G�t��e��W���V֩�<���s2�i�m*^�.�c�^[wwF�=:���{S�������gvC2E��/g�����qm�:�eX��\��n�q��lqZ�������`"b��[�lPS��r(�+�u��N�~7��:���,�$yl�+�}JJ�h4�͕,�Yi!x~���w]�$G����[�	Y&p��KO����h������V��p�q��HDWn�ux G%����]}Ϯ�]u�z��&��Ce�ј���e'���;���
�l�}*f�c���0nX�Z�oN1�Yv�e4J	ԑ�y��r�c�;4��o����NΥ�U��������X��#헮�m��̶wtμ�O2����ǲi(U���u�`�2��tɎIs��5f��XV��������h�����ҡ�r��m�=��1"��@;ʱعTѯ���]�����K��G��^��2ne�6�9Y�~��` f��A!�?ɀ�	�$A�� Y���G=O��̢�*T��d���^�64K�Uu��X�L�֣Yf�1��,o@&p�QYy�d)ZÄtIҎV�����w�gm*���)Պp����.!�s#���c�rʈd:c��&8�>�&1�����H��J����Ȋy����h	��Љ�6Rn����L�J��Մ�xr�`@s�j�b��{��1l�I$�I$J2t׍98j�ջ1��NdN^h��Z����'gtM�b �,K�IàX�]N� �r@$�LX�2D��	)(.(��*;�A �RLRD��ĒLBP�\� X�C�	� ��H��$�I(4\� �P4�t�DKKX��I�����b! 	bX�Pr��,]ĄQ$$�.�D����!3�XBE��Z]0�D'p���J-�����W}��P��ȝ�����X;�MJ�6��ш.S5|�]����%Y�\u�V������f�w�]E�A�L�r1����o:���2h=R�'vh�*5t��g���s�������Cҁ���MWeOw�kgs[R�^o�aM�Sǔ݂�$�-o1� ��'D{qo�y����bL���ze-VE�Y��y�ag���M����3M�!6�V��V���n�PYw<zJ�]�}��rBAV�A��SN�O8���5�~�gK�5w%��^��l/Y�j=��>��w�Ν��˶�5�R�dDa��SݣL��Ҝb-�vWB\��QS����y������G�^y�o�ܯ)�;�o���,���N:=ғv��B^�v���m��fyfX�Om��|5�<~�Z8���W�i�,>#�\�a7د+U�Iz�)��@�R�$���˧+��(#�X�b��L��G�}
	EK�罏���]t�^U���{oNn��ƶI���^5r��]H����pS�?�9D�/�"�`/U�v3�;�SC5��\�[�Óm���r���8�"��F��t9^���p�F��g����o��7F�8_)!�d�^dޏ>�Ae�*��O���՜WYP+�陎f���+��;?n	��a}-�ڜ�V�tuz����W��R�h�}����[^T(eS�]R�^�Y�!Z���s�4�z�;a�Tx�K*ϯ��#O�ӗ":x��	���8'z��B�P�(�eo{�d��C]����4��r��@�Ir��6�i#�(ֺ�hY�s�2/�:�����Ǡ�;0c�:�gC�H��rkyL��YpJ_-"7[J�w^��I}c�j�_3Hk��O{�u�z�d4h���єZ�J=�Mǭ-m&T~2��D��xh���>A�~a{���D�/�Ͷ��[� �{{w�+8�;�qڬ�I�Z�'t�ｑ����n�r^U^�gR�`6�T��<^<�}���=t��޾ӗU��J�	Z���p3c0��AgE���`l��0��,�{�RT`C��EF�Jp����WڞIK���U��j��g_����	�s�Z�|GI���^a��c�R:��n���6[}�~�R��i�7W�{&�z���EjN����y"���ubצeN�5�5uf����Yhvb���X�G^\�L8�˽��8� ��
:��+( 7�b��䒽���&�o�6y���S�ފwD���zYɒ�:ݼ5�G��@�=���{�}^��54�S{�kЕ�3V�I�M�"�\���'�A����W�A_�Ȩnd�7��b���*)��t2�-��%ӹ���lӿ���IT�*3cO@Mj<,Gd�G2��egc*f�B����(hv2%1��,T��t��C0�]=���˺�~��~<��W3+{#�$�ufi2�u��^-�eL�gEL;;����=��5hgJ=���YO:Dt;nb�|E�`����~�n�JO�)����;���x��:�5{Gk�!�H�>
6��5WV{jr�R'�/�!kVε{�[y������!G3l�������ԩ�d��L�+����y�~��2cL��-g���L���[n<�W��zw���+k=���Z�\�S��׼����W�+�,zfS9ex"���xijy��Ǯ3.�)z��\��Z��������{7��/n�����q�� c��>|i���y �6�^���X�ZL�1f�H�U?��S��x�"TB�o^~�)z�޽-V�hW���Y=}6��tJ��P���:�L�]l��q���f����n��=I}��By���	�(���V�g���x}�$����W��W�E��T`��o��Uk �8��;��sԊ�`'X�L�[��ΰ�_�Ә0.Q?T�v�rO���* �ۡl\���)h�6�|�:�:�tB�!iEj�:6I���R�v����ά*ܢ^�8#�����żڿm�#ʿE�è�`Z�����e��*����^�yb���t_�M�>�ٶ;Hxpi�|�+L��[G!��Cp��)ܑw�����6����P�
�Z��o{D��GKCњ5�I6�����1}�{Cgg'OZ��6��,��*�[��c�Խ��Ñi�_�AEW��Ɵ�<ho��#B&�5����`�a��l�d������\1$ٽ�����}Y"낙g9�\V�c/].\{j��΂�vF_PR_ma��Hqwl��2�l,����t:єee��ҹs �����u[p	�q�G�D@ٕp�% �6�Bo~�YقxW���dom\�"�ZMQ2���C,.��{J����{b�Tt-�- �q�����1�NWXt�)�1��wR�םa�P��NI�Y�*��՛�:]s��ɶ�S�U��QƁ���5h�t�)��R���������Χ��^t��6��]�:J�u��ژZqЄ�{-[�3y�)c��ح��ΈV�j��v�]�����(IXfENk�g�/�YLBg^m�r�@aeYV�����7
z\�ӈg*Ё[a,�gO��:���W�!��� c�ڻ��6]�+��Kxr�\�L[m�[�u����G�b�h�3���>��wY���,�z����P�՚6��X�W�rp%�R5�z�w��ƅ-�TE-�ݴ���w-�� };�:.�-��['I$�I:��vM͈��{1�~��ڨ�����#�w��z��,�D��Aq���I@�Y� A@�$�C[�� �!�2YD���  B �X�:`�X�	$��Ir�I �K C�@���%�,� !� �I"R ���ӱ�1�̈$@t	�)&( Q�Q!ȒH,\��ۮ�vs���q0	!�#�<����� N>7r3�ǵ���G'��~�6�E�W,�o�Ӣ��l��{dN�vW��q���Vs�1Bj��zk�ꆳ�}~Lw���M�&a�*�k��'O���w���_�������
��k��O�������ݽw\ܫ�h��"�9���h� �z~��2?b��$��`��j-�qQ���W�#����PD�����ޞ�+�̼k^��@3�љ�Ĝ1�(͋����K�}�U{M%��.�/,�V;ma���{i0I��<�5��fA쌕��M���h�N��������vtwh�=�k��"��.���9�ƽ^��@���yv��kI�Z���iy���~.,�Vm�l�C����Q݁lr�e���ی+�dV�K�N���I���j��r�I�2�^[yyC��^�'���2������zħ��u�ػ�r�
v��墰�:O�*K���9�&ڥHD�c������1��l���(qH�[��
�J��4ڶ`�%�i�n��,���j���E��ńW����-����R���u�7Kܷ�v�T�ܘ�d���_tGa�&ob��̐gu�r����l�6���7�:�����|����d/�4\ꙛ�䘌v��b�H���_�˛۸A��ռ^�>���s.~���8By��
��c��o�Y�	�Jk�2�OVzV�J�}��@�Sy����=rs�Ei�����re���ֺPnҦP�+����赛��^:.��nzVLY��� �3�^3� �O8d���i�F8Y�1n1#V��������I8�>`�+kV��K��')�@��Lp���'YN�[ggKm���Y�m��fA@�P�me��+Fh��q��Ff��d��Uw
:Vx"���T�O���0�{#�<��tAzz��$8��vf���_�g��ff�S��o8��+k����ds�T~j����g��X�SB���G�^�6�u^�\)����9�P��tf��z�U���&����'�}?���x�:i"E�tR�ԝ�����L��ޯi��!y���:���;��=�r_E9�yO�I�?�����< ����ϊ���c��R̪OM}X:�B2�H:���&��Sw�>�*�u����V�<]BZ߱��(�P�s��g��k��.����+y��1Q���B����y:�:����������.�Е򣝢;�6�d.�3�M����+�Yh
���';��F��~;�z :��Xɯq���E�2~�:&lC�)hѢuC7����`/K�OP��7yy|�l^$tax_�g��71��ۇz���fg�6����ެĢ�yB��d@�ݘ��u�yWSe�>���p�u)���u�fmx�����|�l]���1�S֩Qܜ9�	�� �F�ć.�m�9��2{��	tü��_��v�`��;9��E��OJc�>,8`�nGF�D>��:������ʝW���T�2_C��P�G��}h��օ��u}��tR�N[w^䁽����m	�b�ɷ�)X��;!�_\8aqO�Y��7�٣�J�����enaۭ^A�,�j�m)��8�]��S���Vm{������/�p����w��!<ec�R�cH'?ld�=��e�����P� �K����/�����춦f�<�=��� ]����i��׷�_-.滷)��&Vs�Z��9��O�� ��VLT���鑱�(��A��|(�p:U������kޑ�{9�^���:j5�րW�Gf��*2�ڕ�������_�V'wu��l+��{{T�,�E�4����Bo�*�E�u1�b��{B�<�G��3UѺ`(u��ܼz�>Y���\��U��kh%�ɪ{#e�kQ��)���5�͘\��1���w�-����37|3C����?���Tg�!-���ΥI�{����{اj)
��;W{.C'�O�������׌ׇ�^yVg�lL�$V�qF�nӾ��?��l��Ö�^��}q� ���}�i-��s��zL��#5��쐳C����2�`�o�W/_�\�f����T?s!��[�/��7/���a��+r����'ȭz�L���d��=}+8�)ۙ���J�(�O�ܖ�:F���Uv��LЁ�{zX�\>-l2�������0�^�®����Lh:P�}u��b�F��p�Z�>����LAFS�VY�=�Ad�y!�ybk��Y;���� r�pt�R�R�:=U�]�.��0wo)�H5n�<�Ύ�X�Ӕ��	s�-fMߐe��}b�����볚�Q��ۙ��u�殰�ȭ���S{U��yvj�
����9;h"���nY����D�7~s�]�8��Q6���!�Y��n�Q"����m��r���.��uwB�ʗ���1"';m�F��v�i�6���M�+��8�(G�W�o�W�+n�q�%4�ۀ�A��|��o%JP��t���M�K��)!{������6&�v�@TGL��� FZ�	j�iZ0X�N�x���^}6�#��n򴬻�k6��u��0�[X��$����j^aD�}ev=�Ǯt�I$�I!�<Sd�ul��S��涒;�*/���X�	�!@'RK �ı �	1$$!�ĂX� %�!�bD�� Y`��ȀH	&!$B!$�D2!���$�D�İ%� � $"�$ �a3��&0�	�]݉&
r� �ht��f$�f@FfdCL�	������~�V��v��F��ڼ����W9�P`4����/�S�Bϒ"V��J���&o�z/�f�T��J#�ʾ�^|7�mw<G���v�BC��u�,�µ�m��U�d�p���k��8�j�wuU�&��ƃ7&�����>�3��s�ηx�6�)bs�'W�F��g���[�/�0�m8���,`s<6eR˼��1�r���)�IA�܅��g)�sr�۳�=ge��.�̝��������^��A������Fp�Z��`p*��h}y�GՕ�)�����Ø��zk�=��9Y}���#�V5������pͨM��Du3�o��u�r��GL�b��F6屢�Ot�\w���h�_#�Iv�+xp��u�ߝ^X��2�js*^�O�ά|��6`�"�:��|�`��o`��i$'0�Y����`��2g�P�3߳�T��j��:F�)�V�����%��} �`4�we.�����m�n�f��9)>W�>_g!�˘%��������s��L�\h1�sɀJ��z��۽ٹ%�r!�p.F�v��-@Uf���i�<:J��k!ҧJ����Y���udly�W�v��������'��H:�����0�
�rpgml��9��3B�-�ɺx��Vy�`���N����.����{��q�-��`^�t2��7�oY�������n��II�&�k�O���Xx�tr�۩���Nn��v�9��δT~ؽy�w:ވn�^ީ�����C�����
����ٌU�8�M��QI��/���;9Y��L��Yl�a�T�i���=:,�k���֝,��w8fש׽u��e�V�pq�6��ާ��S<��IF�Ϙ  a=UW��a=ȟd]�Δ��H��r��.�X]"%�ʶ:�=�&��o2_� ����P�W��^�{�#�8Z�Yàú�{0�8������u<8��Swl�R��%xt�'ԯk@��ګZ}˟1����aP��<�u�kh��h]�V%Y���\��_��wf�T��&�T�	�M�4q�OX|�|K��=֎�2�26s�� D?ON)�{���.#^s$�7z��4�8�/J/)E��L��T������h��fvTň���VF7[Lh���F��h��3PiV֗ב�n���ȟ\Zz�V{n��;/'�p�_vl�E�P�l��A|�v]���o'�W&���f9�����5w:R�:7�n`�*�a�r��]�����T�]C�g9�׽�ɋT�U�D���b���φf���`�Y��7=9�W~��J��1��}�nk募���'Q���q���v$��~�����4yYI34o���q�W��f�kh�P����U��ט���jQo�Z�1�pT��%錌C��Zk����g�cɄTﰻ��-��7�7!,�5o'둵S���`����l�����1��B�mgJ�n��3��3�]�k�m��
_g<  �d�uԀ���MɊ�����}�qڣ&����j���Ξ�j.����W��b���'[,z���s�9�_uq<o���90e�X�0Dڽ�]�MF��$�\箣�|2pqU݋w躣�0߳A.��a��f�����y����[��K{|���$)��̇c��*.� �X뺓=�䣱�ʵ�u�!q\�Y��j�cP�ت���ff1;�\�Hɋ�"n-���I�X�'�@���5t�+�ݼ!��Q-,\ޱ���
�\e�y�ڴe����Rm����g�g�ʕQ
�ku�͗\Œ�px_6���P���͎{��+6\{6��Hܻ���1����=T����t����kt�e�tFm�����v��,"���=�hq�����ɋc}��H@�x�Q��h0��s�����~����O������*�؋�Y�~� ���h�����~O��;/l�#)Z��Zs���r��G7���܈�#��u�8Ƴs}���t���a�:ET뤂����#���U�x���[�����.�e��ͨ��1�Ύ��so�.(a�j�l�1��j�C��B���7�^E�Um$�n���7z�3�k�����
7g��N\���A:�	�t<�f��g_.�Zz�� ��^�i��M^�R�����`�׫���o;�[������eL;��o�s��i�uų�&b��g���H?s��������vwD)��V�]�WҜ��0w"6���.�!U������N�:e�S�Z�в�r�D7�q�r����tf�Y#o�Q�̧�J������o3v)ܗ2�N�=�E�̔(`�oE�k²vj�����OY��]�-o��U��/t�B9�q1F�Cb�fˠA~L����y�Vw�uf�� MD�׭ .L��:�Y�rT���'Y/+�+���o-5U&���U�%�n_$�B��.W�p�Z@M�ۼ?�*N&��5ɥ8��y�@S�4��0����t�z�uaea��s4�����Q��V��Uh���M⿖%e�G0T5+vm�u�s&>�I$�I$&)�l����ws���N�ݍD�i�fB @�` 	�� �C,ĲH�p� XȄY���$� �`��`�E��ȰE�r r�`�X"	3"`�"2,�@rHC ���h�P���n*�.woJ��*��w�ٿ� 3�L�+�Ᾱ��s��*�N��9�]�پ��c�|��FBōu��t���z�LޑY�;J��?G��}�����f=��[m-,��(*�J��@����n�1��H�77�Ø��pe:˝��[Wyt=S�g�5�9φm/��^������Y�n �&(m\SaT*lہ|�-��!�4�/�{ȑ�k��=@I�;w��.�{��j��-:�ubl��]�"w�=}�2����5��]$C�`�0�Z����M�w�9�Nj8��R=�}�ZHɽ��
Y��r=+�6���Z��f��,��x��j���k=��['=4!�$�!�F.@�ә�5�.����tʾ���`\��R{&i	��<�����0��=wK$ nX]�
t-}��h�Rt.G���Zj^-z��z�\�м&7�z *Ԍ[��C3��UU_fq7�t��x�z+'U���A�M����qR�Uy�T�G�h���C��	��s�2l$�])(�kF����>�<�J1���{Jj5m��V(HjM��_��b�7<�.H��DH���2i���W�Nx�����Z�m�Q�ϺKS��m�F�߮_</���4*/"��8�72��%����ٛ�f�#�.��u��A�� �xF�Id�H�>����kC�W��~��3�![k��e!ďI��1�O{���*�,���s�b��d��vT����Lj 0w�=F���b���ԿW��d�N�H��w���2(o��ʤޥ���e�)MH�bjU����CO�wF�WW	Z7h惔�oS�J�7��ʳ�>�v�Z?bT���H�yZ扆�K�u��د(��8�"e�u�X��~}U� S���>�^>�ׯv�%������rU���_��^4p}�)�VnΊ��ZTF��S�<�BJ���:��]Ô8zl�m�D���������+�?��J�pC��dn��O�S8i���c�x��w.ަ��)
��R�(SpX̻������1AV�X�z�{ĉ�]�S4\Z�d1�N+�H�����%��ν�5����d��`%]��}$T��C룭wX�i��pcw�㧴��ק���3�<!Y�C�i�u�����g��w�d��T��v8��y�'�S�p-]~ )ە�(훆S0�b�T=��w�A��U�K�2KЈ۱��T@��r��Lk��L�A>Y�Y���A0�Zv�׸ri�z���nQ�c�OKr�<R����s��w!�P����y��]��
�Rw���e?yS�V�{�����w��ll3�KGo���܎�J��E^Rq��'�����: ����lA!��I�yGr�E)�gnlݖ�J�0����9�I\���¼��69�n>ɯ
0V�B�_���ia���nuP��0�y-�+����M��B�[O�)��$��ӹ�
¨6U�\FZiRH�y��O.~�>���g�z3ۂ����h�������Ȋܛ<�ݞ�ד�4��V!�����Z�[�$��Q�9G���D9�m�+�_��xX1x,�*կ<�����o�M���cݬ�?���eĹ�	�>��(���"8R���b.,���u5�ӯ�.q`�G��`{^əS2u��w\�AM�Js*�+8�$X��������]�]Wu��|�����>�'O�l�_�[E_x�g#2gm�n��s�/��b�V�����r�@_���.zT4��qp���c�?��>���ѯW�*� %����t[KN�.��ΛM����ª�XB���b���l@����>{:�'���Y�u��<�K���I��'w���j����-��y��^��T8yM�d��Z��ե��Fʶ�sO}�eՌ��v	������Ο�} �Y�T/�e�ۏu��Ea�h�0mu��L (==��0���__��V���`b{�m����`�&�i�_;��Z�q<������g�o�A��N�������E)�����W�㪚z�����<�`d�wW�����Z�'i,��!*mu���{�kWE����2(�ȍ���OA-C��]�u
���0.[4l���]�3�o����.��$��#L/���mE���ʼ���vS[�CV]��W��P\Nm�ӯ�����X���Χw�!�Y���:8�l�P��>$������<�5�^ �m,�q�ܻ9$���R��b���&'j𒓹ԦQ����l�WDH	Ca��y��c啴�}.�:�#�LPF�[�\v��2�)*+�O�5�)d��S�Ȏ��5bl98Z����+��Љ{0\^�B���٥-�Ѹ�yPR.�C@]܌S]���F��t��������m}ٲ�E٬��Z�s��<�ݘ�4ݘ)î���6:�BQ�>n&�M�7��z�{z2�X�œd2`�B�^��Y�V\�&�́�CZ��X�����U@���qc���иr���.z�::W1e�S�������]�c�ޮ�P��Z�5Y�ol>v�"�};\��RR���w����k����ӯ���Eb�:P>�A�6��4kw�ȵN�u1�Fvt�%��=��$�I$�$�̙����D�v�����r�70�|.�_�3���"�9�f� � 9 $3@ ��DIf!�D Ć�!��` ��h,!�$0�KA`��`�b@�0$0g,� �g,�d@ �bCYf�ţ���\��<+���M��ZN��H��
�쑸�?� ���{!h�)�^ŉ�~ݮ�5�L)L�)Ďn�ZS����)i<�\�~�O�v6==�q5�	M�8�5�b��)53<��v<3swֆ�:
�}*{N:��~�^�T�@�G��0�!�՚g��_/^�8�TR����c7�p��{����U�����?n�,k`��ށ�!턞d`O�s�����Sԫ8��rSv2Gnk�O|;&Q�@�^������,�,m��O7����I��r��T�+� w׷Y~�W��:]Y�EӨ�Q�f�{&u�Ә��m��j2zJ�����##�7�bq^{�^��ܾN��L�3}�b�7�
�aV��dkK�Y�Ds�*��Ӳ�e�*�Q6�"7~��Y6���Hu=v)��٫��U-1j��)̜�]k5�:���9_M(�5V�{���G���=�}Y��B���A}�v:�����[��;{O�:d
�t>�ԇ���.i�*�ޮ���Ea5�.��'_fQ�m�czd���Yi�lv�`	��v�ZS��IoMx&<�G�N�K+>�yc��KV�w*�\(!���-w-�N�_���JȪx9;�MK������4C_	f��A_X�\����J� Jx�{���l���/D`�!�e5�
�7�z�%��lx^�T��#w�|UJ��k�k�:�E�( Ŝ�����OrΠچ�gwL���-����󰾘�:��2]{������4�Ȗ�ML3W��R�fcиbz�ƣ9�g	��,�\3w	��[O7���hJ�w��5}Z%1�5�g�{��=SR��j��;W�a\{�+�ٷ�������Վ�A��H*�����'����nq�VOt�u^�^�Q�b�TO��&�Oy�c��Ǿ���W�0O�����"�z�)|:�i�Vm'hש�k�w���8�~UE������O���u �Lc��s��]�B=;�E�[&�ծV>Y�}lꩆ��ߚ�<Ͳ3��/Um{r����=�]���S��+��"Р%֡��5{Y�Y+�H�����{�YޝE���=�Gߵ�|��K��=i����Z�d�xMG^#cA���'�Mn�K�c�1�it�Aw��M�.��r<��W�����;'���}�T�w	R���p�o~wNl'WU���%���4V���r���%W�e�Hd��yL�Vr�=3��;�Y�^4�(�7�D6��d�p���<�}y��7�Jٱy'���$g̻�h{t�Ej�:�#�L]2���׎�<ĳ��U_���P�����擄8�_-6 7��k�W� ����ۨ��7ń[�Yx�I�<1���5�oZ�وon�]N��6�7��[x�9e�B��^-y*$L9b��\�;qT��N����Ŋ��ǎ���Q��":��z.U�0���ǲaS��H��6�&�����#�"D��h0�r������a0<���}z�*�mޘ�5��7�����f������Q ���ͼ�6,@K��^!]�����6�D�vbT"�=��ݑ|o�V�g2� �j�ѐ�9�Àm ��{�YD̅�J� Q>W�3r'�PwI����4��k���,[!wi�u+RO5��R�]�̮����;�G_2}E�㣹��*�c���n�"�����u"'Y�ǥ^����r�.�uu�����/�;���2��ϣ�xf�<#5R|��5t��e�������!㑪�9�=�4��>������k4=��Ժq�k��8����mqr9�+��2�� [�1�f�ZLr�;Z�u�#�j�P�
z�9�h:�^��c+7�:z�N�]�p�듒�������sM�پ��V�u��4�U�1��:(L	o|}{��=����ofH��Veaq)��L�5y��`]�y��Z�^ɧ�1ſL�6Y��E�G:�yOl��g�~e�|�7�:��[S�kV3+���)�3O��\�6L�,��u���{���IcC�x&���#�e��#va��k�E$�ѭ�\L�����5�ch������P�ew��3�^����'aN!KV�7��ư'[���U�ҷ��`�<�d	Zmet���zh���M#J�����	j�o�9	�Zy�O�f�lrɮHi�]Ư�r�f�έ�!P��cyJ�,�I���R9��=)��]zK޷W0�Y�7+%K�AӬ�������&z`�+CT��N�U�iu)�j�\_q�F�������W�M�Ŋ�\=u���M��dr��hV�-�.3v�y�[��[��ƽ ,uz>�$�u�w��4֎�c�x�5�,�3t�ey���a��K�b��q��5���7JX~����Ac���ޛr�T�J��v���j�S@I51���Zp�2��n�Ƒ �diAգՒ\]=2�e�����$�t۱�l��Ob�I`���;U��u�i�-����;S� (L��Z�WhQ��] m�X;��m����o��wm�'�/B��Q��۷��Rm��W���ݭ�B�!,�vw�P/�hv�rI$�I�I	}3!�r��}���[)���!m[�4fb@E�!�v "���0�1 �	`��9 A�Y���ć �	  �dXC9g,A�XA�$0�XA�9`�D@E�� "����L��$"�9sD"�����s|�l�	��Ql>��tk���?��5ɻۿ�1P�^�{�s�w�ڱ��κ��;��YՙQ���[�*���_lc�^F�����;�pPgc{~ŝ[x}�0��-C�����d�����01�l�<��yh��S����ޜ��*.��ջP<�(k��d?\����A���at�ܵ}~�&d�q�O�9xL����h������/V.F:���=\�����H�N��d�)�Ӌ�H�7��[W~s� �#n;(�ov�U�>��}Jy�Tn��Ä�-;�3��U�w�zwz������k��^�&aD���Rꎨ1|EH��|�*�c��z���,`����#�W�����L����.dqըp�WS�3�XSI�2�Q�2�:��r
����-�3K��0��ctR��T�/2�\؝6��Pl���@�����A�DRU@�Y�&mr�D}4Iwo�cA0��|�o'"X��|A�\��9Q��'��r8F�ph�5��?bqrڻ�`���,�m�^�����0`!����t��èFM���<ܒ��-��{|Fm$W��z���E�vl�O�s��Lt�<�%P�M��}���Zf�������Ϛ���ER�=u�	�x{��:�λ��񺍓��3xp�C�T_A� Ow].]6��3v���#�D�7�U�6�!.�����6���W��90C>�WF�w ��:ʾ=p�*3`����C]w�y���^��޺�㲂U0i�O	��4���=�Dӳ��i�ތ�y��C�/��l��R��qj��*dԦ��A�/E*XcW�v����7����%Z�$g���@AՂ��Nm���^�re�X�N�3ssዶeїВ�[���x�[V����3�'���K
���^^�8P���Kl�j��2컻ۗ�����Jl\)wX7kFt�O����J��x������mZC�t���/�J5��JwgM>��`uu�7AI�nM1�m�o�rMw�CW��\s�,$+�>Tޫ뽅wFa��P\CT�,lZ�׉�[1+#��u�i�Y\�d����5�s��$5}]ٮ��|�U�-�O��f �L����$&��7x	�{�:���[��6U�
�0؟=9�s���{���l���{t�,瘳���.��Ƿ�I��y��gFM�De.>�G8�T���)�ܴ�ez��t��R²��͘�������N8ۜ���k��X�~7���4/u���m�Ǽ��'���,�q��>��B0����l���Rs�D�&k��2�"��]+�4�f#���E<��L{ɣ��G�K�qb|+���j��)�Z�8҆N3�=ݛ2�R.ҋ}�w���O	��[�.�^�'�]
�f���<il���0)��?h��m�c��Tv����!K� ���Ր�"���^z6t���xpS�\wi0_S�k5�[bhǐG�ڻ	�PP�s=�e��5l/q�E�r���OژVgv���	���<R��N`���v�(.��Řsҕ�9�XFHC����C�I�_}H�e����%M��f-�������=h����Ş�tr�>��gk����h��~�
Y-t���d���*ٞ7�sw���e�R�8r8�0,��
����}�V����o�o!/3�ܕ��|�#˂����u�4�y��6�/�6��=�N�y%旞�S�3q�RW7fڒG2��庒���7z�.��">����㽷`�Վ!یu�v��z�����t0R�����)]w^���:���C���y�Cxa��F���)�Aiᅕn��8,z��@w�n�x]=�dd�纸��@�}e�7��Q�B������l��s]|/ׇVB���-|:'��s٢�v�;��
��1ҞH`����!T<�]���[�6B��J+zz䤎�^\"/\�,��@��t,�3����,�;Y��UU�ӧ���yO��Q�}++0����]��{�F�O!���'ȭ.�ֺ��^������s��P��S9>�[�=��hT�-�����/�d�:����q���F�`q�}�����F�eE���V�׷4{�C,���b��d]s���y�@O�ȷ�>�Aד5=�J�:�%�-����� ��l��2�l˾��m[L
'�	Z�����lm<[��GE���
���0�ٟ:@����5�e�w�-������X��Q/iw˃��+��I�5;�����i�j�5DV���jU��ml��Lj�Z�Rr��Nw�;��c�b��Lǃ*�wc���.�v�\gդHN�U՜
�r
��6�W"�m�G7E��ޢ��
�8.PTa��1]�|Ebk)��S���YK��/�=z������Vwp��t8��ځ��.�S���Itݽ�k
�J����H��B�bn]YV.%�ѻv�+�9��W���E+(�ɜԛ[�\v���Eb��]�wh�{.�޺ z�on
�7n;
��d�$cN��2��Y�}�6�qN6}P[BT8��q��$��rX)#��EgM)��.*e`�YE��F6�Ȳ�[h�ȴ�e賷�_5�C91aq\X���+@Tl��y)���p'�[IAk�1!�_m���Y�i�ŏ.�}6�mYY*C����I$�$������r}���s�S��z��3�0�l��aD�\ H%�l�a$0h!�X0��C"�)A�bY��X 9H�g!�� �Ifa@,!�,��,�@ �� İH%�,K1 2H3Y��`�A$0$34�Ȇb�9��rI`�A`� �0��@h,Ȱ���E$�HX��}|-���O������ٙ5N˫<Q�@�&.Г�����7��<@�eF�9��Z�s��L�X=t�3�\�j� �r�j�T�����*�����{pu\sY}<e����������!Z�c�h�Xfֻ��R��Q��f*7�cg�ښ�n]�%�����Τ��-���.��ʅଽ
sU����ʼaL�*E��]<^v(�;#�έ�B�b��l�3>Ec �wmk�����{9�����A`D�E���C[���{���;d�.CUd��kX�a�sa����K�.B%B�{xV���.(�7W���q������$[��3�QC�p��yޢ��.�P�%����"�|��ټ���k�g�KX��B1�8�p��ɰ2o���}�k��s�xH���0����dmo&�5�9G����34��G��/�ʫ��]\��Wo <��0`�n˒����J��A�:�us�C*j�Qٸ"�9�;����x	�%癫�3~)-}+r�i&���C/6�خjo�-gO]E76HH��Ohx���3�g]t�C��ɚk(܂%��RJ����n?�yye::/0�8=9����7¹}qJ��f�L�`�;[�o��MAR���7��b�a.�����Q�}%�}�u?U���=��{�Pw������׽n�������/^�.�o�{�}9:��|7�+��{�c�դE)���E�kO}̋�G�sLY�Q[��Źm��s|��\[��U���HܙEc0h� (sy��*cJ5�p+���[�� ��������pޝԥȕlZ����"#.ΆmvSdʋSwӤ���j�������6�{�},="O?".,�u���1�=׆���c����\f�қg��K� �8�W����m�9k��\n��ҫuo1ĵe���v��۩i�ʧj�d���vj�S>eTU0�7�uJ��#8׻g]�ľÉu��-M�.�ޣp��0kTE���bn����B�^l�YS%��B
��pG|T9�{����z��f��ASXW�(��호c�N�@,oN�_h>K�������qQzNz=f��ac��!�t��4�0�5�&+�+os����g�n�8�p3����Bt�r��A��4S�0?[쏽�:�����n�9͕�����_v^�0��0����N6�-q��\dƎ���V�I����\o�K�z]�_S��ջ�C�J�'Y�P�N��G�P�W6ȳ2��DYnЕ��kQ��{x�,c �ٵ{`�^����2�J3b##f����F���&���.�(b���p2��ɪ�ػ��'�K;��_%�C���"�=���Ck����t�0{�x���Zt�B��[����W��)��0��ԉhv�de�9��ۗҸY�A�ބ�W!�<8��c�$L���r�gEϟ�M%:�#L�r��㶗\̿h�3G��q��0ѸB
>)l��ï�ł׋����Cb��KaDA}xh�l���"�D�HN�v^OJ1V�C��3s ��15W��_��ج�<�Af�@u��r)��݌%'z�q5�y���U��Sޢ��>�&���G�,��9aa��cpu]�l��v("�H#��zи��g��C<�=�Ҩ��#��2�((�;hUz7=踇�u�Ҵ��ƑFqq�6Q�KQD����ÂeA=�'Nj*r�U�l�E��{��`ϖ�#g\g��1�5N!���Ow�8�:�8��Ș���Jw�O�S����%��������T���dW>KK��p���)���n�8�EC�l.D�Af��o�~��^D���E�Ǖ-~BK���{�j���1Tƒ�.�� M���}��3(eq����|j�.9ֹX��{�r3()}�����'�yԑ�><���|!�
h�EZ�ho=����΃�L�6'k$Š���wì�K�Kу`CN#�²i	(��.�>�o#�^���r7#Df!D�t jh����룑�>w��5I���"�6�6҂hTDr�x���q��w�J6h�J@��,��Ny�<F��}y"mw��z�x�M�"Md��{�\u�Y��i��Z�D�Ӧ�R�����&�g�4�������qQ�[~^��7����c��a
�}4`j����Բ���/�S#���.AGVn("�l����Sn4
U/+r�3�fe_CCU���eŭ�vQ�`�ت��߀��1:�g�@�����w(#W8��/���xRF�;�dI!ۊ�P�/d�w�_D?�8e���Z�"�D�:��26�����>���k���V|p�D�HB��I����q�A�Rj-�$;Bh`"�5ӕ���3=2�)9G�Q�p�W8�x���s�Y��!g�u�Z�R2\����n�ȉB��*�|��8A�>�8��#�\��駇n�J�����9�B�[�l�`>!��2"%C�\���!��J���Z�3��5,ܺ�꧿^8{w�s68m�d`}Na&���P��[��uh�G�6�fp`�F��;���U���o9��2U�["���\��7�R�솢F��9!CzgI"\#�bӛ�b��W�-&0U�4�ֽ�UF��z�V�
{\�A�mw6�ŝ4�v�z�4>�2I>��-�@v�ՓPl?j�GNn��d.y�\{]�E�`�/ 䋏��jἻч��[a1"�0i]V L�I�S�B��0�!���:3�(b�D��RT6sZ�㝻|�s��Sd�]M���M�u��ܽ�=����Tc}��6޹A�tu��n�<�q��+�E�6���[�R-UZ�����b���'*��
\�x 9ka���m�3Tj��GJ�g_DG^�r�z0"���Cqv �܅�u8�ˁ�+���h=V4�6�vZ���8�����ȉ��W`��4�(]4�E�`�QA�"2&��[�S�73�Q��-��;��N�Q��<U'Q�#*��w�E���u�]*�����Vּ�vj�$�I'I$%�y'��ً'E��Ë���]US!��H9@��@r�	,fX"#	1, ��X9dY���aD�,K�C��9�,��Ȁ���L Ȁ �����D� s��`K-.��Z
,�K IY��@ra,�L��	���r�4�A!�̖��-�h-'m�/r��VɒU�mk�ꉬۭ�Vf�� �
&{��#��:p��>)Y}ځZ�6�]�r�)��<`���\�r���C��/�y+1�+/�n�ƍ:�4\��z#m	�~2��V�����=hQ� =H#�_\UD�S��1���)x���܆�I�0�-r�0��=�Qs��`�!I�uB��'=�J�=�~��2d�5�L+$ޡgj�c�0�/�-���
��|��US��q�ϐ{sn����8h��$��s�B��-��G�ɉ�}�o��(���P����䜊� ��C������`�W�X<�j��U�Пue����ئ���x[�eL���}�u���Ћ�;�����jM�|�����>G���:G"£p�EjgudW�S�n��2 �6�C�X�4GZ�ƈ�G�!T���|��<�Iψ�X��q����d��=��g�����'�0!���eR� U����]�u��"�))>!��\o-𛴢s3�;�>R�м\���$��/�>��B�v���i:덙#�
଴�8�@��C���g������8�<�4g�8D�Y�	�m�ų�HW/b`�W���{�iI-׵�}�� #Ʋ��u�<`��Y�H�XGLN����4}#rz�S�C1\��a�QɆ�1���<r�<�7��,��H��'fP9��x�Ey7"��\��TF=�u�|�!7E��S.���3�Z�ϡd��F#&��;-�
��Q�<�P�譝�o�dpه��K��Xl�uG��\�����٦i��+R>�ըd�,Ѳ �<����أ�S[�tJ����n�����B,/h����5쓤A���q�VKӉ(��$R*,�>�G��d����L���(�4�4C�ޟ{=9��9jOZo>8p\�+S�4�yAB�#�x��G�)�9��j}��D�6i�d�PP��ǔ(מ}T��J4�n�9�U������r��ѭë�����-�k������j�6�dD.\����V��5f�6rP���e�6j�w^�>6D�Y�i�ƵqR�`�{�C��%Q3�I20f��Ϟq��s�Yd��liZY����>B
��M�Tlm%�MQ�kv��Z�Is2�P��+I6��w/��aĚȂ�C��˼�o �%X�Q�t�$�XI��	в�0z�gz�ք<��x��H!��ii3>6'�k�Gj�u(Rj<�y!:V�9C�y����7Ǐ��
0|B�ܡ��*[��?g��-��!d1Q�&�Y�6Wj�M$���C/`�D���3o�W��_.Y��Wwc�����G��a�	�vsE�����#�'^z��y�'�a�C�-9p��$騔s]���X_#ش��p��D� �睘��R`��RK�zY�q�L��0���>Auљ��,�Бl��>C��l�ˉ���vZ}2�Ѻ��%$�<E>?<F��s��]��d^��T���Άb�$m�:6�7��%�(�s�7hH Qm1�&jn�2�ϯ�����}0�/{�F�h�"K�G�-٪Ֆ���S�2w��ͥGBP3��sbI�W��T���{r'뭹K��ȯ�p4EΕ�p���r�WKoC�&^h/��K�o��ظ��|0�!ڸ���뭝�V�,���8�xb�����i�D�;�������Ŝ���m.\*�rEbe���8O
C]����jSaDO�#.���������t|DZF���r�:�]fe�$�4��8yC^�d8�>�da��>c��#)u,��n�W�PC/<+��C6�x�s��h���rD��Dq'�!��)�;iT�Fi�>��ސ򇋟�Q&�B-���l�d΃3�`���v��u)#�����d������nK5U�|�&�0���&�'�kݚU��Ϯ�P���]�ۘ��%����V28d㿝�c�����"�b�ˇf������P�#�}�
��1>4v��gLQ�OMuv �.��������8|����m���V�@����`���d�Ú�P]��~ʚ���F�D��>2D2{��`�����^ˋ�✠(�2D�x����\Y�1��ۛsiqOy���Bg����%s�>�谌3���&�n8l�4d��$\]��z�cQwB9Q=��{ȣfȃ]�<C���� ��$B���6D�c�=cujn~�� �_��~�v��C���`�e�#D����7:nD�GN��̂=�F��@|��n��P�<\��0�0��f��oڞs{}��nKiFX��'VB�(�1<E������C�k�����V��V^P=һ7�ޣ�Gz\!��x���gM�Y�	�P��P͏M��0� �ߎ�c�i�C5�g��U[��1ޝ�u7���E8��s{�M5������ye΢0����#�<�}ɟ9��`>�X��m��F�x�D���{���vW�v�B��g��Ba�7�X�+���׷�Ρ��)&� ��w[�=���e#�d̚�6�lU:��`�n�Yɗǥ���[����V����Uit���j�y
�fB^6p�^B�p��˼=s+'�˖�A˝��W8�\p�C��:M\�V%��7(K�g�r�yW�T�!��hf=�`걜��I��<D��/y��3"�	��N'y7�&r��MN��.h�qz�_MvQF� ��g)���8E����?���;.^4\�^}!��#e�sOY��"M�8�B�I���;TF0�{���r �$�4z��l���:��~Mf$i.���N8���gy	؉�3a
�~�#j�O�9厉�n���N�e�0T�7mk�.�v�(����v���<C�ǟ�����6�4@�(ˡ�΋#;�����pz%�ϐ�B�N�e�2[�n�콞���BS�6+eHn�qΑ@�(4��ٺ0�XG��ˍ����tbp([����"g�l
0d�f��0��~C�i�!�3O\�8(�<�$A%Q�C�8�ZB�>�utq����W���M��|1
�v���4}h�S��)�w�%ې�<l�Bm(��8@��m�}}�6}�����F���+ɟ*���۾<z��C���-��*�[��l�N�G�NK�3~�C�5�#�L�E���2[���#���ӝu�h�����B:�C:d�؃�L�>N��2�9-u���۵} � wz��t�>�m�[.��=)]tE�-����u;�ՐG)�@�{v6��c�=P�'Tzo�iv�1��YTk3i�r�����Zdb��۸t|wn�ǯJ!<
ti^�\����&�wq_W�i#lz��L���V9Hݺ*�tnG��P̧���}w�֔ģ�k�3�n�S�Q��d�+�C0#B[��6c����8�"�:�_}o����=
��E�L�+ o����e�$w��`�o5,K�E�}��A0^|�;����LR�`�2=�7MO�"�S@�k	�l]�]j�/����Zt�n��p7B����`��\�&_vQ�D\e���᝭����D^9�@�d{��8��g�:���c絷�	CJ֍���s���ŬR�E,8��RI$�I�I\�N�u���2l�ȱ�wf�/C��g ����.X�e(4��A`K�� "Q@���	`"$�	h2X#2�9`� LH�r�9Yː�@LI�N@	� ��8ba2!̔\�	僤	bD�"������$��
PFJ0I "ȂQA.\�.A"!\B9L: )P�&`8h(�A ��`�:���,�s/��0�C��ke��.�̜H*W�O�Ƌ�2^DQFc\a�#��z�{����(�#ƍ��"�.C�)��S//D�4�s�)A�x8�x�.��!�-�&���ۙ�{=�"y�Θ9I�Ԩ��n/`E^���>��͜5���r�s+-2�����ddv�x�!�n:W��4���Ťa�d�9G�;���|AP����,�$��C5
w���^ޓգ�	<Z�?��B�V��'N՛Uzw'e��$�-�sP��4�%�h��"==�pZ������`��v�@�k��z�i��ޤ f]��^)`�H�ʺr��[n�R3��mk��p$c4윳[�{<0�.$��/��z�!P���*����.���9�8���p�i0d��� ^ӳ�t'W���E���Y�w:&�=�x��Y��9�'�=��k$��}e��QGq�ha����*�.p��i(�O�s�;}(��O�NC�dq)0�W\��5�9�S�7�^���9s��y3�T{_���u���i�}n/�>.2Df-6=o�{�|↑�!���D��!��BuY�]�ȝ�t%�٣�G!QN'W��Ƶx���&5%�|���'1��:������g�f��jt�YWI�kB��ﬣ�f	b��͒5�7����U��[ǧP�����A&[�A�׳Ų�:C�j��߽w9{�Ӯ:�{�-E!�%Ы��8��N��'��q�����1&��fUϖ�A��l?C�Z㎟C�'aD�����Wv��,"aQ'M$ϵÑd{&u�v4�4C��
�B��W-.[Ұ�K)��aR�0�`�1
NF����������և҂����TG.t�K�ĸ��7���/��h�Ow>� P��N&F��.�P�&���"� ��g[�Z���^M]pp]��fr�%~W2�܎��3@�u��I���c;<��g����v�.<�r�'-´i=5-��}���&P��J�q�&�>ד7���]z�<}a$����f��e��r�V3����d�Ԇ�.�џ���W��8 �-�:W��B�!Ȣ�#Gwc���3�!e�9�BA��:���;H^��V�3���Y����	0F�:nQR�:.\\?�x���\BÉY^�ރs�n�u-ܺ:�R�%��ln�5� �a��p��F2D'K�(C㊥�zL�k���Ng�L�f�M'��e�E��BSn<���g+�������x��SR��:	�3.�s:��m�ר��ш���xO�@��Ӆ��	��8���2:��N�=0���+�c�0���)��+�����xΩ����yi���&��X4nԖ�O#+7�#yAr!����#1Y�TT�[��#'Hr;B�m�DE'.15�,�#}�}��"�����)�%�!�O��{�S�^r�C�Is�#H�L!̓��O�/m�5�k�����M���4@ޛc�`�M�=��M���vU/hY�&���^~�S�����s}����A�78�K�X��)�Ft�K�7�K�8�Gbc(�7�s�7ԲW.[���ڼ<oQ'��[��n(6��ɑ��@�E������#E���}0EӸ�TeI�G]A�O�.����1"\��FXW��ۃ�s4�Ɯ��z��F�g8S�Hy�o�nu�c�(�y�IӇI�ըYEBn�{��ٶx�$9�Dj������ј�JN����>-���sp�Z��y5j�������p�#��'_K��N�I^�z���\s��Q(RZl�.l�B{9`�z}Y�<!���;F��I�+#H�L�������T�WO�Q;��o*X�lj�����n
0�1�swJ��b�1K��9f����+U��.��ٻ��<|F�}�N�e�As��NG���m�h��u�� ��\rп ���FH�f��C̶�wzB���׈�B�Ì�mk|��#�H�p�*#�HP����:&�b��B���B&Hr%&)A�TwSj�����Z ��c���3�X@�,��8�ѩY�:�|p�:|h�W�S+́�P@�I����[���PG�3��^��u!�+\HyYQ�/a��AC�m!R��\d�&�t+�^�E{<a׏�!0��"��i�gBC+2�ymTw�`�+��M�]���#>8��� 9�um���[��bO������h>B���r��KR��v��5��p�㇈�VF#�Q�p�FQ펙��ߟ�7�	1�K�d(S�
t%���$����>����d�0�n"d&�"�RdeVP�vE���i�A�%��XG��#e�_ny�;.�Q`�eI�D�C%q��{�6�%���vE�F��܅������)�:���&f��!�`�E*HiƑU�qo���W�t��d��EM�Q� �"���1�P��،��3P{Xc�B�h��j��#C�r�q��9��On����7uf�Y�ř@k�;.�lT:u8$4PZ�f���@�d�C�xo��O���:r��G!�����ǈ�ohQ[�\�|��!��a��x먐�����>2l�5ˈ�R�Fr���k[�#a-�$9|^��S�i�Ϥ>���2Wj'�t��"a7t��֚XzQ"����.-a�ME�
���W%v��6b�Z^���p�"ŅF̜�l�'��I�:�����t JhdKv>���I�3� ��@�Ŭ���%9�<l;�ןҟٸ-0D�g�!M�/G��~�{�]��Kk�H*���Ȗ�ٲ�h��s�~/>˜���WR�G�7��Lơ��iQDM�|��w}x���U.#��&ZdnEd�������y���l���:C��CA�2Si�'Ar���N������GiI(FۄD�a�}���@�Q���f!Qo�2��6bu����O��p��y���/s�Ӝ�7B�_;��r�rF˖�3-���zޑ}�t����W��2��w���A�,�����E��=����8�����X��`����줅2�����zz3iC=.0��Ix�'��dQ_��q5}�l�ȭS(A�D��M`)��6C��{%S���>8d*�韫���ѽ���蝊w��Vvƻ<'��3�ոr�)��BvN��2�;��!ڲڲ��L�{�񛵽
A�5��Ѽ�/��+S8�R��|!W>
�,�@�7q,W�/'F�e�s��R4��N�5���uv�qcR�F�ʵ&i�`���܅��2fv;��n��އ�V����'�!������޾�.1"K���őR� -�����YF�:��j���6z�q��6�:���B�rʖ�[�c�|0����n��U�}�%�ͺ�pۮy�8�L����x�-(V��n���f��u�܁f	�j
ov�[e)}����2�B_tr��1������QR��1鏀����ӹ��5Һ�i@]Ʌve�z��6��oWb- 6�^�{�+[�WP2�Ы�c\���!�8[�r��Җ8�8�pS�J&GAub�S:�	��l2�Aw;v0]�YSu�]ZȮT[�p���έu�BdU{v��3*�V'P���^
������2�=�E]�4��{^�\�)�^z57V�$�I$�D�铢�i̓�L{f6T�������ub��˺�N�KqFA��QJ!I�$��%�,K"�0@�RBI 	9`�H�Qi�vX'9%�N�L(�Rwt��	�1"RA`H%�b�e	p!"A���a, ��!ˡ&bP�X� I09@�$�B.�#�HK�	(�|n�����x�����v�4Υ�7$�9$է#���f����𷂗�c��.���Z���ћQFό6�߬�ZbU��~w��˷u+�z��sECH��dasD��R���f49Dwy�Wu�)9st��L���VX��z���4y/H,Nr�K�;;�8ErU~�{��ώ�
���>9h]�@���'�%�";��e�������"=��V�F�."x���^U���ӡDx�MEyQ<�E8�\`��I쉧��.Dt�d�%�(;�����t/=����>j�q�ϱ
�v�,.A6Q��3�t�63�ߎܛ,���&��rXi���5Fhdv�!���񂒔�K��J���if`�̊���
��jrT�୞�w�( F�κ�툗��W	C_H:�j�ڇ:q!�ƪ1dn�P"iV�R���V��^A
ۡ�Q�Hh��&�B!A{S�@�Ӈm�Wo�<|Z�EE�� �)>�+��*��x!�w�hٓt�
0x�K��w�Ρ�>��O8�H�"h�&T)�3�>L�g>?�7�>2`��NDU�A.7Zr�F���XÞC�[��D;I�o&�H����sc{��E�r=\:b���0����8�scH�G��,�;d֏C�75��6.�Z��0,X+xa](��Y�ѽ:X�3c\RH�ĝ&s���;r���S�:ظp�pȝ#��VOX�3r9�'�$��y���57¼R!vԱ�{!��62�>���K�\8���{���ڭ��-˻�|f���V����2��pI["����m��C8h�L䛣I�����9�k��:6{�|}Ow՛����=iVes�A�j��d����S �O�,;�o�vrҕ���
3����]��]���+E���(�TQ�}���=4P�����J�g��T%z^��oj�wW�W{E�M�/
pj�b���N��WՓF:�SJЭ�[�x���4�O�d�0-�q	a�J/un5���������.gY��pj���"c�M��/�uN�����S܌��G\ɒIu���e@PS��c��}2�J�5ߖ���K����r�^*+�]}]L�!ީ����!���@���y(��E�`�ɮ��ӣ�zVc(X��Z�x�u~r������7�(��o��g��HU�su=f��h���(�=:�!�σʚɟ���o)��n9��on�0���@I�ѭv�M]B>㈐�������8)��[c��o}��v�rb�w=̃ܫj���6=v靬�JЫ���`{s�%r�صɘ��ɝ��뗙��l��.�&(Dԫ�=��^CQ��ʩ�}�51��4b�;�1.�7$;���M�p� �h5;<d��Q}]���E3���21?k�ӥ=�%[�u���|�7�OS2�Y��]��|uSN�����"�83<굟nb�ww,d����s�l��M�W1�����v����Ȩ���l��E��w�p��kW�+A��*��̮���h8�T�rQb̎f)�	u7�wt�5n�R��4� o��콥��0B�E�Vțf+,r7t,�eƷR�u�I�����A��Zw�$�R#S���5͎l��z0|���YE�(���os��b`���W7b�3���_�4�n^��1��GzJ#�Ƀ!�ϩ���s:GR�v���q��5ʯ�.�}�������%����18!�c��@�r��|�kl�آSYuaTCy!�76����.$y1%��t"��2�̾���d}IG�K��G�����緓�:�sb��Pn�l��F�j�j�uz�No���7j��J�.���3�v�P��8m~�W}����N�f-󇳇H�,F���̙<O~��>o.�^�
����q)���,�V@���d���	����ѓ�E�X/�l�k2��fӴ��U���=cS��#a+�л�|f�\�*�xW��,��8]k���Ӝ24����7���yb���,��եݍ1C�m?D��|+� �]�/���5tвvL��G��>�K�۞����S�i����ohpQy�
0y���N���u��}0p��V�#���;{9r��n�]���;yᓠ��Og�`.�%dκ��{'OU��0��sl���y�Y�X�N�M%�ޙ�^nj� ك;+�&��c�	¹�����qIC��z�⥊ǃ���b�z'Sn-�k㈟�M�geN��b�9��~2'o{¹��Z77G�Fy���V��Y����y|O�v@"���1a{P�:����&;w�V�ؗ.�*@07Uom$uGn�b4"�����������I��]�7fT����x���? ?����AI$�I?��@0�3��� `0f���@k0 3a�@A4=�Y��&X� M��>��4�ł���!zû2* @� j!�` C ��f�������|&o��<���5��������r� ��~�C�-e���~f~Q��͆x�@v�������H8�!��?ګ�8� ��*�_͐b�ǹ��o�"Fx 3a��=�����w��A��Xo� `�0�0@� 0f���}��K���7��1�� >��7�h��?�����?����?!#�!� ����� f�����wo�X�@��8�#8�����)�hd+�N��� Hc�?�R� ��/���������?~Q�8����� ����v` f��-���������Y�f`Ā���}�fff�K�fA�>J�����%��	��?�� 3a� �A!}���7�_A���C��40_` ���6� }c���4��b7�Ä?!��d?���wx��C���Y0`0f� ��b���`>����>�Ň���(@C����|Ӂ�!a��~��}߈������̈́�?�}����|��3�W����>��3 0fS����A�X��3�	���a���r��0f��?` f��@��f#A��,?�L��F���f���3��ߠ����f�3
���H�n����1�0�63`��BZ� �h�@����8)�E�b��a,��مPC�0 9 �,	������ f�Y���A����0F` f�������fb>���S0�A�������� �pc���|�8f��c�@������7������,?���� ��>�?��@���3�~-�|��0 ��� ��~���1�����3��$
���8�a� ��h�������a��6fq� ~��T��"���a�?;3�և�� O���<@�_�a�����a?����1��7���?/��Y��3
����@O����.>K�����������x��|!u/��!�������� �3a���0�����fC�7������X�f����x[��M�}ɚ��	��X	������"�|� ��[� �� {������"�(Hk0m 