BZh91AY&SY�";��>_�`pc���#� ����b�  �    (                                67� �p z ( 
P  
         @P�    �        gǕP����@�P��*�
��U"�@�J����TH�	*QQ
����)JQTB���� ΕUQ"*T��
 �F�@�Z������R���2(e��Z�U+XM�DM��wB��ހ  �  ���.� M� c� ���
d �n���yI� �@��� �7X {� � �|� }�))T
P!AT$;��)W�;� q�@{�籽� ^�Ϣ�W���:�� �0c�p� ^�; �<$U� �� A�    o� � }}� ۊR�� �9 .�4� hww n�"� �Ðu�� �� �( (��� �T�JR�E*���!� 2�� t2 \��	pz(ݞ� ��C�i�t)�� 9c�
V����  �{� � � t���6;��R��z��8z�c��4�.�����a������P�#�7�u�P��(sg� nh   '�  ���I �%R�@�EA����vz����7gOZR\yJ+ :���ȣNl �^����@1�J�����0�n`� �  � X� 4>�u(Q�Ǆ�� �y:����oX*# 4������ݎ@;��%;��yؠ@ P �O�y��HU%UIR��"��*^ H� ݃�2�.`{ǀS�	@9@�� ^�
�^�P��A��� � �K� n�K�g��ê�݀�9)Wr 8t� �P�A��    QE��
R�0�0 &#M0i�O�d��*       "~MT�S��Oe@h�h 1  �*��)P      z�"T� 2h     �=F��`�Sɤڙ �#&&��Ow����������
����ptL���玛�`�
+}��(��"���AE��� El��^�8AE`~��I'�AW��E��PDW_u��>�(���1��0�/ɀ�@
`�ɀ���(�`т�0_��  6��l ��Pv� �@l �U�@6�Qv�v�Ev� �A]��P�]�TlD � 6��Qll  �U� ]� ��ClWlWlP�U6�U6�Qv��S��� S  6��P]�l@P܄A�Ev�`"&�"&أ� 鈻`.�#�튛b�0v�M�Sl�6�^X��킛b�
��أ�(튚u����< ��m@��,H2Y#��?<�^�\ool�!M��ܮWvlt�����i�|7�g%Щ����gn]�����G�N�^�����=��7�X�ѫ:�kZi驸���_NXw�ژ���:1mȈ����br�	Cͽ�)���h�ʤ8�wu��N�1�@v���Ad��L-v�������d�睉�B�ˢ#�B��:p֩�d�g+�T�N��kbk�8%�3T�D���7k��ya�j�f�)�Nn�"77r�]���������N$�5ҮpV�l��R��Z6��]�/d��D|92�k�00j���rr9 R(;7t�,�N�c��Sb�exww ;ƭor��u��p�r ���W-�d���b>_v���^�~#Sg-X��:��n�v�������t�0*��PEb�ו���aht���ٲ�,fr�q�4,Qݍh�e삱�e��C7aX9��-O�}6A݅f�2�*2W��m�Mp#f�;`v��y�t�y��b�p��&���1�mW�q[7z�z�V�Np;�QɳR{*�[K=Ŕ5H"x�������(+���#�����"�u�e�:s���;��Z��Ç3�8)#{��8���Vwa���`|6b�=c#9�-9�Wvjy2v`����op]���c��dd:���-�{�#��qxQX���3�/,�Gwg>����^����;D{}t�Վ����y�f�ӿnu�/c�9[Ͷ^K2�51.w6{	�p�׈���i���x �&�ŅR���R��^�R��\X8)fSi��g5A�5�Ӻfn޼x�gB4�;��_x���� �^�Mz��$�2}Lm�"����=�r���=���{C�oj	 �)�2���ۀQV%��Yt�����wK��q�D'��2q�m&�T �h̠�)�iS�[��W�)���ܻ�nZG�w��nx�~K$Hyhy�W�8d�����G���N�-c#���`'�a��1���<C�GC&Ke�\�,XV�t�\�a--}>�현X��p�H��:��&��T�Gdw;84H����h��A&�t�&$��/^V>��ߵ��UH��ׁ|l��D�"�s	�緛�9���Rr��]9n��]=�/v�R-$ջͱj�7D���2+9�q��Ր�x��ϒ6t����������^F�>,����L�@���rY����:8Xh(���#yj-[�7/_�9�n�����ƹ���V�CV���y���P����q-6t��X76������u��oUǼ�s[tfl�	�v�V,%���vs��5f�oi$�� {�b�@���:l]��|q�*k����.3�vs9#�	�TQ�[����#xс]�]ݏF��d`��V���k/qMV�"��E��nRZ�7ՠJ��=��l�f�vn�-��6KfL���x��gLق�;��W�l�mͱ�����Y��n���S�Ċ�= ����[���ڷ��o{nˉ�{�q�y<EZ��o�C��9s9��Y�52w�� k�=WHBP}&X�qa�';J��f����t��Fl�'2���c��`;��嬅����<Y�â��B��]͵�w��ܶ/�	����8�a�s��2Q7�P�q+V�����';Bƻx�����&oLY(�4B�K\軸;fBl�T��mjt�D��/(�H8a�/��;G�M��`�v����n�i�@(f��\~�A�� e}yi���J�κK;�XҢq斆��w�7��l��ѯ�p�(��]�Gh�"��˻gtEE�v��w�n�Ѱ�5�Z&��7��Qv3|�&��ՌR���LsКh��V�x��I����YK�Qe�G�(h��L�n�Y���Nj[��{l�x𝓲�jfĊh1�b��"�ƞ7�գ�'){6dX�,�Ah�Z��vpSN��,z8�X[��vI�S�o�}9���7�)�Y.Lp�$1��@��,?U/jaN�r�ST�<��f%SK/o�H��F�T�2�t��'a�=���n�'v�T{�F �\��@��Z۫k��v���z��T����S��v�<�3�wx`�h0r��&�g��k�9l���d�#wt�є�@4�v�=�3V�쓦��Gp%go6l	h�R���rd���DY�))�*J��0w;7[��¾U#],qhlj���1��n�wD�+ư+��ˊ�{QYfh��:��;�$����6�D�%�VuTBt��jbn]}�v�&�-Orq�\磊a�@��v%�wu����tn�`4��*��ܸ`%{9�!�T:��8 �@�Ok)��d�J9r|��7���y�ҝ#�Ia�p���npX ���C��CU)�4u|����P���b�h�FV�n'���S4Ϟ��'�T��C۞0,=:3d���犻[}�Az�e��Kw���v�%ēŠ5:��Tj����\ܜ,ǌ]K���xr@�±F,���7E�`,�8�I6n(u9��F�)���3FB��N6�u��u�Uu���.'V�
ln�n��F.)u�К��-!̝�t��uʖ�K��r��2���.�S���ud͌�(ל7떳�3�m�Z�~CTI�U�Q��Y�ܶ��ςwkڌ�Tl����>�h��x"�۷fn1� ��͓u+���c��u���ѽ�Q������`=���iãva��:s����F�L��l��կast��������4��q:�C�X1X.غ�Z6F���;�1��oz��.�h�'��҄�ޭa�z���; lӽ1��*ۉ ��5w^�e�S=�y��G�i{�J�|ɯqr͕�����ˁ����y(�u��v�ΛS��[�����SӚM9;��~�&��B�ư�N�	!�c��x�m[rSI�`��x5����e��l=�kRV%��խLܒpi舜���Ou�&�s�h�x���&�g���d�Ga���0�s�'��gk[�As+�8;'ay�����{r��_�X�68F��Y�s���jİgnj���L'Mt�����^_��y�Ew�4�w~���P�I�,f��;g���.�⹻�8�{�L'��:���ޙ�Z��k��ggh��e���uU���O�'�0�k<,�ov��h��}��v��;�L����h��o����a�HR�g��d��� ���t��5��82GV<�A4�Z5���M�W!��k�w*y��5ac���������SN]����Kh�����mG:k
s�-�&J�j\�qQ�i��h`��^�����v^�o*y�@�T��0ՒhnlD�H�z�4�����tU�^��|4��"�	�l�s�m���t�ŵ��E�h]c��#q"&�9�=Я����Y	Oow�1��(mM���U�E�1�k6ƹ��@�n���ŮgM<yQN��,��P��'V�Ǹ��=�}7A�M�M��Y�[ߜ�Jp��צ������h�\�|�Bc�v����+���ۍA�e���cz@�-��Y�/��k
��e�e�d՚R[��Bޛ��]���}��7��#DF�� � �]�)��`��ʷ�ir1���e���_����3x��R[���
�g!VbEk��V f,2Ǽ��7
[�s��1-�T6nn"ͺP<�L�t��d�S��ٳv�[t� Ro5v�)� ݖ7*/�^�s�'�[���[��AP�ٔ�o4�cND��dM��{�%�7I��/S�*�I��oe�>:����bΜh@|�0!;ϲ��\�՝,���|�$�oX�tWq�ዯ.M��׋�wm�l�v���I�����96���F��c�t�l���p��N�/-(�m�#f�r��8ukol��x�&ǭ�b'S��]wx�;��9�ŉ���}ܚ��$�
L�I8_�����+On��'.�ωeǋy�)�������D� 0�b��unv��7��-nĲ,zl5�|��;ܸ�,
�s����}��P-ۜ����"yi5\�W0-����3�J	�RN�8�T닟���-�;V��OSbM�Gf��`��ٹPm��)$3Aݏb��r��Q�jX�x�aw��Ѕ��RތH�v�GQ0�7x-�Fua;gi� �^��\7-�u�E��%�r���H �n^���&���A"�&r�E`��Ǧ�g�S�n�i�p�C�h)��ǽ%���[j��Nwn�GK�����<�Ҟ��J���|�bë��>`'�*u�ɐ�G �Lf�{��Ր9�Ud�w���2���mw*-�y#m�f;�/t������#d>��3539���/�o6/�vLӳd�gb�4Fڊ:u�ٜ�y�[߲�ܽ2f]J^�x�$`�{�H�i��Ŗ|iXF�6���Υ�u.ǥ�!rHvmzݛ�s��̓#��ǐ���`lƉǽ�ӯ��{݄hU��bL�[XF��A�8z݉^���<#(�CZk���0u�K�W0l�SS�g�s�������77
%�}3V�ʏ|OWr���+�䴮K��ܳ�s��m:�!ƫ7�!5�Ht�X:�£�v�-u/{N�y��U�t�}���m]�d��8���˻���Ҟ��'	�m����\������W6nsr.�7ٯ�l@K�FI���L�I�.PKt;����U9c���:��N!XnɱNPn�8��x�F����i�r���kJ�sx�l�A!�rn��M���� ��t>]�+���d|���ƒ�=��d�(�R�M���w{L3�Նn̛i;*��U��[��˸=VօכA���*Y�T��"�́��ˎ���5�r���-�ę1޺�kہ�L܅����ި�. ;v��MǧwL�i��W6�oj�j|]�ۛ�w��n4q&9��ݭ�;A<s�d���*1�r��swqgk��#nw�9�5-��иUA�����N�Z�z���;q��ʺ:�!�Y�y����{��92������d�ˁ�S$bB�h���U�϶K���7`���kM��d�`�e��6��ʦI��Yx ����vk�����zy@��$��씹Z=�(,����5��y|�ݑw�&E���(i��f�l�3���7m��6%���F��=�V%�d�6LO:F���&�MZV��-�G/| �6��xl�s�e�
Ż \�;��8w+�q�{��t�oc�6���pHtq]�y���:̵u��_����ym�b}N���܈}y�7���/==�yS���n�ӚѪ�aa�uQn夒ܮB��f�	�5�X��V����2u���tN���N��☗K+eG�v!B~<�z�5�aZ��x����/���k�S�p��nA��U�oY��xޡ20!�L�༗4�g>Ӹެ��պ�I��i�3��{l+�>��͇�Y����-�\Aey���FW��23T��3�4����	�:���m�)�Q�x@���pN��q��7�kŦv��9���.�q��GE��U�=�p�U�d]�xZ�wEø�a4�������8��e��=4����泫�;{���ͯ�F��^��')�y|��`�-Z����t��p���]Ƿ{5���;��/ �`�x�d��&��믂�i�cӹtk+��c�F	�\�	��^����V����&:����U��B���C���x�gr��Gn������v�ط�:A�Unp0������5��^m}�J������8���˻�9��Z�y��Z�l�̗�2,yFFaoWp�֫�k���.��'<�He>��ـ�k"0�E�_A�';goFG=��bZw��2.sF�Η�����#@{�٧��<N#nY�������Ad+7{s�3��FD�|�iA��⛀S�[�x^-�:�qُe�,4�,=����{��Ֆ�sd�C�1w>:q-CN���%܃X��v���d�4qzMaǦW�7��e�0߀�[�nzIݏ`�{�hM�N��l[e
�#S�y�.��$8g
9��#+ٽ��j�]�Z'r����L+5�ʳ��+_X"�1�r77y�i��7a�E���,P"V�f�_D[�;]�Zs����3�z/�=��}�y���VgZ!z�}w������R����P-�`˰K�d�1"�=�a�Bඑ����´NȐ�K����7:���/&q�����#É-N�c����d���t��9w��9v�)q�ӭ��<��n��6v�l�(vL��{�-f��.�6ݼ��3t�c5�i�L��^�z
�r�����N�ag T0E-}�5��Zc14���g^�f�QN!��w|���p�9��~KOlk���$4�;���:�}ٯ�m�ns1��{�z�ocn����Ŋ'ǣr�y������z�FjPфȸ;Lg�����cm	�N?�%�������rFjۄ�'���us����ɛ���8��+�,�>g)F�F)z���i�:��<cN3j���	����Bpf�;��zZЗ;:��㽓��$�����vǦ�6�6:m�N�B�M6�6�#m4�i��4���4����q�:xm����t�=��M�Ƨ�_�E.� ~�ޓ���>�r�z>�y���L���w��Řpf������\1���;Y ?�i�58�E>z��R��s_j�IJ����_|�vtk�,�y����<��IH��[jƶ�Z��գF�UF���ƨ��j�[UEjƫ�bڬZ-h�lm6��[[��E�h�TUhڶ��Z�kEmZ5kFը�km�j���F��kQ�X�lm[F�-�E��j��Z�[F�-�֬���m���F�Z���Z�mk��5��Z�-VƬ[[Q��6�kU�*���j��Z����j�ZڴV�Zح�U�Ս�m�kj*�ъ�֭E��V�6�6�mTU�*��E�mm[Q��UXֵF���,��H2*/Z綵S˲�^k�Λ��M�8>W������	'=8�����>6�~����4�橇m�W2�c�c��~d��¨+���  g8�w�r��>>�@W�b����=��_�a39���&=��� 7���.��rn�]M�w��s���w+�*�o��:+�#\������四o%�d���)����˻�|z�ێg#\PA��;9ȟ`:f��<�/5�x�`ea�S���p�s
�Y�����][s�1N��ٔ����M�V�!�h����s�����S�����+�_{��v�ޡ4���{c[:e|)��2���1g��٤���g<��F�:@�0^{�<6m����=��Б�$��@�����S9����O2��V�M=� ����%�rh���	d浿$�3>�a��J���R| ��XP(E�Fy�<���D2�;r��`��^�hК�������1ݥ�]��F��r�E���+!��<q
.�����NĬ� �9�ɫӨ��6wG�j8�
�v�C��7�.�)ʁ8BU~��T㌚1=�3�jN"���p,-��ǝw��޲��]怪[�{����j���	�7�l�k�Eq��7��/]��X�g�n�'N�N,��>����<O�yD�c<6B���C��VΞ����m>�v�Y�ّ˼����RyxbE��|��}���=�(�"Y�J�'k�c�~>;}�R?zwԁmx��p�ٖ�Ո�sE����cja�1���Ӻ�q��\�g��^�y���&�ad���aǨ�l�(7*�5Û�o#7�z1���Ǚ�$,���	AI����"��1y�<}�� �D--"M�A��b����MB����;ӧ�˺�+}�w;�p��K2�o5�ܱ�T��}���[��3���Ý�g�}{ěM��U�τ���D,��޾}��������Z����/^얤��Y���JnY������Hs=R�|��"^za�Ӈ��o�v�?v?,k��y��M�}�%���G[�G��k)x*N���^>�Ѹ�ù�v68���8,w9�׋>�D�)�����t�vl�K69B���$c����'�����Op�E\�͌g&V'�g���3�v'��!�����~��:��n�.gY�轡	����o���1��I	��Kg�g�
ؘ{��5h��$�#=�A�7Sa��Pn@fp<�"//;&�o("�'@�5Y"�OJgn��!n�r6 /��������弴3� ����}3��9��Y�趇����_]wI��[��A�}+��W�>W,��I��	zݾͨ�OX�>����B����Y��+����hV߄�5s����]Ĭ�������x'�ɱ�$�����xv�m�����(_<�vX��I���8����7�����4�
���3g/0=�A5���=�{�\~��B�^�v��xj�I��}������%�wn{���-�ɐż���|ɵ�^�6��5��ӑ��'�~[̢6����L�8wq����3��xl�
!���>ʡ�%u��¾��1_��z�^�A���も��g{�"ld!> 6� �	ǔ+u��6��xzw�u�F����~G-�3�t����_7�|d�� ���j��=��y+@V3�E�%�c��?i�{4%��x�Z8p[�µ9�)��q,*��/j�>������m��ݳÓjk>���~��sۢ��j<N�4����o��/F�Hdy{:Z�3�(*���L�3I�9|_	C�n&��h�y����9G<��H^�j�c������\w	�im���^RMQ�I�� O�?n������{��	xK=ػZ�D�`rN& ��eZ�#�BiCY�Q��ܹ�U^���v��#jΛ�����u�7X�d�-�P�̓t���&��7*}Xgq��+[�Ч�X��ywõ;gF$����e\ӻ옪!_0n�QfyJ�o��'��s��K-p�
}�t��=5=޸�=��~�}R�]��r�9x�Jl���|TԲ^.wRfޱ��$�m+p���@�o���t�(#սɟu���ImX<}_�'��;�-|�C�]�I=���;�
�z����g���y�D���{O��]��=�s�$���9�>����ӽ�[�{y��:�-+�(�c9>��UI{:y����V=�,�=��oqYuqBr��oE���-�����N�=��<�<us��3��*���I���op�G�^�2{w�Ź�K�s��ghy�L������}��-(��@Uk�1G��Gx�wBa|��4ϮW���#�F_g��b��bou{|jõ*���������R�-���F�>����N۳�{a(��/E����=�z.>-'���	�Oq��8-��}l!��8��+�����]˪�&�ݮ�zN��� wpf� �N��ec�`���B�z�j�_nu�h����L��2p�����m|��㻐���"Ǆ�@Qc9�[�-i����]��9Fia���=�ⷽ�͚F���)\`�-�����wW;�vn/��]Ü,�A�|}�3��y��l�F�����62+�R��75��ۯQ8_T�.n���7��o_9��8�"���,�:Ʉ$*{�jMw����#DW�9�'�r9{L���'���=9��{��T��_=m�.�x�����n�k/. �'*+6?^�;z{-m�ߑ�_y�A�ݏ{���Y���W�:�d���n��������Ȑ�7ۣ[��!���Y���34A7"|��Ug�r���?w-^{y�X��#�=�k��=���[_n=�=�H�OW"��9�v���N��|������`�;�w|��m�&��f���y#�;�3A���>��I�;[��w7�yvÖ��1+>��i�.�CBv�((_6��N�|.�V]<\X-3ڞ5ٯ�����y'��5��� }�Z�|�'���8"=�?{"�4��!U�Ac�����m�����\�^R}��x��g�Ok�e�'��v�`Z]��6��C�bň�,y%�G��A;�����p�{�C@>/e�noy����{e��b>q2|����Y���܋�_�+*d�>���a }���Ξo�y����մo��wuI���W���YY=f-��軾�R�&2�G�n��	f�>C�yM��^����t�/��2��95v��L��W��u�z��7<6�s�߻�_?P�M!.������7Ңl���t�	��ȍk�\�r�nGu����xG�:����b��w={�L�˚��w9sG<�=�����_�&�||����j�[��G��������G{_�	�L��=�y��h���)�F��j��O�z`T���~'7�h���uD0��:�u0b�>#шԛ�s[֍�zg��F&8��7=��a�- � P<v�Քg٧q��ͥ��\��<�zj�C�=�yd<��k=�N�g��j�HS��Sؒ�l�MqY0���M�Y/bѺ|}�2ISP���c�7�4�*�～��Q���W���{p�({�rKY�g���A�#��tE�g��`��v,9l���g�[��hܙ�f���z���I�{=�R�g_�-yxZ^=�yOI��|��Y��D��p"�+��c��G�/4^�4_�;1|��S}�s�w? �!�s� �a)����b�T}������a��{)~��d�ܰ�;(��ѕ���ZkOo�sT^�����T���6��=�{jc�,�δ�o�i�w<���{4q��^����w�g�-�����s�	(�ˮ��۝؆���%�QbrЌ���L�*�A��84��� ���q.)��2L�a�&���J�z��7˶h�:y,�Y�$\߻Ǽ��/��y�'gg��6�*Xb����.�-yW��� �@��s��Pt*;�����w��Y=��`Өҹ1Yt�f�������Z/�~'T��jQo�f[�׷]{�?�;ئ�>R>�������x����c$K�8�Q��r2�a�-�O���;�i]�7}���Cա,:�oL����(��^�n���Q�7�%�<8t�b��=�y��^Sp->J\*`��몡����.�DFk.�}\��⯕b=tL>[Ek���>9Gm��U��Ny�����U��9q+ږ:#�)���Y
zG^��\���F�6:����x{;�L�#�������J`ޞ�:19=r���3�-�B.������fw��I�Y*��yt�ϐrg1�b�	��
S�B�&Mܻ<�=�m�Зr���n�U�gd�F`x.��X.T���S�>�0������o{N{�vY��s�{ʲ3��=g��𒢻.�a��}zg�( 2y��rϞ'C��H���h���z�Os�솓࠵��0oH����4E�0�����4n��=�m��n�O�	�7�7�ȉo �t�����vF�� ��C���>����ɗ<�'��J?���d\�ܡm�tݙ-�:�q+6���ڏN�C����:kKJ�Y�B��r@�N�.�W��La���ÞS;a��^E#�V�t߸on���[@�̇���R�5�W84�%"Y�ws���a��� ��_x��2l����s�C 9~�jw-���\��ueZ���=���n�����V	{SZ����Jp�B�H�E_��J���lE7���d ��;o��#�Y��Q�7M����=.m��;غRW��g�呣xu�x̛�xI�H����
�X���r�v�Y�1���{®��p����}�t2f��)1����y�Lc�=����F�Iۯ)�G�����G˽%�N�~@�7�:�hn�)_Q����ǡ�kKޞy�n��<V�|h[��)����d��� �|�M�}΋���7��]c��=�'{��^���׀�0nL>�8�Oǁ39;Ů��b�yE�2�;��H=҄X��>ң�����ғJm���o�iy�#;���*�{�#�u�O_��ݏ����[pK����OG�ނ��z���#=7L�/�rݚ��]l����㞮G���h�O�>������=�o��E�{�";ze
Dy���D�y���n��zL�h�kP%��ƽr)-&�T�]��8��
AY��.�j>-�!qI�pz6tP�.�.�,���o����~|������`��d����4��1��|����*���?K�>ُۈ篷w���{�u�u�4M铞�G����=Og���"�c��>��ȷ͟#؇)��{�f�!��`�c盭��3�n�Y���l9D^�Ӣ	��ݛ�a9�0��Ad�<$�F�3۔���{}_��{5u�w(��|{��d�3��}��Q$ ��Ě�Q_�G�^9�y-PJ��B����괓�zO���E�E����Y|���.$��j�ʠ�F�Y��c63�glL��zC7&�SI�2�J���'��k�t�:��:���u�vվ<*|��I拧����c&���V
�,��!���8Yѳ9������]Z&�n�/��M�1��v��v��E�.vĪ]ѝBq�b���Z���o ��l� ?_z�g����W��n�{�����t��|F�r�zG�t���9��6cq%b۩���y7r���h<[�1sI�縉���������c+ڽ�^5�<�\����}�ޫAO��
�6ߵ-�����hGb4����9�zQ�ˈl�w�h�F�hDeS��ѧ:�{��vx|A���wkw��$x��`R���w��-�_q�A<��9S�G#���7aY�2��^��{i��פ�{��8��{������=���{F�E��k���V:���cK�.��ojӞ��dz1VK�w{op�gko�h��w(��Sf����=��{��T�'}��d�f�E���Ǉ���w/uh�|�޻��"�5���j�b[pu�Y��a���G�{7������{�f�b�}�^��^�x�y;�؂:��
��;�$=�������vw{m�z�RH�Zb�F���g��_L	��Q���&��#3IM�L�R%4�Բ�
!�g,�ȉ�ۜ��F�7���_������I�><;�'"}�
O��wr��Y��"f��!om�EEg�~p�cz{_B�Za��;�o���j�泄��}Hr���s��p��7,8߶�<5��2�yK�;B��y�#ޟ��������Cs�vy�v�%�g�*��U5���6�x����E&M؋��](�yzy�.��t2%���0x��<�z�|\�����5��!DB�逹;����O�W��֏n�N�m��{݌�������A.x�6Z*'���Fw���簭�H>>¦�m�5v��:ӧ�/o��n���R��Q�c5���7��cF��kVo����z�&i�W������4s� ��z�sxM,u��O۞��u�� �P���O��:}u�����`�� 6��{ǻs�҈ ��w0�ӂ�+��z��F읣}�����1
�^A����	�{������yl"�.��8;ိ� �w"��_)�������r���S�|0uo�eߎj#����j���f�]�ƌ븅�>�-S�u�:��w����pK�����;�d����&��V�g]�]�x����\D��|�<J���)�
|�+�S��S�hUfr��x��t�w�Y,�����d�^�;�5^��y�лl�l���^�Ǘ�4Y� ��K-T�eK�pJ���*.����t�yUךx��/?%�R�v󷦏_g��|��Fu<<7��aN��ef�I�;:�׾�{��N�|Z�E� iT��N��k��^�#��!�yf�kw��gz[1>���a�T9�8���}8�0�������Aĭ��ś�����M�.����cG��2�!c`v���]��M���b�"1������ݼ�O�
������+�c���\��3q�طGE�w����O�����AE}�'���������U_O�������~/��\�á��卺c�<{�{��m�UUT.jv�������U�^\nX5�.�KvC8:ng�;$ջK�7�z��Mzҽ���/Vvn�ͺ]�i-�E��9�G���f��Qγ�Z�NG��ӎ��t�k���x�3mZ��&H��t�x��y:�v{���.ݧ�vg��ˢ7c�ub�����'-^�7q����I�:<�m;ź�,m�{�s�o���/�w�|s�Kn��kUɎC{�����=<i�p�������6�6�P,��v�ڃ��Mpz��v��۞/qŷ'T�����O�rnt�x�;�{=`��tn;B]-3���z�x9�v�J����Nዂt�Ŗ|8;F|��\:��f���a��ug��{���s]u�L�]˶��nu<��r�1{G�����vR�7x�uzŹ��Iɶ�ȑmϧr�W�I�m�᭪��b�܌`
���d�0T��u����n҇;`	�s�n=�aۦ�5�i�z�6B]�r5�<d�Yێ<%q�ָ�C/h�.6���J��Yu����6�WHt��$8^N*L���l$P9Sѹjnz�nݰX:�/NA	�^җnY�T�[,������#6�7S��u�Lr]�\���ɫX��ޣnJN�O��A�:����\�ǵ��c��y����Y��\.��K��Ɖ�����y�8�6`�Gn��q��s>ڝ㎻��q�z��8ܻ�`�>oo���</-�����k7��2{�n�z��X��!�X�q����u=mvϢ.p��`�<�ȼ;������{Z�pQ�l�+�֯]�y�,�c�k���q��bI�y �ێ��<�۵>��&wj��\��c�a�yZy��:�wmG�X�������@/����;���D��5�pVj�q�b�gO�\���P�/Q���G]�����ÇB`ӂ }L�֥��͈�q�ع+�G��Ol��lx��2���v3���5ƍcW@��!6)v��a�Xn��\[\`�������9�g����&�݁����,�]�'3��F�K��}� ��f�wR"��gv.:^Q�;ZS�IoZ�Ö�un�7t,n�=�A�L�[���7h��m�"YN�)�]�4��wE7uњM�؁P���3Ѱ�nН���6��96�x��r=�ꅞmlNn8;WktU����^=Ǒ�ن���6����_�O�#���s�piNF�������.-^x�snֲ�V�Eq�A�^\����=m��=�+��k��P�`�yuN��-�F��76{8�ܜuϷl�a��c�t���6�i�������]���^ݴ���Vz�ۺ��Q�v����^��Ɉ�սmf�B��k�%�]����|\��~���Y���(�k�]^�*�Pg���Z�і۸�ڄz]�"��q�1���d�$�c� �o!n��qnz ��<�7��;����:�B�����dZ�:^�n���:�G<�����v�ւ�0x��'�8�\��Df�8.ʈ\ۊ��9��X�]������|5vw-z�lp����ڹ +;���b�]ơS4Sݳ��l�cU�V�b;u�5ַ=�v�Dm��n�׵h�Z�a��v�>ͭnA�ۮR@B�մ��j�f<�� �9�E�cܭ�!#�O#���J�tq��n��_}�׵�nٕq�#&�W�E��X7��v��n-�%�>5U��C�E��lxӞܙ�Z��X���g���u��79�mq;���mj���hVvL=��N��[+�.���gF��v��<�e�{u�xw%��kt�ў9BE��o��v�g�����R5�er���z����g�rs��Nc�:���	%���5���m�M�Ξ��C����sN�f���3�û�����
D4��sg����ۓ!qbE��c��w�L��h�[>����rn��"�J=�5�Qw2�/I��e`⺶N��x
&�6��~G��룤#��p�jz۪�z�\�V�luf�tx\�>z��-�N��e��=<ѵ�R�n&��[��<f�<��;�����̝�9�벜�2�֍c��qNʫ�K��F�f�%_kj]Rk���] ��u�����a�ݲwl��mr�c���i4����� s�؝����9�-���M����fZ��η/��X3�{O�8k�eH��|��\����3�*x�q��*q�[r�uV�'�ⷞ��s��۩�l����k�;i켛��f�¡v�-�7����tpZ��l�!��ꓝ=�������]���1naB�O�b�⻳�R5��불|��i��6�<&sWOGf<v�tB�1՗U��lUfY��ں��9�]l7(]��2<�.M%&7�̴��<cq��i�q=Z�S����ܝ��׀u^��ٱ3������p��l.����q��Xф���Z��tY{wY@2���{
m���>4��:�NFy�ܕ��G���sO7�8U+��غ]u��`��4�6���$�[���X]���<�ܾ�]�$�x&�sJ���j��ͱM�7���׺���6����] "�P�Mִ�����;�&�b�`�ړ'U�ϳt��B�����`��1Ӌ���� �K�3�Ԩhd�����j��[s�[���˶��73W�u���P}��q���u�A��q�Y��o�������u�؆JB���s���XN:�h�N{W6�󱋵�h9�]�Tzy^
s�,W;>{,l��ֵnd��˞�2]��n�����L�R�\�U���,����cv���::-j�9���!�#���,y��(��x�?qY����b�#�2͊�^�ƻm�^$�vd4��F��l���}�F��k�S!����G��x�v�v�!�'cQ�ö�h	�x�k��vNˮz+s�e9�	�n4�n�۷�X�<i����i���v��'Hfpg�w	�p�Y���p���8���N�x�w�%
�n�����[�gQ��Z�ݞ8!�q�$����/1ĕ�c�uۜz���wT�w|O�O�)OQ���m�TiS�Q&p�;c�U���~	窍�;F2黤c��;a��_|��;���՟Y.5�wn����1Wo�/E��B���xb�v��;7b뤞6�>�8��6{{U$�r'G1��/���<��h������nX����wꇵ�km�CO:(����yV�z�*���.�q	j���wi��W�|vգ۵�o\�&����n	;v��눨�s����i���-s��S��{˶�V�7��N#0�d��/0C�v5]ü��ʼ7��luK���X}E�o4��ۛh�j\�t���9�0|�ً�n�#���<[d+���{=	n_h
Gf�xI#�e.L���tv�>ݮ�7<��7h�[R������ѣou�żC
n��T�=�@��2I�a穴9Krq�gu�n��
��m>&��u£�n��in�=zڇ�˼e�+E�۞���m��Iܛ��u��3\t�����<(��L�M�n��ٸ�/��s��O^�9^�K����ѭ���s#�뮴';p�i��i7u�_a��"��[+۳Ea՞��<��RF<�%�5<4gl�����@ڎ�p�n���a���l���i���f�ש�<��'bw77'3g���a��ҁ<m��p�Pf����AR�|���g��Gg]mp�]�3٦���s����Q��t�۳�����=����hv��$��郛�ბJn1V��[�� ��a�E4Fz�ě]��g��v�z��rr��S���DǮ�"�s�#zz��<���8{1wW^�0�u�p��s�n���]�`�xwX�Ρ�H`���6�{�^||�}9�!�;2#��c�ʧn��j+�ݹ�������\��!m�=t���������k�g�ܸݫ��f^*&���+�D<����ˮ�!֫=��1ij�|oW}�8�;��:�n$�D�j��ְ�٥��{bWZ��kP�5nh�B�3���]���$�6N����q��u����1��9���ݺ^��]�2絈˽X��ݮx�o+um�z˵�{Vsu�fu�:���W��y*�ޔ�s��uwP/N�Y۱�<E��N������y��G$]�cWs&�o#Q��8��/Jv�v�Jtt�=v�:�c�@�O��G���lG���6(o^����p]��b⸷'n���8�]t�n-h���&�a��Ǯc�*��ׁ0��\�!v%�v��5�l�WC��֕]��.=n�ӏ^Ҟ��d�jp�El��]m�n�R�uĲs�vԐy�)�n(8cr�q��9�ܲN�b�=z�v�ps�n��}=I͛�O}�_rngP]�,i,/�.�u������t���%5�F���mq��[��[��E�XN�l���5Z�^w��f먱F�6û��x[����K�ǋ�F���X������t�V�N'�����4�nF��nb�k����	�[�p�l��q�c�׶K][��/�q��:�ю'`t���H+#��s(�����n��YJ�u�Y:�����V]O���x&��V���FK��Ev�`:���K[��[ulMG,�^7� �m���ɟZ��'�K ��9�x��nqj�#�{:�����x�cU\އQ7%>�m����b3�����9������X]��]op�sۚ�b��/^|��C��秣#m&��1���\y��uhmm�76�a�:鼼;D�M<��BR�v��i�:K�d��\�-�{k��J��h����kݭ�t�Q�]WUv��]n���-�U�Z�UѪup�mi�-q�ӛ�������j�u�G]�����f������������������D��|��}��|��y�aA��F4Dk$j���������Q]�i�ڹlTZKx����U��D�nh�F�b�Z�_m�׍W_�[��5�k�4X�m&-�^���E�mw�x�mm�FlQh�(�j��*(�F/�.j-���k��ۑ{sk�IX�cZ(�%���r������$�J4b�3c!�h��\�Q����Z䑱Dj5��}���h5�ߍr�c(�������d�SW��N:�^�Uz֡(����k.n���Q��W���o���y.v�ݼ8��H�խ�\j��x�2�z��^Z�v�g��ꥏmy���=�4���M�t�ׂ��X=��<��i��u`5c���]lӹ4J��ݧ�j�B[�1����[��d+�c6��m�ݪB�˕���������x��N6�­�������[P�9ދ����{�㍻�n֩6⠺��ѓ��\H�p��hު�[���U�N�Ί�v�]^�L]^sjֹ�5�7�l���c�Y�g����i=���3�ԁ��ݖ;���m�7�$����v�Ǖ���2p�e��^��+�r�r�� �nq�xcilZ�&�v�-n��Z	�jD�ţ9�8ޢhy��X��PQ<�s��v�����κ;r��p�����x��nB��{BŁ��.x�W]n{vC���g�֭ҋz���ۆi�����غ�u�i�A�h�[6��v�X=^b5u��]�8��n&�Ǎ�k�ۀ����u�v��WDt�Ek��Nx�� kz�U�u��=lu��=�a�����IkՋ46�I�kچbN�������� 1�ulQ�OG�\m�۳kcT�%EΝ)�@�io'��LY)�li�9�-�����h�v���ѵ-YJ�K//Fs\�Y9�Y�s�\:�E��nL�
���3��f���ςg��݈hnT�.Zv��c�g����q���qǵ��ݻmuz�6���	�E��냶C��Cq�p�m��\N�h���ե��pn��`´�:#%">�!,s�q�3�u&򻧄Fy1Ŵ��lv�/��6�8:0����{T���s�O/9�=��q�X��M��൑���Ia�#Ӻ�/F���`=�������N�\�����u�+F�՗x����.��r�r]]U�8��հ�uUUU\q�z���y�S��=��rw4%��nC׹UǙf^�|��C̷/��[���S�[�y���|\O��$��H0�q�wD�B���/W#�Mr���'Ԡ��}x�C�NQ�U*���O���W������t�r\��N��)y9��G����E�����??6��񱘺�v����6x;x�;%�n�h#�I�%#�3���񶬷{�� �ڮ6yǜv^�f��R�����Ywsv�]��LdA���+�9��3h�j�m��9)�j������<
�3�/�6���㽧�?�:ܜ�ޘ�׺��i�����xN���v����1�q��٭�.�N卍��w���S����F\���~
?����Z~��m_ZJ<*��>���}����Mܧ�_���m����0g�_�~��+�ebxH,�l"MWh���O1���h	��A�e�l`_3�~�j�;��n�uNk��ٶ����|��Ӛ�5�D[�f��u���p��.˝���7���ݴi���^X��io� 0��}�Zہz��s,�o�����jE�`ջ�`Av��&��.K>+|%����\,���؉���W��_-ǒk�w���/
lY![_����\��6�j����6N(I��6f�Se�)a>�����a�$��ƅ�	1�"gP�[va����U{�f���)9fmk�3�m@K�W��3�-�>��i�׾��5��jM5���:����[��}ȷ��i�۪�;�m7{O��L��5�^���\�h �#�n�̓(<6>D���)``,]�q̷����`���u�F�]
d*�=f�qmC��o~9��_Zm����x��~���S��p��v��U�ĲY�bgEf���Rg+gf0E�u�+[�mwo�v�8�>�yM2����p�)ot�k)d��X��ݳh|zt�_����Mf��-w�ѠBU��3�������6�8�{���5�n�'��d+1��ZK2��2�|ˋMv��v�l1�c����ۓ�X.�� ]���'ef�F��2z ��� mB�X@�t��]�v���f;�2����ҬQu���`���V0���[��������  �z�GK�]������O^N)�>;n��B43���Xݺ�g�����ߏ����|.�>m��eo���e��K��EiN��Z�7�{�2ڳ-�*��{S��U��]�9lh����D&�B���q̔�v�����2����m����k������Y�82]+WT�S��q/�����.�]����vۇhd7�޿��>m��uo�k_2��%�]���|:3L������9�d��N��k+g��o-�O���|F��C��#}�*��`�Ǳx���n�{P]��;l���~̾����>��
��Ҹg���qR�0��E�m���BV)К�!0m�{w�?B���M	`'߃ǌc-��bzb����n:��S�!���!��X�"��P����Χ-�v�x��WS�sS3�oO�h���e��4`��/\V5�]����lj�Gf6.n�Mk�z�zw6��-S��)��_ؘ]��|��kv�xq�u�wov��35b��kPٍ���'J�:[�-W>.��.�]��aݤ�+w�,Tz��[z��<A٥YG$�&Y���C��c�j��HzS����ܻ��`*���S�f'������w>^&��ܸ���ݽ����Q�z���������h�@p�1�����`�zFw��<ٗ_�Q^2M���*��^��7'w��v��� $���-oϿ��|z���>�x�����&8ٜ�ַ=�ݻc[��n;{�.wUc�g�;m��:<�\K��.��]�f9N8���3
���r��t^:a��U{ukZrIt����vǷl!�N�p8W�(!;t�-��p�Խ��p�3庆 �'�,cd�v⎻p&��i�\u�:ؙ�:Ӂn�]��ꧬ.{s��x�c�8�P��{0��f�[�����|�/~q}�Ȝt�Ms�U�qd��"��M��[�݅� u��"`����M�p.���4R���ԜBB�	���0�z�d�Y>l,z��v�ް��C\�գj��k�}��m�N�Y���Fe��y��RvD2����b���l.����u��ӗ�Z�D���������S��j��m6�i쟸N@��젣_5��`74R�ȭ�)�!6��ݦ2IsЇ�읫�㖟�ھ���#hƨf�.�"��l���Va�{�3'����w�YQ�J	�C�}u�M�zb���q�k=���uΒկn��9z�m5X���E���xв��S�V$��2�[Q��f 7-o]ۋ���-A^�eM�����Lņ��EC�B�CHS���.��=��e-���%�'�pż���W��V�����!/�d�}�/Z����2�;R��)oU�wQ!���lK^�y���7��v�=wtT_�/f�D�P���VvI�I���Ui�Ӗ��ߜ0�=��X���;�2�ͻ�u�opڝ��W�SZa3#��S��)�m�����]�Ԥ��*F�:z�'a��P����E�J���b�z���qv����X��K@���y�;����]��!�MY6^�8�ޮ�l]9_fk�q���(Oൽvޫ6�T���b�kj�~;FC����,�/���e����̋�XY�f��[{7U�\f�\j�zĒ��X޻[hTC�m���5���v��o�R�*]<[��n���VX|�8ވ���*�D���7	���tkĬ�	|kgY�Ѝ�ݜ�Ʌ�׵4Sˈ,"H������4	�Ffնd5ŉHUhl[���oӻn6������05�b�d��[���o���Mt~�}$=���N�~�M�O���vۧ�h�U�}ۊ��X�S�r���6g�t�~����h?� Z����>`7Z�l�W9��$A�q�����	�@M< �O�w��,�����]��%N�{���$*�'�Nm\�ї~�ofc���޻��YRa�e�X�Zf%�3S�@קW�0��Ӎm5�X�ܷ�M��˗[:��͞�oW�p-7��]��]�4km�N`J�Mݾ��m�jĒ��ܺ��O�Ֆ���?xʨ5zLO�3�����Кw(ъ,:B�nXHNn���E�55�{`��;��ދ#�;�3�:�`�<�̄�<�����̜|��.DD:�-g�O�g���{w��m�t�v�ZL�Ľ��Kk�ڲӖ�K��_�H~��ۡ��S�-��B� me܁wt�����/��_L Wc�PD���O��Ӟ\���/j�4�8�?�0�<j~���O����p.�4l���UUh��Ē��#HӒM��>^�[x]�ݷ�(���TW�Ac
M��1�r��
ä"���awt����li�o��v=Z��]�ݿ�9C/n^ss��������v��M���mws�l�U�w�y��i���f�7Z��EE�$�o����GZ��X��m��ݽ��͝R�M{��OY8���.��9��n.�а�=���	�<N���y�b����Ԡ��l���ö0O����XG�i׊lLys�-��1b���Zp��E���CVO�a�ۈ����T=CѬ�uں3����L�R�dwOg��A���������Bo���̒E��ܢ��Vv���v!����֮z�=�D���:c�苭҂�QK���ONz�ǝ�ڲ(���ƻ2�3�N��GI zh��xԊ�n���ꝵ�ܕ��{:�^G�:o"q�n�%��Xcn�[��X���b���ٮU9�[l{��_��ܘ�����Lպ�.�Hr��u��|���/cE���, �����觭ymH�H3��^�=����;5��&�]"�a�Kv}V�w@\�ٷ���X���|��b�n�MV
��V�h�T��y!�C]]Mj�I¶��`.����r�����)vC'M�B��7!!	Y���6�\5ݿ����n8�,��Ɖ,10v��&�8���'a������GO//S����֜�m���R�ش�vLvmf�B�mJS�Jwª\bk�۟�u:���_�u��Z&�!� 9�a�n..�h��5���O.��U:���<m�,}}w~³]��ٽ�yX#Fd%fQӡ@�f2n6�ՍM��]�^	8I8o^ù.�P���\��Z�31�^B�x��e�l�D���Ї���D�a78��+���ь��x�>9�ճ�5҉�w�}!�.�ۜ���:O�"�	��lz�n]�T#$�A�A;,��Mv�v�]��d;:��Qyɫ�8�L�(�5/�<]�����3Z���s�q��q����1�]�B/rq���ږz9���O�mY���y<�ڝ�c��;���m���C�	�^,a��]汋֚�37�!��c<0pėh1EK��)��(�H��7(lQ6�8�����m�Ww ]��c�{��#qB�4���^�p���V�=n�hv�=wn.�����vv�e!SO��ln�kƌ�N�{����J~��=�'�q�iϽ��efQ��M>�8��۷�z���4w����A�Y����{�#,@�=C��K����)�y���'Gtɷҭ�-0��\k���ek}��a�<g)=6�9�(���h\�8}��}�泫�c<�W8��P�(>��X���<���dػ���X7B���Z�K��ɼ��i�
�;%���2{��x���,�w,v{�ڶ^����.y��Q�i��
�g���z��Kc,P�vdȅ>���8��Uٞ�Qٱ���؝ ��g��Db��j��s�)�G3�@^�����	|�M6#q��Bͧ}��9��}�׫4ő�^�?h��ͬOzN��롌�{2��'������n�c��)֗@��]�9�ozٹϻ=�yp�,�ҋ;���=֬덳}w]����菶,��S�SX��Tܮ�q=f�����)��y���~�/�w�g�����ٔW�X�w7���	]�k~&���N���\�Q�]�m��N�GL9���c�����X6�����m�^���V��{�=��g��ZY�==�|E�ٞ���O��nS*� �b��ǔ���V��F��w�Y��w&�|�!���Db>ͩj��3Ӻ��U��^��|Ɔuo�®$��q;�}���:�3Ad;��W���p[�;�R:��%V��]9n�z�.�90o>��1�4�w��=����kă��\����g��t�"��q����T<ۘ=��l.S�}��7�ܒX����ݻg$�wx���n9Mb���q�ihN�y��\B��/�c���7vd�F$����J���ם{�d�7�ۦ,l�I� �����[ŮTlE��.��<�mj�h�չFk�Q^���k%żk���W���m�ۦH�i6fj4���X�����r��h� �c��`#Fe����"�j��V����HhLF�A����%)�Ѯ[ �J�Q�1��m��Ib���\�6/��OK�B��~��l�Z�fl`�J晉��ι�c&ĔT$����n����{�+�D�ƾz�H�ε�
�_Ms�IA>'�|cߞ�9��l�-�z��
���k#�\AI��
N��@ŭ�Q��I���L �`?��"���	���s��s��+�R�R��nI�-�QW��g�_w��n�ǁ��g�	8�RQ�@׊qx���p�?�����[|/�/�YmA����E����q�	?�cmٽ}��������x1��c8�h���>�8��J�j]�N���Om͒�q���~>���9�M> ���DF5ؽʙy�?T4`�V�O#l�3�}����A�vǳ�Q'�����% @%&C�i�\�&_�>��x_���c_}����R�R��n ���یMx/��? 3������a�P �9$㾹�/{��з���%����}������^0rIÐ�@I���ٍMi9��s��mܿx���9�AI?�"����jfv���pp�n�Ʊ��^��f�b���.�fz8¥a�S���{�[�x&o�w5���d������u���v�Ӥ�*��ޚ�%Q���I����L��̱0-e�3qyB��34��+a��18pBI��
$��Iz{�[�P���5���K������&�n^֧m �t���8m$���6S���y����DbƂX�!����E��]���.�ݣ��z�aa7=�<u�ߝ����L� �݁&��p��_���y�e�í�[��lF��9���Fo@����
L��x����qܽ@�0��!�-�uLN���Yq�A�AI��Y@��@���wBK�^9t��A�p���G�oKG[����.���.W/	��KqV�>�8)3�)'�g#/"�Z��.>ݶA�\�RO�����e�n]d:�b�q�`�>���������<o��
L��
I�'&��3�6��tL��]ӻ��KtuT<��1Y��'�q��G^G�aD$���_�x�1Pƫ�j�n]_���+�<�=��=�ϵ��{~���}��X4�4�R�>�ɿ!�&�į'

������mN��Z.0�`�_��K�$}�x�d8>v�v0����\����(q1�]�<s�Z���9�ʋmՍ՝���4���M���/i���ywQ�	s�m�W-�xn9��&���q��=#��1X��]���8����y��Q��e˸M�㘇���6)W��x9�����Fk��kz�I�/�S׀���V��՚YW��ny���=��X������������~�켌g���^3ٽ��u˶9nj�x6e�Z��%��E|9_����`K�����)�J�r�_d�x��!������^��o9Z����o8)0r�({�g��L�c���w70k���!փr��Á'�-$����o���W3���ݏ��Rg
I�©�:[9e��T��OO�xEN��>5���G�aD�� ��V)�p���0��"� G�o>��w)�Ы�'���!���[���G8�k$s��n; \�Af�g ��8 �%I�#rsw�OL^�9c���ԣ"�i� ��'IDx����XP�p#�CQb�y����]NջrZ�xW;ruG](v�8t]A��g.ŋ3>5��6����1��ǯ;���y禩��&pp�ޡ"雭�3
>��
LIÂQI�����-�Wߞ�h��*�q��f��/{_��<�JEr�<��ŗm4�yt�[Z�)m�i.d]�ۖ�i�`��|˺c�3�Ay�.z6w�ꨏ����K�qУ�'���!���9o ���H�L��~h��\�X�Ƀ����&A�I���q}��ǎBB�泣iND^�iq����Rp�!%����H ����s��7j���*��m3��RO�wj�ETk��<%7���zp��h����!%�JL���I5�7��q��{��2k��ӡ?:h���!����X�����q1�܃���A٢�; C0�ზ��q���^��E��eb�i=��n l���[�R�����	�`� �{� ���	0s5��cGxuJȊ�m< ^C7c�D;'�{�a��G_@���3���1�gZ���E@D5N$��v�z���h��/�Sq�`���� �]_��e�7�q@�0@IÐ���	8�7fӃ�3V���׿Ӫ�۽�k�L��j��O.��{ �*�"p�j��xo��y7;��)8�.�ˎ�{�i�n��[�̝�匇���ɭ>�:�r��d7��cq�B��?�$�BL���!hs���j�#2�P �+���
 ���Y��s;�b�C֋�� V�r!D�l\�?2�~#�G����)3�)'��=���{�~��Ê�6E���~�Z������y�5�y�S��A� ��
LRp�{F�z�vq!�%��`<D8���ܷf8/C��7��Bxŋ��v7O\�������� ����G�I��Ƕ=Y�x��*W]��DD����f�U>��?��8�x�	3��LcKd�i/�o����=��[|�㨎�;K�D58�V�p�?�p�$��Gjѻ��{7��i ����Zo9I�����)�f\H�˺�޺z����|�%7A��� ��I�
NJ�����q��v��0r-(�8��{4V�̢Һ��Lf���tfλC>t�I�P�6��W�K����xp��?G��"����/{����@l�y�&"��d�Tx�L�0�1��~pH�w����f�<2��|�A;^I��R`�+P#�&Dgֱ�ԁ�ĭַQt�,����	 �o �'BJ#�$�}������������z�7l�I�=��l��ʔ�zў�T�
�ű/cvtX���~q�~�o�����%$��W���n��`���Clc�f��2�����s?�I�������u���%���~"�<u?��I�ͣ�ŋ)J�v;p �� �7\����N�bt<���	�`���� ���W�)���:�ȷF��S[����^�M.8�0r'$�I��L�liNi���R{��cI��DM�{rn�4�6��o�"Dn=.a���9���<��v��w�vrN;��G�p�$�s��{�e��>�2������J�W���|n�w_�
L��
I�-B�&m�<]��0��st�PYp�OG�f�ȉ|���2���M�f�Q�4S�G����F�D[��F�s�O���uq��{��������nђ���Snv���:�/,uӸ�n�V�m"�Q�ۅ���WF{Y�닙��6dۈ�������޹�\�ŴRsEv'��pq[[l�.)����\����ڝ=/�-��/Au�*�G��2g�]';�������\�Oa���X�����wM\.C��j�t�ORR��k��mx�3;o-n�x��n�]�7;�w�m��~�����xM:78�K��]v�[�9��^�n�wL�sH�s�d�_�?��>1��d)0p�+���[�٤��f�fx�I�n#�(�a8pB�q~S�	4�	I<��L���}m�s�>9��:fM_h�ءw	���m7x��ۯ�G�L&�s澣c�{)��ڏv0r`�!%��������R&�e��u���;q�'_Ѻ�pRg ��x��&��K˵���[�!]G��� b������΄�����N�0hR�U�ϵw�E�z=���&�İd��T��^�2���q<{�D�!���%(s����o8 �۱�P!&7<���|��L������=�9���I0Sm�\\��Y�k�m4�d�+:Wa�GV�z�����?���]�}�Lͽ��v�FNM�m��zٳ-?�[��͸�A�I<-3�	I���ӛ��"��$:��1�>'<��:<=6�WYȼ�?dy�םf�"�O�n���s��'}��~�iL�͙��p�)���Ȉz�!إQ�����x  �>>��)�ǵ���8篭��B]��1=���10pI47�x/`�8=��ܓ�<���L� ��{z��[�|\X�u�=�G ����vly&�N��^��of�iv6��s�y&�P*�z���d͋W���yO ��UQ����[ ���!&pA)3��� �s�:��#6T��_W&�9�\���ƴ%���'��:�8���BJy&�����_�v�p��9x��nΰ��\F����2��Ξ6{2om�z��0`�;D������8�>��|�޼}}7JI�L�q͹��4�A�m�Nj�2��Ȇ+n���A�NJ��.Fehw��/l���n��t�z	�:���>Tؼ��n ��S�ci�MN�PD�2�|E;m0pA
�\���2������=VR�70�O�|d���y�3п1��ٔ�=�9�V��7�-ȡ����f/8i�e7Ra���(�CVP�x|G�� [+���f��.�t����F�BJx�D8)3��pK[�ޅ�O��0M�89����׃5�������+�������a5X��8��d���rQ $�A	8	.�B�{yk��6��}�[�O�/+��x�<x�ky&�RN[ �3<(���S?�[���'����l�v���<Z�vx�gx8&D���39h�C1��?8%[ �܁ ��Γ�m�;p�
�r�`:!��]����ȸ��-5�Ӈ�{ I�����kk���Y�9������ǁ�r��t��C���y����
݁ ��VԳ�<��F^DF&�L$��z<AI������9oc]��_Rט�Ob�;w��S��5��O� ���p���nw�:��(Go@��/�`�R�\']�覷��o>�f}�9q�n㱰��<{���Z�<�P�w�}5����]�)f�S�ޝWι���i&qC�"*�[l:�u��a�F��{�|G��H��{�i��el�+��y�I<$��L��4۶Q��C6��^x5[�g*uw�1�������{݁ ���)8������ǃ��~G� vE��A�=a�(<;n�,k�����vx��fm��.~��������},p�$�<|R`��n����xT�VW'n-�ps9�0Ry��M��&x�;�&Q*��|�n���,g ��/��`֛��Ȅ����@$^3�Ƀ��*�B��#*�*�����b��>8��$��I���';9c:g��h�{J/�Ȟ�pA\��^�!&pAI����@W�ӃlK4z����R`��Zu���*VW'n�S��'#�^1���sq�}�a�ܷ��x��O�� �pm��&�D�qC�S�=��ح�j��^[�뀀Al��?��w�P����01�6������Z��8,�6���Bϩc,��f���x7���=���MO���$K���{o��G�%�se8(�}cY�{� I���.��"��{���h}����i Q�$y��u,3�1�|����7���?n�8��E]��3�׸o�'���C�LI�b���2\�6��h�pl�QN�p����G�ϴ�wn.
��]�Wm�h��8�����<��4��ĝ�Ǟ�e}���P!�=H���Ї���_vz �H�,Xx�����̶]\��6a´h�M�y9�;<��
��vש3�9�0y�(YB#Oe�cYC�g[
5�Q��uk6
�t�M���4������w��食��ʳ�@]z�c�E�H����B�uE�'`�H�I�\y��M�j��G������������D�kf��
z���{��4�C����-�5=5���g]�5ۓ�\{ro��Q��Ō��|=>�`úW����w����\��3.��a��<�eHS�A��)���E�'F�>�Aȩƒ��
7����6����f1T�^;'�N�gi�u�&�|s���C���3��7���Nn�yoĸ������^��<3ɿ5� �ܷ#��!���O�nu�yD]S}3ݻ��x�ޤ������I��}�}]�����"i�&?_M>:=�M>�=z���Y����.�b7L����癈��r��]���U��Ke�F�)�U<b��Q�2x�� ��N�ı����5����y�|��F|~/���󚸔���]Y�%�#�����GW��>���E;��=�DbOnb"��"M��޻ǝ�h1�F����b�a3���r�cw��b���7}��۽N$ӺN��ǊNW}��4������9Τ9��\5wuݺ�r��>V�{��9�N���y|���r\�AuݹÜJ}7Q7�N.r�wJ(����&��˲���/�7��6I.w]�)�5�'�Ě_}u ����]�i�{xFC/���`��ٹ؀JL���f7��	d@��[���&�A����D��\� �I�g��&�f�F)�D&2E5&2L��� I H�!$�¥��/U�^���B�WA�@7��S��ɸݔeLYy�b8�gUql%+g�8Mӵ���mg����88�՛v�x���F�������\v���u�e�q��k����kk��l<�إm�1M�mǇ����A{D3�Nu���y�����ۉ���ہ�y�Ɣ:7�6�:�g�)���nD�/Vc�s���G��mXGa����4�¼k��hwb��<�T6��R㪷Ot�5�@�f|7.��:�W�+[�Q��T�6N��:2�ۭ��������e��� ��s��e��uݱ�u�L^�*\�,;�q�\��>7kH��U�6mtEq��� 8��s���p��V�1���������r���<A�nu���d���6�(��!���i����[��rD#���,z��y:grW�v|ux����s�n��d�m�]�옹=C�]"G)�G`�U�j/���q��૶��#nص��b9�ۛRw8ۦ'�v������Ŝ,s�u�;��I��49��S��)Y�Ӻ��ƽp�C�ͥ�.6���r����,��,>=b�D���w�O<񡨥�P��sg�n	�0���^3�ur����Fyľ�������)�m�n�9
�����q�	aVv�]��Wj�[Ou�w[6ϥ8��yݴ��=��q�z.�e+n��d�7)Ӂ��V�j���r���$�:�mdґ�N��'p�G;tV��\Gn�����J�x�f��y�q��t�n�X����3��8�6�Fv����+�d��P.{f�<��rO1v�1ԛ\��Q���O���<��b���۰�O1β�l�%&�^C>��حv��懬��x�����sZ}q͆{����K]��;[���y2�+u���ka�^�m�lf�(��h�M�2������u���&�1r�y���mܘ/kC�ۚ�Ib�Q̺��nc��۝�&yd�ě�Ǎ��=u����KqƊ�}64Y�MSM֮�:�ڦ����|;�`;��J �b�-5c*�$�P�ORs'7TIZl���6�����j]�4��7�y΢��ܖ��'��ݎ����ή|v:C�ݙ��v�>�X-vK����gٶ���<�;0�X���l����{X�J8��u��ۄ����']�2���q��Gmώ�f`��aU{	v�v�����{�n�u����Nn���q�G#�-�l�Ŭ��;n�m����s���ĥ�3杽v8�:�3������]�;N�n�����߀���'5��zJI񜩼;m�������������a�ٰ ��pAIÐ�����<��H��%��?R�\�����v;�J�;�Ԭ!S����
T�A����7�3�&���z1��u�����)(I�������n5�*�=Y�q$�l����ePt[�^���NJ��?�L�lRo8�9.�x�-�[�9����<A �OU����씨4�w�0�V�r2b%�JFfgm��a��N��@>!&�$��[L�QK��n!�F��l?T�°��rf�	R�<A�C�Rg�'7Z�>ė���Ckkٔ5q�j˰�ް�vy����n�]Vzi:f��z�!z���r�Q	���3}�ނ�>t�9[W`����TA�y kD��}rM�u0�s�#-?�oP)3�����7o�\�SEM2� �DB��q�V@g���Yl�}u�Si�̟�� ��]>ۊu�ո���y,Bو�y�r�Ov�M64g����#���}D�QP���f���[�y�s][�s�}�Й��������@)0��;ۼ'F	�B���a^ ���I@���F;[5�8:Wn�*��V���L��?����&��	3����(��	��ܶ#n�@=��O��tK`����%<����`����'tqۂ*NM�G��8	4��I�|���Ri� �>!��{����z5NX�9�Sp ���^��R`� ���&{���}���7}=s�H�i�^C�n�F�4Yv�R�鳭�ѷcG\խ.��;����q���.8��p���@%C݉�峵1�
і�����I�ip�]���Sa�8 �RW�B.�`AI�ɖ��Ík�gn��� �N���[N�'n)�輎�{�8���	&�՛���_���C��Rh �=�^�ȇ&pA$��`�|�69�sT�N
jP�gP��ljQ���aQ��<q�.>\���W�Vfn@�l#&���,����,��;
h��{�A}DI �@$P����y���J�{������z��9{E�'I8w�3ӓ��Zm�� ��pF�G��ɑ.�u_l�DP�j٣�[�AM� `�k.[��ȳ��������3�|��#�l��M7�x�p�9������0�d輇�h�������i�2!���;j��O~&H����0�=���M��mZ�pWX�����x��n�O;�W���Ǆƾx�x�$�>)'���}���YWpipT�FR�h�-�e�!S�,4_G�XP ���I8���Zn�r6�#�u�v�v�s�HV��ukqo��9�I����1k=s��+o9�`�!$�
LBN�ϳ�mg�Z0s���$-T�E�p�|j�9�����I�I��R{0��R���87����)'����ٽ79mvRॸA�`�>sW���#*�Q����m;x�r������@� .@����K�<P�ś��7	�/��hPO��~�q���t�}L= � � �#""*�~h}�v��7�������p�����Z���o� {�5�޼ݮc���Y���N]<0�
L�RIOߏ�o�M���c�Q��x�`�2[L�ݰ����E]�NA��lG; ��������,}ݐ ���
N���XNc+x�K��y��m��1�o�X� ����������x �U�CJ��9�qk�泀A<��ELd�.ދ�7vRЌ��Z��>���=]�[Pg�4��`B)����O��.A�N���dFTOP6�tX���U�^�SVv3J_�A�C��9��E8ase���bv�CU���)8pon��3�3Q�Gx
.EL	��u������x�m!�)7��$�E$��$>���[[40񸗁�3��++�\a���_�zu��E�9�!k���6�Z�=��u�&�0��@䖔�`A�r����s�M�|	zs���ﯧ��XN�d�i�)�%��[L��(
��fZ�Ҟ��H(H���#Z�V�ت�lkh�6ۻ�_'~w��p�>e�M����磦..��yڹ��lq�i튮��	r�h���E��L�d�J��r��-��j|�P�+@�!��u�:GG�.!k[\�l�/k���5��n��ѳrѸ���$;m�Rp�J���|u��^�O���'q���k^2�Ȫ�v�ܸ�*��Vz���7p�; ��E�^�os�N��w.�[|��~��N6��p'\�{�`�탞�x1�=s=�0�������w��>�^���9$��ȇ�Ȏ�k�<*dɫ;��������c�m��sH �RO"���	�w��uQ3��4G�>�a>5�vq���(i��q�p�|Q��N���Fw�����h �����C���RO�-b���Ld<�r���.�R����ΰ́|� �P-�o]9G�x��E,�)�������.��4�c7@1x�i���r�>�� M��ׂO��L��@(���6�f�cd>��p�n�ζ4N�l�1ӎ.A��!$�E�g��v����_�K�xrC���X���b�]$��#�\�it����=�i+��q|w�������������A�I��m�q�aJЋ�	G���>)����T8��IÂN Qp|+.[f{�jmp�ۋ˕V���'24r)�2],7S�c�d�޵$u[�p��A��xvj\1o�j�a˛�&&�`l� �9�{�=�h��kZ5lj��d��-X�l[h�%[��E��RkX�5m�cY$$@5�w�y�Lߖٜ���[׃�U5����oq�O ���8)1շ����BL�<4��{q��
J�85�[�8hup�ӵ}OZu�gr�ƴ�sޏ+`��ÂQ>I��&r�V>����]x�M���g��L�C�۸��6�����f�`�-��wN�'x���ݬ(����P#�>)0pAIÐ����FEF������ƥ���f�����L��'�s��I������\I�$�?��°bM��p0�L�i��lfۧ��,�3�n�Ey]v솻pl��|~?'1��B�&I��.󙺦��N�������¼A��RO��I��RO釤b��װM�4��"�#;*�CFPT�c��ְr�
L�%�<�9
��� �'�Q����ƋxX������F�� R�D���h�m�p�R9�����}X�������|�g:���B��pq�g|o[�a�5g�Pd	"�b�k�+j6�Fք I�TI���9�;��'Ul�c93|A��ǀA�pi�x!&pG1u�&�0r7u�x�0pA�N����/S=j;$���<��/g�jh���$O(������A9��A�8)3�N����Ͳ`tw ��������Oz8��K�;p�k?���<R`��q�9v��@���5�㠗-���8��W��7��^&����Wa�&�P�����}�v���uÂQ>I������7s��M�)����#��c���ٍx ���pwY�%$�'��L=�X9�,n�k����A�p��o�:��y7fI�1W�c��0��m.�2"q���{&�� �n���?���>)'�Z���5�Q�Oy�h��+�;p �e0p8� R`'�P l<wc�4�D.fA�p�u��$�__Y��zj��Fv3q��8�����a�q0n46e��x�l�h��vۓHde���������6)ްT���l�GZq����v�JE�P�o�lD#��{�� � H*��o��U�����$��g$BJ�}]�����4��������MαڛF+Ja�b`�!%��ƠY����~�X|P�~�F�1�]��5c��k�r���uQ��:em�1�Hx� ���?����L`�/��3�BI���'kb��ӕ���Ev�g5� �(9�0	0�I@�|R`����l㽜�s����ݨ�-o8������:���=Fv3��#���)4]�&�6�W/N��^��A:�9$�G�I��BL*���im*��,����/���$��5��'BJ#�'�y�C���K�(>�K�1����N�S*z�3�";'�����`������>���i0pA�NJ� ��9'Iw��&�*�Om�3���^�kj�n�mW�����u��v?��� ���6������2��L��w�^�V@O���3�A�[��q3��M.��_+�=Dʿ���c�gz��e��ĒI����ﻗ[�ЧnU�p'�P_PA$@��WC&���VU�>�!��4u��i��>2׋⍙z<3X���N�3ڭ��.��:���9��{��J�����c��v�gv���ۍk4ZK�����<�u���W=[i����V�^�0�^��4n�Nzۊ:��x93<���:¹.̙�$����v��2W]p���;e��CF(���%j�9�k�䆜Qk����̼Wl�mm���;�?܌vK�g�׵5�.�@��3��F�x���/��A���|���}�#�&)8s{�{�;ғ�:�hm	.�6n��Fds]NnЏ$�$�A6�ǈ��U,Y��b�xl���x�mM)�zΰ\�N���ӌ��q ��^�2��86�ÀDe��N�I�����	?���ضs��J�cE�\^v3p ��� ����)3��I�f4�l*�۔I�{\�#��(���w.]ܕG<��;�Iw���5��L�ɨ�?����A�)TAA� �����Zw�}��[�fU��En�vQώ�����8��"�`AI��
N5
ǭ���~��j7�Ǽ, �����zv�L���]E���#Ֆ���C݌f��1h.�h�����`g8pBI�'��W͜b3��
��9����.`���ڵ� v����&r)'�oY���>ݷ��w,Q�N!5@���>��_��d�D_�~RA�׹����3o!ܝ��u��=-u��6O}�Z��q|�\�	�(��	 �=�< i��&
����e�ur��y��w�iw��l�����w˙������� �k�!�:>I��RO6^�'�ro��7*j-w[90��u�f�(��� ��zB[�S�]\�9T�q�������ȇ�+�9�!�y����v���f<��E�g*s8�3l��^<�p���!$�
(����Q�5���:��+���˖l��O=�F3��V�.#�!%<S"*�U��z����Kk�fr��#��&���z�x�vi��V�
��6\��rs�/߿��A+)��k)3�$��e��S��WNFG{[����9��3ِ�9� A��I	'&��`�i�.��/[O�:�>*�3����u������6�C��Ο��L�h��x �l�!7�-�u֞�S�u�&6�n<9�����3�X�\��J��A��qR�wɜ;�N��K6h��y������S9�o��2�$[�B9~��QV;���\�7����-Z�z-g{�.��:��<\A71�G���}��WkQCs�!̦nE�}p�=��;H������wЉq�?B��x�Eᳳf5"��t�s�{�th�����U`k�{Dl���\B/g�A�_��$���ǞN�[EE���'��}Ė,wL�u	I�q����NR���G�h��wH}2���6*l����	ڶ�w`��D0#`������������Qح�<���PB�
���w M�n_]Z����S�g�G������.3��+���.�I����?_r�Jv?ߨn.�l��h��I�i�h<Z�3���R��8ǎ�������iѽ�F��/��o�Ճ��_{�9.*j���nÞh�II�zj^��ɶr�^�=g����B��|��&�a��V�H0��NS<�/�dr�Ȕ�pa��f{����'������
>����8Ş]l�=�X���H^��7�T���Fp��o�>ٮ�:������{Ԍ�}��s�]���ݝ/7�]�4�?{���k��A����{Z��Y���{q��L�m�d�eܾ��O'�����[�s�X��a	�{��1��t���Ay��^}�3��>��^�\j�_�*�c^�!�r�㇒%�f�վ�G}~:���Nr��Osw.�[�ڶ���n�%�~���r���Ȳ2�,������tG��{<��w�;*�3��듨N�.�&K�����:�Ȱ��(&	�"e)G:o��$����"�e����"#	���D��zw�"d1��v�&&�~<H�޺�LK��(�zW	d�4�:K�;I���#��>z��#��n��s�:��#��&!���0gwC�v�3Ri+�I���3z�d����X�#f�\h7��JDf(1}�/]wws�(1�e�F���B�̟r4�M���ݙ��#/�lf)��D&��ٓ}v��+���b"(��"���*��M^"/����d��ȣ>�q`�O���xxx��܍����v���-[�?�BNJ�Ȣ�I��5�ф�����A�C�L�RN�YQ��,hQәQ�Ks��dKp�vS���
[Dx������P �.A	8	-�ӗ��1F���d8����C���sY9ɛ�A�0k��L�>V������43�����p�_O��-�u��ϑĠ��s��*q�ks���xq�Y�.�q����߽��}�o��8����
(�$��wr�Ω������M�ius��Q�N"%����#�2!�M��I?�f�9�|��h|�4�3�nc�mWQ���ٵS�-����k�0a�� ��\���ۼ��:`�u�(��)8pBI�2"biM��t��\C�`�&�3�7��x�Y�&r�RO �vgo����	�������O�wrm승�=g��6��c9�-G+�ց��a�=V]C�&<�헸gx��zq/��͚����,�S0MS�虾vn(����c1��i�[��	��l=�3��Lʗ����<=��@ }]�!������:�']un��)5[�i�]l��@��暜��t۾�0����u����݁$�t�voj�[\�����@.�!� 3�0��3�{Z�kEώw ���C�����lڪuo��������㏯����7��I~�ncq9�7���.��u��V<�t;�|w�9I���RN�"��`�y����mw�(�l�r;X9��G[��xWY���M��|h�i��A�zT���K-�}ǈӶ�}K�#�N��k�]8wi[/ԃr3	V��N��K��(Qr��I@��7���B[i��P�F�	��z�<BdC��j��������L������e�1��c�����ou����LI��%��c7��a0͡{%Ù�Zq����p�1�Vt.A�N���	��ϥ(s�NϒYs��3��ͼ��#R���ʄKY��d�b��^~��8�kC9h��
���w�Ǫ����D�`��}~_��ww{�����N��_
�:<Ý�2�OGs��E�� ۊ��;A�|̉�%�Osv��gu�M�]k �[�og��5ֆ��At��<���.L��avG�z�m�6�OZ�Å��n�M����6��'�WOG\L���:b�j_7b�uA�D�iۈ��m��̞twD�:����<�ݫm�n�C3�nϫ��(��mm���__ms�=�¤�����Z"*�y�9�7i��s��+���GP	|w���q�����#_�y3O��Ok꽙y��,�B��[�:���v~�otT� ���.I��P#� ���>�H"QgO�P!]G�x�l!��������c�&nڱ���!�Rh���[�G�/��O �<C����RP ���BN��6Յ5�
<Ӝ:�`��/� �h�Rp�����dC���E�jM������ZE6f�����6�e���e=gA;��3��V�������ٯ"7�h��k�$�_�$��IkS���n�^<�CΥ������c�[7�X�:ȇ)3��I�)e���
��8�ҹa!�t���(ƷO���ͷY�i���N4s�f0�� ��Ɔ(�⭃�s� QE� ��8��7I����e��_@���N.�q�`�"1�[��	�I���'��R�c(�}��a�5I��Âf�2cO��	c�����Q�^2.$4��n�ԁ>z!���o���N���^�
���}��������z��8`�@����z��>3�9���=�gώ��WY�N��8��7�
(������x)��X�p�V��J:\��8!%�Ȉh���n����q���r�93 8�x��9I�$��N7��޲�G�f� �\z̟]�q}�K��0�D>���@$Q`Fz�2�w(�@�ˏ �`��>)'�)0r�K�2m�۔4��:;d���V�WQ��8&�k`���8�F��/٫s�%��ȶ�6��qF	��wn�z�7B��0r��wv�Y��=7�����I! $�����;������L��7m�ҫ���&���%$������0� �+��:.X��+Y�#S�������,�!߽*��	����8!$�jČ�P���7��v�8=l� ������I�JI�l�g冩l�-Ew;ETdKLfT�������!Mn�������޾
�~�J=$��MECȫ��(�FT�cmfϵ��B+%�  <>{�ڟ�$�Iھ�a)�w�0��`�����?�I����@�zZ9;��'�D�Q�Nvף��=�v��MM�3Y����ǁo��EcSl0b�;��&fa7��\��	3�⒁ �MOKXC����,�OU�#�[:5���#}I?��� �'�P#�&G:��M����[00���M�>I��Дm���sūv�R�(^��wnŜv��v�/����{~c��0ӤG�c?� �c�d�'f�=q{�~0���O������(�r`�ZP �>h�]��F=��]��8E�fq�OQ��v�+53w�&�?��
M˃
%EP��x�uؒu0pAI@�QE�AI��Oۏ].��a�1�4�>�-p�l� ���BJx�ȇ)3�������h����#�Rg �
I�u3c��F)��х��x��|i�Z���P��3�S;�l3B�D�V��	J�lD�3���v��
r�+�A�l1|�~y8��7~����;�_"3c}��e��*/e�-�o�����z��o�I��.A�N��MT�<}2m��;��C��wn�1�~.��g&nX�A�6���������~���?����s�u��qϯ	�:�i�Y����nE�Z��O�k,��{4[���`�=�?�p�|���[�&:�_�C�M�0�I�^>�K`�!2!�Rg ���&k>�LSխDYT� �ǁ�����Ъ^ۇf��%� ����mJ�_
�F���A��� $��!%�:*d\��Dq�v�=iݺ��v�Yɛ� �ǂ�poH$�I��W:�1���ȶA�_@����$��qn����ތ/޻�
L�U�	|��F+�"����$�������>Ժ\����>�>=���f�)�5���c �� )0pAI�Hl����d�*�U��R��U�g�.Z�\<�#F�\V�cc\F�EJ�o=�t)�������(8w:��w�m[lrǱD7~������ߺK��p����{ݷ9>��籭D�fy�ՎB1#ۢ}tk�q[<ҵ�T�w!�ۺ�6��(2�h �/V���>ҝ�)[v�ha7O,���Z�P�7�-9�;���v�3�Z��ζj.ݎ�Tmcێ[;�L]#��P�A����lA6��E�ؠ�{tn��W�D5�㫝u��f�mڃ�Zw������������)ͭ��__������!l���<�nes�.!�{T��i���,]hl����������Z�ȴ��7��b]���z�wY�7�r�����u?����A$�I�$���N=NdTՋ5�����+�覎���1ޫ�6�,x����qk䓌ߖN_,J�`�V�I���&s䓭/�J�:�H�*ojYS[`�q��c �٘�<R`�f8��g�'�[�s� �x������Z��ny����=�qM�@9��F�-fmd�[�)��ps�>��BM���8IG�0�����0ww.֊~��\^LGz�x@ �`�N��G�I�ܕl��:�*Bj�݉.�I!ػ�µ����+���֒���g�x	�����_���{~|؂/���8>I<���-�/��T۷��gk���"�ۊ�!&7��fLG�c��σ�u�TvMC�Ax �C�Ng��[m�Q��8D�CC���������:��5��b���I�y����f�L��[$9�<� 2)�0 =-��{o�1����|���5Ã���rf�+. �B��Rn���I���NL���A=���@����}��ϵ����z�.�q�ޥ��A��G�o9I�0ws;3^o)E���8 ���c6��`O}s*-ۆ�f�A;��fd���f��mf���� ��8>��NWP���;-��e��ժ�k<�o��5������k��L��
I�R��L�cGC��>�)����?L��vof�`ݱ��)���X�R�j
y��i��n���<A�{�~�����>�$�8�Ŝz�z�k8���^���,9����K=ed�XG�>�q�<|nlǈX�p��J��E���*נ���u�����-��g�UÞ7A�`��AI�t�ٙ����96�<�!&BJy&����9�P�$����Pw���O��g햓�/�m������%!�?���Vo�
z!Wv�2��=�C9ːs��?�S��6^'oC=�⿔7� �yO �7�Ro8)'�BL�!b�z�&p�fa�|1l��t�8���Ω��W��ޭ]� ����fJ��Z+�%�#�^�	0i��O� ��U-#mQ�UU�q��[��Ly��WE'sÁ4Cxsn0�Y<l��')��%5�m�Q.��i�j�m\8U�2g��ZN��u:W��ڣ.\]��f��N�@�Q���%Q��ȋ]�z#�'9�|�{	��w�^�F��M.��Y��g� �������GC�ʧw�6_�z��o7gUt�y�x��^��M.A�O�8!$�n�]DU�i�Pz9����|�)?��g ����^�^z�5t�69�8V��>��� ����
L���@�ӕV��lad��P��Ů�[�'y����R���f8�
��gCz��ڟ`���7��rc�%h���9O.��3Uo���֢�xr2NMO��f��]E���3�9�.L)��W��/�|c9�;^<BL�����JL&��GI9L���׿�]s���4t���G�0�H!$�I�hedsYM^TK�����ձע瞵�n�f��zqn�iQ��qv��%Æ"����=<����$��	I<�h�A�=�:�7��tsh�y�r��2�ю/��`� �'BI��:�x[A���7����y�fb};ȴ�de��A3;����v��ng�8Y�ׂ��H ��AI���i�����uQВ�|F�/�R�����޽] �I��m8pIDx�'���$�����ݵ��*8u���x籸��矶Ӈ����A�`��w]Kq��Ӵmb�цi��B�BJ#�0pBL��_Z��+�:YM
��p�?�w�,c�S�ŵdb�-��c1���)7��$��=�/?������Ut]�O�n+�;�Y����=7����5i�������i0fy��w��v{����y딼א��;v��|5�D@|�y�Y?{�w4��ͧEs��׽���>��K����|�Ӿ�������I�U������:]Sl��ak���Orio.���yS`]��}zP��{��۫�'e�md`Ī��u�׍�I]��#��+���de��y��\����AP0_-W�m�g�B��*X�Wn�%�ț(L��t�w�8�tj	�{����˾;o!7OÁ��ԏ�{�����|��󔮫Î猡y��v8Dx	͸��C��};n+�3����j��g���	{�ȇ	�2!���t]d���FQ��]���>�{b�W�8�;�o{�4l�o���s�O��w��ز�X�m�b�ooķ��.l�~A�����n�M��t�������8�ŋ`��s��{�#����.��!��o��ʎ;��Ҧ���y��MP�~��C�a�����[��$&q��ݫ==;ōXj��=ۚV���E��4����0�K�%�������&�*x�791D��i���s�/�@ �վ��ܞ�lޘݕ�z'*�����ũ�n�&��?"o��}b;^�
��'|!�k��%�0H���^~�e	O7ZqţA��֕s�1��O1m?�>���^źO�a�9�J.�穮��1�����/��F}ѓ��7��`!G�o��;��=�"яU~<��gd�k����5Y��]q|�͜o�hF�<G����A��c���53�E��e�,�?���\�t>� 8;�:��
HdA��d��7�y��2�0>��︔%@����j��m��4���h���	O���6+��H�0��E��E���<��x��/ۺjH�$��b�WG���P��b�2c��-A�(�jL�/�x��I	���(�d�GuѨ�!F�j-3D���tb���/���fS��!&�xۑ~�m%�|\W��)%�)~uy�SMA�������x�����w�_z�� lbW�r��ѸY�U;u�W.r����O;��qŎ�,]ы2/QΟ8M���݉�-g�����j6�� �;]��+7�y$긱�7;n��yg�b+9�g���Ƌ�.8��8�ς{�qC^]��ۦS�n����g1qE�ܔ�=��X���E�΂J睶!��y��[B%��v�Bs�8�8&������9��\N�]�s��yu��y�vY���^�vPͮj��uԴ��Y�q�����p7Wl�I�FSЖ���s�E�-�0��U��;=u*��vy�kD���q]�nLx�㨀icvQ�^��BÄ������#�:z^��=[�u���G=�aؤ9f9;==��0�vL�E�\3�k/]�]�rҵ�9i6������.�����<u�v������ �v6��4nn7>�'�W���w9k��$�<k�x969�>�x��p2�5X�`�8z6Mͩ{�qFb1�cky��](�������J�m�ݪ<z��ݺ�����������G�sV�h!�r7D�K�Z��ݶ4��s��t����dZH�^���jE㮓�.�U۞�wf�\g�j��"Y��t��j�{up������c�[W!Ś�k���Lo\����x�F��;7k�-[�}��H)=z.�`�ݰ�t&�'#��}Յ�Ҽ���"vs���*;��qp�&�3���:�;/��۲v(���v��I��ݜ�LF�A�C��eV�#j�rGO5ru���.Gqcn'�O�nqcs��#^��N���i�..8�q��v�{&��Gm1�5��؍�evz�۷d*���][����3ۧQƐF��]�'�<]��s����ڮ��l�P�>7du����pj� �;�-�-0���5��]��d(�*ZC��{D�Ps�:,��zq��G]�ql��j�u�َok�"�5n�dG���8zM���W���k�2���o���-b�UZ�UUUU0~��u���Ȗ`_\9L���k����8'��#���;�v�*;���F�!0"��	Ӽ/��@iݸ�{r�����9{v����;]�^���(������ɮ|C�87Kl�g�؈���]��gU�L�ۓ	��ٞ�]箇�`�CV1��N��Mg�T���F0C
�l�lu�bṓV���9Վ�SU��\�3W�]�1�[����{���T�[V��x⥸؝�n�^�;�{n����?��L���dy&�Nwg���J��:z�p���1�]L���hG�o9I�@)'�Oœ�;�9�f�{���1��?������P ��z���K��>�{Pq��A	8Q)?��y���D`��۬o2�<�e�.T���,x �9I��RO$��#C8���+��L4�� �#�8|�:��o�����@�|U�pzΐ��K�f�`�����y�L�$�x0`���I�&��m�J�۷��&�i��6���Y����1G�`)'��g/s��!?Ǜ����L��k�v����huqr��0s��E���v1��#:z)�-pO�'�X1W6��R��z�[I������u��t53O����� �RO��1�Nc�G���tsĖ��/s�.���m�U&>��_��;���ȱ��ּL���"��`m7����q�wYm8�賍E���26S�=W�z�����8�S�F�����}W� �6\BN�$��6��Q�	�o�}��r�g ��"��Rg �������d��t(x��a�:/Ä�#�� �b� ���BNJ�M�,}3�y��L�qkBXs��:��z�\���O�"�h+&��� �pA��O�U�&A�J�<��Zʺ�7,a��t�>f���Q�ެ]����	8	'�ȃ��y��n�i�ܰt\#6T�d�Q�;�(�Rh���-�f]��������c���[q
L�i<e	mؼ0y�Ӣ�8In's6!�cj�w��V��A[ӥ�)8y�`��(���W*"Жs���o�(�KE�ch��T�*r�Rn �T��[i�M������ٱ���0E��q��
J<�4!'�e��s\�C��:S֎K`�X h�,�C�N:���{u�l�c+qJ�v=ď}<=��3����+C��8���|��HC�PH�!e�81��<b���+y��F5��Z�G����9��P#�ɑ�M ����5۶�s7��� �Y���	I<m=�cs���8Ib8�G?ۋ2{޼�e���$�G�Eȴ��	+T�K���T5�������FieVNu�p �T��oX8&pA)'��n�5��5N���L��Bq��]Mkm�R�7e�2k�f��{m���"������o*`�@�g ��wa����/����w�k��$~S�e�1|��?���<#�L��r�x#^�^�h&���ʛ�wS��8�9��n�np|u0	�`	M���f�-�78Μ:�amN ��$��I?��&p�Z5�n�����}y�"���ہ��� ��Rg��<$�3�S��ܺ��sy�"
��#�9y'�����ss�M	�=�K���|:p�
#r]A��7��$���Zf,Ь�1ļ�H̙Fs�'`�vW/��o��gԼu蟤/����6c���I�⺑2,�o�����	!]Ǆx����o�f4Nf<|s8)2�O�*S��7����������;����0�Q�G�I���#E"�y*;��~���G�sv��]zי�ѻ���s�s�^y�d��-߆��B�7�W3����IG���8���n�:o�L��+o�G�g^  �s�9�g �i��N)0pD�����3Y։o3��{/ѝ�w$Ю�޻�X�"Ӏ�����;wW���A��&
M���J��Dl��K4��ޡ�l{m�\�����E�poPIÐ��@�9�y�w��GKIbp���=%&{�6�o�:�D��V7x��<��v�й�W�s8 �}� �'$���(BLˤ�+G�Fo8�R��}$M
�;��pA�\!�e�̲���41޺�ɲy�7UuL���;k���bT\�E��Ar��M����s���-c#��\	�nG=vq���,�F�}�8�终�������3��r;)#s��a�����wW�n��3�����g[�����U�Br�-�`����8��e�ݷZڹ����:R��]��M�Gn0^U�gK�O#���I��.1���ݚ�P$�ܺy����[�>����,�uƳ�:�lݬ�98�%���E�<cu����w#:&�ݵ�X�f�o���|F��9{5�͝T�whȕvmk�����جZ��<q��t�& �ІXu���u�ô]����������`�����ݳ�d��z��v�x��5o���u��A�\�o7�����8$]��r�ݹ�s0�9�s	ԛ����Wayŝx�}�A;l����3��M�a_5x��%�֬��)z�ˆe\&c��dU �6�s�\=n�n��Y��T�ȣ榢Ʃ�.��������A���M> �v��Uj�znZ�8$ʿ!3�pʪ��/�;g<PY�Yp]���lv�Ȼ@��D�w�����cn�'��N������A1����7l��l�fa6�i�����!�9sH�qع:�p�t�[�i�sW���\�zָk��z�?;�����0D-o]��n�罞-�u[w�9�N���j�_[0�F&�7�_��_J���`�&o�����z����TU1h�HeP�3-��؇&a�	�A�Js���H���I<��f�)"YC��3����~ '�#�n��'~l�T�nz�D�5���E�7�8#-��f��-�1�4�S���u��)0�g���p.�?���p岦9���<��n��Nfu�q�k9��s�r,ۆ�Rnխ��,o\9�e�>nձ�}=�	�K=u[w��Q�D�w"�8'vk����y�F2!��8 �ݷ�[Y�wn�WP|�t��`�޶�p��k�ᢋw����x�pl�p"�Ƴ�Dc�u�{v�{Hף4�_PZs�8�#�6;]���z�=\i}��#\�˴���2�L�Nܻx޶�.��Ct�j����gjn(�����H�]���U�̫8J2f���e	�]#|'��80���F[뭷�z{�޼��0r�졷M7�������+��v�sv�A�l	��eS9S!��4��҂˧a�e��3fT+�B�gx�������i��l/;t���A��f��^�3/#�8�=���> LK5�m�����7�3�X�`� �N���"�ÀEۇTa]��&�8��L(}��boHo��=�{�Ѵ�r39�ڛ�&5�[���N���gֲ�q̠�2�fe�9�vo���,��SvWtZ�0�|/�y�8 �A���n����ӝ��7��;�s1 �h�
<���&�n�y�.M�R��{��s�[���ۈ�_���X�A���v�A7l��n���ᶬ���� ۴O�`Ȯ+��x��㩀�`.����-l�ݻ�CrB����wot�m*�gv��Lk9m��`x�}��M��\�iC7�;����V�� ]��ѻqL��(����*e��^��
8}���v�?����H!���x|���s%�i����,Rg ʾ�i�׫73Å����0s�'g����YXY��av1Bk�5h��.��s̑nQ�r��T�Z�l-�����r�rK�YAжƷgǊ	�Rn$��Nw��;�K!:݆gBd�l!�`]�eJ{�h������C��ҽ�ڥVxUe�Z�>1�c	휂n��^�~;��������Y�s����7Mݼ{v����v�M������q����_W\�r��8���ݷ}*T�E��g85�1ϭB'"����A�Á,7#�[�gv��T^b�� ���a�s8R
����:h]���Kp;��-ow��;9����W�����Ê�a{	[����"���&���:m�O^;��}�w����\��Lk9�0sv�A7l�v��7l�>N�va�Z����v����㽷}*aL\��g8��T:�ɹ��5�s�pDc��A�`���oAI��
L��y.���gXWv�h��.�w��p@8��p�]����U%gtl0�,X������۽������7���n/!Q������s��J�^��ޢ����'/2�����2\����`	��D>�WSp�`�G9��0��:��i���f���{6o]�Ξ�}�p#�kӫ,���\�d�s`95H�u�9m��nI�p����ۗ"�:+F�э���� ㇳ����&��/ �4@��z��v�㑩����*..�fzc�hƇ���o�v�S���qQl�$��t\�Q�g19�w0��/v� 綳��CBUٵ�������ݻX���uvǄ7m��;nmv��m�M$MÀ��.�ǽ���/�x�?���˯�������gs[u]\��u�}��]P0�Ӫ�@�n3a�Hps��}v޳r��n�8#�&��5�[p@(��q4��ݵ}ja<����y�:l� �8vz9�p�ئ^��?�s?��&��"|n��ݶiG����!���9�v���(U���^��w�Y2d��9�.�g|L�xId���HN��wݖ�+!i׆�f���������kq�k8"2�6�m����}����+QV-8�i�2�X�Kk���Vۣ����rn���N�x_:����Uŝ�e�̦�e���v�߫��?��#��L���,�(6q��7f��͞yV)=���U�=�s�{<���������~}��]���n���J�»�\Л�G����-�ŏ=�S>�qFA]�r.��f˂<'W6Yw�+#�q��(��7#8[�ޭ�fѠe�2L��zc��Qb���7G��P�;",%b����j/U�1%�.�#�������M�>�>��m�j�W�e��&�1���M�9�g�\]*���5x�8�9���v�͛>{��<�[ͳuMU[<�Z���Fs�h�z�Ȼp�6�C���G��u�@�S5S�N뷑�$�2n��Q2�]6�\�-�	��ȫ�q�6��{q�&)z� ����m�6d�v�Ȼ� �F�5؞{�k6�tm_*ډ�"x,U}���cY�"�p�8>�ii�ed�3sU�Yy	g,Y��$�3������Cg^���#vy�Bs��vM��/k{o�|~|��s �\�Ȼg$������5Ry�}��q� �Sg�����n��n��&휄6�Q��&L��%s*�jܺ~�qb/�6����L�a���2�5�!��)0t��̲�f]�fQ��O/O.>:��5��lټɹ�F}Iw?�RA�?0���8���t�����K�`����v�{_j4�߽�Є)�3�o_zL�ٽfC���l�8Ӌ�������|��go8+7݉ �|�O�Iw��^75m^�X~�xJ�+�I�m\j����;/�ny�qŷ}2װs^�ٽL�u�N����f'�|ugd}�����u���9����^���ofw���Ã�� ԃػ+����������nv�������?Xs_ڈ[|�!�'��>ca��bՍ��޳B�yM>�\�s�1�R�w�2<�g�o�M^��طj�/Gh��og?_y���-�D6bt&-�fl`T�u0�٪���#�nA�G{^��{�uå��вr����t��/z�Q�{��}���Q��<Gσ[yV+
���鼧�
��<��-���vC�D��Μ�����I��}�Z�}|�-�`�%��"s\�z}��_���~��\�ݞ����{��c{�W��N�O�]���M�_��eOA1���٢o����n��WB��	���3�L!���?L'��K�t҄�qR�-,������۽:��ۏf��M��~��/)������Q���Yۗ=�k�b.�i�A9O��o��_�('�_�t�:����{�n��l��{ٮ����q�LCt��$��+�˚�]�]l����>��{Yjg���-�B| �hYι!"�vY����=�g��gOY�#չ�����t�o[^�I���-�3��h�'�<2��۵xb+��}���פTX�cP[|�Qc�wj4cG�WM�Ƌb�B�cE$�65~7귈��ۘԛso�x�m�ۢ��t�����I�2A��(�,�����I��5�ab���&��wj6�M�p�rۘ�F�L؍E=��/m�(���b}��ADDm�x׵�Ѫ1`�ɫ��ӕ�\�Ҥߊ����Ę�r��h�}جd������T�:Tg���Qoj�ǌj6�4lY�����	�^-ʍQX�5��ZQA 9���������*jw��b�؛�Mn�!	�t�W$̫!�-��<���q����p� �.�8��혞���tU�y��p�"��$���bw<g��|�_
h�-9���`��1I�ï4��]$a�cY�Bl��j�-6"��p�����8 �sfˑv��a=������믤�U�Vr��pn��=Z�r�:v�5R�Q�>)�kF(�K�;�~w\���~��uۇ��!�8������u�k�7�6�/�to��x�m��ud!3*�M�2�!�������ђ7X?��s�g��j�*߼���4p�ծ�ԍJۺ�d鉈9ށmd?��9�7����z��wN�g0I�kӷ�m����N$�$�y�)0pA���fH>�p#�ltFwA���<�u��
 �Jp.����k!�f�Z�a�h����v&�A1�=u�9�����vL٥��Q,����n��쳐 >�E����!��Ͻ5*�{=Waײ17�/���(���y�4��
���k7Y񾦴U��z�n{�!	���#�A�.�9�e�-��T���2�_�V��*���+y����~�� ���� ָr.�?������wr����^�
�����ݗ��\M���h�/9�@�퇳��smz�wot��z%�����Ռ�[i�gv�*Z�3�#�(Tv&�%�~�Xݽ2rY�Q�u<�er�#2ds�^sGT\���}��2��|�H~��|��5��Q̫]���5��)��7m�;�n��}�B<�x�S{u���y��͗]����;���:�R�3*�4��jO�}���G�G;��v�2�I�M�}�����[�A��;��n��T�lmk�LШ��,�#�S�����wC�2�%�@5��|�ˤ�2�32�!�,�gz����s<��[e�1�ƝzNe^n&�xƳ�(�n�� �v�XNW?[��V���,�]=�Z�X��v�zIӔ����1�Z-�%�?N�����4�tu�������{��ώ}�￾� ������t�=���p�a-Ǚ#x����ɫ��^�r[OWn�����v��:P$���N�����#�L�^E�ۋr��/9�5�!8��x�`}7Gd�l�s���K�E�paA<�ݱpO,�]v�ӓ\��e��i�ť���iF2�4gu��!28�ۘ�G2k����h}^]7Y���q\�����師�}�}~_�u��yn&���v1-Y�h�tl�ě��1�A���U�^ݿ��G���{� ٲ������n1��)皓��{�-���7�ӓ�x� ݸr;]�f�sv�]���m�[F��u��d�k��:f��e�	-��L��Â=fͮ&^_;ﳐ֬�o�l�ɒ�L��ӑ�BdD�8hg6Kۋ��q��ƥy�7�Ʒ�Sin��A�,۰��|��l��w�l�S�<t� ����:���D�t�I�Ϭ88}WSto7M����Sa�y��p�2�2d,����ֵ�mQ5�oZ�ﶛ*(�D͉��b4Ir8ް�I�e�7n�Y���>��?��k�^$�we��n�����O�r�����y�Θ���|~��c��;�����?����N��ﯯ��$��J�v�{sw2��!��9�휋6��`�ßQ�F��L��&��;�Fq����8�LU�b�K��N��-A�.j/�k��DViS{zm>r��H�ٛ��8��آ����ŜB�м��xN�>:~.!|�O�ok�x��������>��+�A�p�]Ć�d,^���3��w�[I2�&eXB2��������k�Q�7&s-�����A��Ȼo]��E۸��ˑ �-�Ƈ`fm�9�����`��Vs5��}j�R��L �ޗ�Mbu�+��T�>>�P�Ջ ��+V,i���:?����L�0�ˇ5z�Dv�Q����p|h�}���"���[Y�g�J/��}�?WϷ�W����:�?퍫n�q��+u5E��J6L��N��ۦ����`{<�����߅�A=��ݳ��n�þ�^Êޛx�=���fNp���xU���O�8r+��l�awp.��;���
St\h��w��*�Lx�;���}p���άn �y�|o[�mqI�����-Z���۸'5���p.�@ ���-tc�k�R!?6J�U�T�D��ʑ�qL�a��wl^�ұ�^S�^��r��<����o�b��s�t:-�m���͂�����?T=��|��)D���σ��g&�e73(�����6\��7��V����g�l���|�+zZ�L�[w�pp|oX?��}����ntQ���L�|��"탛6\}v�]ي+,��[�D8�{1���_y�M�1��M�8��Zl��aл�w��K8�<�k��V��sn.;W�e,v.���u��u~zM�`|rX�$ٲ<�v��m�ckl��i�Ϝ�"S��>��,s�N���k!��g���S�eT�'�ݲ0�3��L���|\�t��i�������A��Ǎ�3b-n肆c�pFk������X2U��-8γ�t��\���桗�e+,����x�M�9ݳ��y(�k��hn��A��kz텈��ͳ]�W:��d0��� �:�3�:S
@�RHu1hk�aF`���P7�^~<�LJv�ٻe	��UI����3G�۾��!>�������3�U��7m��z��e\s*�E�2�߬��Cu��gg����R����m�M�	�����I��N�Fz#le�q����sm�- ��GN���9����w<���曻�^��\�,<⬄7ՖC2�c.�8=��1����m� ��ND�1g_&�z��n�׃y(pAI��Q9�m�N�� ����:���MWs��qL��F�8z�]�Jz{�}�E�_
��B�d�噿a�`�2���&AN�>�Q�K�[V���&�e�`��8I����8��^x�:<�u��L��ݬ4�,���F��o��<�pȨ�l�{³:m�NK8>���uӻ�w�@�d�1� ��&�|� ���a�ms�1Xv;E��n��Uo=\F������`y0�Ð����q�ݣ�G�G�mO�&�nϧ��׊b��{׎��'�屢=�Ϩe�����|�rđ~Z�ڻB���z��
�����2��?����|.9��귮ۡ���[`�.w �G]z�Z�oc��e�j4�G6W�1��h
B�����/��J<��9��׬=C=���Z:x6�c��r/]Ӻ��!�n��1�'̈́:�����n�a��d���׮��큽O���	��Ԧ۵a^��`+�z����Kr A�l����أYh_,���~�W1��n�l�.��5W����<��n�m�
�^9��#�Le��٤��ƻ	�F�U(��RU_��������]G2�c�O�}��=z�f���)����
��_K�#��ss��Y˲L�.�N8�wH�כ�G]���C��ѷQ�3K�����rM�87mOY���㯅�pG}����.�9�e�>�prS����N�tj�Rx�)o���#m�����.�?��5�y��=�+wjo7���9��7l͓״ݬbj��{��8 �`�Sf#Y=&9`�+�� u��-�8 ��ۇ"�.k˓�4�l��⥃��r73O#�����g���p&��LdI��/�����4\��c�� ��c]y��mƽ��t�<��gwhf.�o��pN&�	]�����<dr|��=�)�%�l�>xu]�sϖC�h���m� u8$?�7l�r	�a��e���y��pͯ0��(
�`�E�o����Ͻ���T<0�8M�-FZ_g�HG=�U�0.\^[{���w��ی����Y����>��s;��[��p1UV�}�����L����m�/��)��va�H[vw�,�Ҏ�V�Y�XC2�c3(�f��b��Tnp���hг=7	���o]���n���[����"��.�G0L3�v�������g�wL��,�����pE�*��U7]�An���v��	�g �v��[kD�a�����9����+_A����X�����;n�]+�a�{Z9W����6f�#� �Ժ.��wjN.޺����n�C��nB�-8fۋ��5� ��r��c�w/�j�KRηm�4Ĩᘧj[�\a4���,��	\޼oO��g��ۇv��[Z��Y]h�։v����r9�2t7O*m��o�;�	79���e���7���k����q
Jk�g ��k!��8 ��f��ܭj�4��xW�r ���	�1r���b��&�^�n@�Oqs��;���1����*�f~+�xz�%�?iWٲo�Y��~�$�#Ϻ��iU�VF�4�5c|��o�!����Y�Z��,�w_���F1o X���w��y�뷙>��3\1(��	��C��&�3�^�Sg�}��E�8>�7l��n�oDbkn�Bo\8=L�t�Q�,�y������8�qp̦��u[�y.q�d�<�l`IK�����㞷Kd3�83�Vΰh
�Yӳl��i9��&؆��`;_��| �g ���7m��gȊ����b���f7��v��칮9�\ �Ֆ�{��2�a�e���Y����;�n"m��ޑ5����b�ˆ%���3������v0���]���-�3-̣�fQ��.˃/����|�����͝���`3H"���o��<L��ɕ���g�*���gv�2*k��8����ٍ��M����@��R["y�9z[)���$�@�^b�n#�ox����c��%9�ۛ�y��5�Gv1���z�����z�D'��l3(���\3(38�S�ƾ��@��2����a۰�Q�-��⥜��O�7l���pl����{c�,��y㠲���nF��E��w^����:�;1>g��#�SY�n8pn�9]�y�K[CW_W1�W�~q��Nk08�9��x����?�����m�A��8"'{n�sɢ[����gn��T�n�F�u4�;1�n ��"���ݰM�&E���w�Q��� �'Eۿ��!��-����[Z"�v��J;)��n ���n�Ϯ��l���O���_U��˸=��/�	������!'6��|tS�w[42��?�-���܉��A�y���sv�&�� ݿ�ݵM$��ĺK<������x���q��[|�M� �]���t�ӏ.=�_�Q�����]�g5����	���ӹ�pU���n�L��2��K͙��[	�y#s`�R��jT�����Q7r(K	4�9/'�\>u�!��7�K�e�wNތܣ:N�޼�g�w��F�j�O������wҔ������z%^�l��3�×4��y�	�;p�ؑc�$G咝B���� �å�f���,w��� Qw�4u0n��ͽ���Q�����s�&���_f�
Tck�]�����ٮ=�k��˵_1i���{vAyeD���c���k����n�$���� h��頳��,8L����h�����O4��^@.-�ly�|sw�����#����p�
���'���os���k���Olʶ�+���g/;o���yV��㑦ICU�0n����|�|�<�\����ڪ�E�{t�����b:4ckH��^.Ѿ�된��</�[�{���޼�r�n����0�)����O4i�b��Ӳ���ǆά{w�"�y�;����c|\(0���8(�����!
�s׵,��v%}�p����}�[Ǝ�|b�y�!�Þ��=��q:��}���#�������������7��N�I'����
/���d�y��]����g�T{;F!��R���d[�iA��K7�Y��}���-���xH�mm;������,��-�������M(�4-O��o�?./�=ϼ��>|iJ�)"^H�
-6W�z<��<��<�o7���a��EV�5��Dr��!�b��]�/g{~wc��� ��Z�j��qW��}�$^:V	.���\�.mE����5�}����Q�������m�Տnm��i��h����s%ʸY"�2Z����*�ox�k�X6�v����ۚ������j5��[�э|�,j�Q���5�6�nE���b",l$m�UͱzW�;Ź�b����F��*�%k�n[�|��E�a+�b���ٚ��kĕ����Z-\�k%Q��U�z^-��m\����s���r��^����P$C�wK�n����Z�z�Q�;S�GD��x�ݱ5d6]m�����agc�<�؊W�n��yyW�GWgg]\�����o9�FR �q��Q���g��c.�A��Ȩ��G]e��sq��5�^�M��βa�[\�n��W�t\n[��Tv��Qq�mK�8(��^n[��`IE��;;�t1�`EMt�՟]�yn�e��][�z,������Jq��gv롑�ڷl����k��8�rs��R;���κ�u��-�g�*=��]-��f��<0V���ܟ�8舷d����S����j�:��ϥ��s��X��:��I��yV'�9ݺ�e�\�nOJFq���Z�kf�j���k1�qX���vl��v�抲��;�Xݞ�1��m����0��F�q���9�)v�a��S�\�r�E�3���Og�g��GvD㺮12��G�;ƺkp�1۱�0���]]�g�A��i�=kkL�n0T��Ae23P���=��ͥ��oB�8��q�[�N���#A��,c��t99��=EGG>.v�1s�勑�r<�ol��o�\h����*��m����OU!����ir�]\��\�uD/�#���lO�@��B�E�0���𺮶��5�T8�K��v����I�;B�[uť�*����z���9Lm�zC�^89�3����\��#��]��n�{1�m��mN՚Z^�Zܓ�t��"��i�
��s�j���m��_]]�!��3kn��A��S5���v^y�:�i�1��'`��O'<֮<�^�86&��W��j��烓�,�6"�@\��p:�ۡ	R�=�K��wV�%���cN�����v�cZ묎�v�;Nb����cf�C��@���Z�q�v>���m��6��B���Βt��B�m�-�v��P+��6�p5Ň-s����M�C�Ƹ)Hz��Z6���Qj�7�s�)��םY��f��.����Mj��Z����p?��������VZ\^t�v�[���61��&���{q�y���Dv"R�ۄ�8n���hp3��=9��IF;ӑ��Llh�-�KQWc���{l#�F�S%�թݒv����[p�7d�n�61.��Hnu���Y֎W��޵Í�s8X@#��vq�K�B&���uE�\��ǒ wS�չEٸg�k7���-�0=�ć5�m����?��5�c]���.ͧ��t$�.s�(�
����0����d����?,����,k�?����"��3C4�X�?N7�6հ�Q�K�ݸ��a	�����g�m��`��5�WS؍[l��r'Ex�F��8�lh��޲�ʻ�����!c"��K�';�T�<����v��>�o?���n�Ϯۯc���کg���i
�+1�nz�8Zo]��Eہw/�T`�|�3+H ��<G[y����9�)��Zy�:O�M�����<o�K����k��I�g��r.�� ݰpA�ۇ탧���,�a��<����eݔ���p3�����Eۀ��oF��$����)Aa�X��"�q����j����7������u�l{wdo������'��x�-�퀻h���Bx��ٓy�����ř1V��}��8����a$��\n�8><�Z�C��n�����w�qN���b������߫�E=F"2y���l->$o���}��3� ����2|#`�V�jZ�ꯇ�^;�����g��l���?'�I���|T��q?��ݶv�t�c�<z�W��al��0p7n�타An1L�	�F�V��WGrsm�O{�:���v��.���8t"�Lu�2 �/_���h�8���̓�ڸ�U������"[I��i�/(`�	0r��`�1�Z�������@��g3?@�� +�ϻ\���m�L��t��ہ������i �v͝L�}�_�־}4���a�9�4�֮3���{�]=;Ƕ��A����b]�C���A��]�x�����;�Z
��~%��F�z��9޻����՗�̶ٙV�v�ǆݣo��l�x��OVoZ��s<s*�^�f�|o�8 �Nݰ-�gMCi���8%&��9n��a�[�6�W
��8�$��`-��㣶5*BM��HՔw�;m��A�}w��zĄr�yY�j�l�Ј�Bj�R�L���C|a�zqDb����t��M��&pA���9��z�]}:��~�:݀�v?��I���0vj����-���2����Gf��n����,R��6��7��h��L�!&��6YL�6 �q}ם���x�]��� �|��>I�i���՞�{&�~�+��qo՜l3��ٮ6�'l����3W��:�lV��v11�[����h8 �pA�4 BU��M��Knsb5<J�P�O$�El�~��К�#���u�]��v�A7l�>�S�V(԰r����'U��q����e�p|r�8 ������.æ3���=��A9��9�g�ݲnY��-,�Qή:�̻Y|7	�`��-8sv�]��Eۻx�+�q��o�����t��F[y����U��kƧ�]�])�M�K8>}��������o��������&:njjm;����O1���e%g{}6�`U����[u��X�X��x�+�5��\U\A���?o��>�f��?|�BL�v��m�c�=3|����|C58p���	�ۮ���9}��r�IÑv�qV�|{�e�f���L^��$�;��x�=�67Zfm��7��V�v��n۪��i�x7��d�s9q��ݳ�}v�9���Y'�f+Y|1��m�C�!��#�/���ocάC-KN!����\t�BA���+_���=�k>�U׎�)�M�1����Kfֶ�v+��#6��'9E��e�3(3(����L5�ks�$�TEE�b�2a��0r	8r�j̴�ܖo���f�Go�|	c��si��n�w5Y�Q�zFb���Y���0r7;
��3�Th�i��@������p0Zq|0Z�`�|�ˊǡvI{�k���ok9�Y)��t�z�p	������8 ��gn_�Gt�=\��][F��"B�9IhK���{(g�Ko���y"zy�����oޏ���a��X��|�.�ñ�$z||��r¼�L�grF5H[m�������b�tj��Kp[8,m®�J{s��Y�C��c����5Vkm!��{t�o;��8]f��ڞv6�v��u�n��:v��Ϥ�!��= �*t�=oDk]��tW:�[��v�'s���C�g[���%Ԇ��y��ٻG�D+QM�787\5�.�m�9�s��\jU���;w��l�����?��n�8�ʯ	�^�Psn�Y�����K[vG6�/��|'[��T�pA��l��ҷaq���uVqw�s���\%s	�Lx������9�^T���1��b�=��3�A�g���R{'�L��kf�7�����`�iIu8��]�xf����7n�zE��z05vgQR�����]x��hJ-T�cq,��l�pn��A�f�0��=Sj/ ��Cwu�!c�Å�]�uu��7�B����ާ���\�\^�nj���(�ഡ�`�K�f�B�w}0��O�
�T�9r���tt���X�in�o�ybP�VU�z��C욾���N�?�h���uϮ�սVJ�uܮ�����r�r ���h����pN�>{��?���q7%�L���S=X��*z���11�=/u��O+�XL�[	3*�d�\̥�~n�#P%e�]U1#�4
����B���z��S�~�(����pO�A�|7%D{E�U�sq�u�{�{(�.��p������B/�%ޓG�9�/��_�<�\5�_z���d�p"���"�2qs_%/2P�u� 3qw�
�A�hł҇֗��a߁݅ݣT�o�t���X�ib8�`� �Ӈ6l��v�ȻwFsp}��b���Ƚo"�Cm6�͇놎˕
g�� �g �녑᪚�#��!&�W�efQp�e�2Y��Ҳ�@xq*��Rؖ�V��b�S�d�pA�p�]����ȇ�;&nd�Ls7��a�9��2�����!�n۝��
�e�`�C�:��	���n���5p��,&eY	3)�dWkoޙ�w���k?2��O7��E1��a�E��� ����r��g���������;xXu7�&�/[5f�B��z���Ӎ��T��E�!��n��"��BN�9u��ln��l�n�G��!�3flEĿ\�"�D�����7e�]��^��õEBd�M���^C�7b�`Ǖ����Fl)xyS
T�v%�����Lj�QW��K���&��Ӈ]���v������}�����r[�m ��H���ӽ1�V^.��{5�x�mp^F��O�sdތ"y����\.��A�p�"�'�ۇ:�w||y�?��$�z�G=ڋg���)o86��m$n�ncv�>���z�ۤ8wgZ꽢�au/�f4�#hװغx��ۮ;�7E��Gy;� �|��E�8�2��W^�{�)V%޸��oF��UT\�!�ޔ�A��&탃v�A�^��;�U6�
���!����uo)o�|�X8fz��z�㸸��0�y�&Q�CyE�󺰄�-�e��C�b��z��^��7��b1Z{g���	�(`�x���� ����y�~�J�f��9��w�O�GeUv�3s��fWz����L���y�n!�ʏ��M�A�{�+g_l�"��&&���8�!�,�4���'3݋����k-��ۯ���]��Yk��o뽮0�̩�z�y{q-�� 1�0�?V?�Į`�ݳ�A�g v޻l���阖��'š�@{�E�z�a�J]����;��]��A�ۃj�/,�}�2\U߿~z���Z��M�U�F�<��\L����Xͻ>g���kR�����f�e��|�~n�!ͻ�v���˛�D�.���N7���˓�������Zn�X���{�ᒾ"�f�����
Y��>:��T�O���{���D�yŧ�57ͅ���������ɽ��Nz�!fS�\̮2dQ�������T��V���=�%����0pA�p���rۇ]�p�O8eݝP�o��r�9�?�7lr;����b�OY����%��#��X�����ݽ���	�g"ͻ�`�n6^�y5�ڧ������/��|��=�IE�Ӈ]���k>�J�Z^��T&�qz�����fn���NPp\�R����m������\/;��w����.�6����z�a����������@�$���MǠ�؋�n^�ս`ݥ�sLh^����ڟ#c�s�i�;p��Wں�����N0���Lu��q�-�S��ԑx��r�9���s��݆(��z5�oH2n��F����1t��'9�^;[n]�Ə��W��N�#bfi<�ꃃ��k�T��nzՙ�]Wgr�"M�Y,d�V�,��q���+�l�m��}�1?�w0����v�âtn{d[��'$LZ�w��2O��~_~��,�q�����Dr����|g�᥸0|��C�7�8�	���⏮�In��l�r.��0�L��o�����{V�w-}�.Um�B6���cY�6���ti��e�S+�5��L��� ���(��]���kPꢔoM+e5|,c�Wz�h��8r�"��pn���������e���gx0lm>��p|�8��b���X�9o�p'y�+�99�L�jU����E�����]�pM�.A�p�]���dVui�!���b�զ��ڗ��d#o�A��g �-�n��}v�p�f�f��x���$8�0�1p�a�g1��ݫ���m�m]��{q��O]LV��}Ϸ�*X8��9�e���'��f7UGAV3+�s�����ؔ-���Lm�4&��Ć����V�bWUW2�"y�9ol�M��6.�|�cr����M����!~�>C���4l��� �0����wd�K׼��rWp5jc�
�ߒˆ1D��,�xDA7�?���ǵ��o�H�_w��QƼK������8sv�3�ߤa�w8pA�`]�r.��v�Xd�a���f�h���AR��{d#�7N���3���fU��fSu2ty��|�u�X�  ݸpαZ;�k�+��޹�L��F�g�s��x��3��k��>vރ��`.�drΆ��sʯ;�ǌ�=��9��Ď����\��9�~<Z�8 ݸ˘YpZ2�q�uϽ�?� 6cX�xl��� 6x޽&x��wN�g�+=I�66ҍ�����~��z㏟ۮ���E���.�븥s3�m	䛁���ʇ2V��4�
���p��&��]���1#�כ�J�I�q�Æ|���='��G#'�w���T��֜9o�����f�$l�Ŀ����o^e���l����8�����Ӽ�W���5q~�[>?.)�|��[�9{Q�嗦8���f��u;��7�M�?{{}Gk[�c���g��w<�N�Q��znW��ɛ~�VoO0�������b�8�ڱm����i�ǩO;���w1����v	��=����
���is6>3�ۢV9��� W��;��I=[��mQ�{��!9��M�Oy������>�n�t^��{�i�jQ1WXC�ќ�,(��8!h�*�]�m�{��~��c��[��o%���T�����C*5gwS)�
P�W׫����ylo׉��2R�	sg�K�T@�����
�<z~�܌C{8�_v��ݚ����`�Ӈ=c�>^��H��[s�(�[�״��n�CV,=ޚ��q;Ԩ9OlZN�Z���X��=���*y�����
@�9h�� w��-IS��K�=�p�o����1p'��|t�dΣ�W����7��<g���h���+����a����W��i��q�ׯ�;���B��7[��뱿��zy��ES�{�q�i}��4��@��;P{��C���왼W
�!Q��C�h���t�����>.���;Q^N=���{�'�o2��o���t=��7���
x8�Jx�����O���Ƽvl�:Ȱ�<�ղ�L�V�&�ON�%n��w
���*5j����/yŖGs�(	�ܙ���Y���Dc�f��m���N�D��>�|_x��Շ+Ѻ��n5��_o&�mr�]Ѳj0jHܽ��wϹȽ�Ǫ�=ܒ���X���r���� 30Km�냾9'UJ�
�@��"HSnj�wZ6��5\�r��Eʍc�[���ή��m�Eb�~��E��6�x�[~�|W65��-FѭF�}��o��m�h�r��Vܷ-���[���*wm�kr���|Uzk�=,�M�ks���nQr��Ilj�-sFɊ�Jܷ�^*�M�mrܷ-t�ܱ͢|V�m���Jޚ���^+żE'WI"*2#Pk�[�E���cX�9���5�g�ڷ+^*׍��5��#�Z�U�Ex�j�w�m���%Ī�ۉ賎:�o{�d���%��|�A�ݰl$����NM���L�VŰ�B��w�8Ś7�w����1�'�7	�g3���q]�R�/ǽ�i����v�A타Anݰ��#M��R������rxݞb�����U��)����w��z^Ϲ'���{s���q)rI�cH ��p���Og:��r�hN����,�'�w���?|q���E���n���<��;���TG9X�f���Sۓ���8�p�v���	;�I���XSy�����_?��i��֥�x��=���c>S�|?�[��S�Rh����+�����f��"�Ãv��"���\N:�(��YL�m�;�pL�A���o��87m�+kv	��ljk���A��v�����Ǔ<�Ĵk7A�oz��㛉=2[r���0��S��o1�хj@l��w�kw:i#�ӄ�l��U��f�,S*��ڊ1�G��g�O_.aK_��ջRy�5I�=��B�}��0r�p����v��7n�����g�F��p�?��op�����+�7��cz|n���v���/�c�=h���q��`��my��WF�9���)��t�K����ݛ�G��ue]5�]�3��,��E�&e��:��=�����S޻a��/�7X��wE���p�fe�LʲfU�����Q~@�3���g���ǻEy�5��n��0r`���5�_�BEg6�3yAfe�˶��}��gWZ
�u��%Z1��
�M��rY�AX��d�ϒo$�E�����`bi���\84�9�n�f�GOu2{V�*;�|���`�p�=&��k�n��m�W�wm�2�fe[LʸL�nfW�|�-���\�� �3�T�v�3]f�W����:��'��	�]��sн؊f�#����e�f�711��e�1��1�L��z�y����v-��WPB͞Kg�[ω;#����[�~o���NE_���b��zG��D�v��=¼lv���]sw@�'���N��:��ú�C��U۬��٧�Y+��ח�&��;d��s�.1�v8��T�^3V��"��{v�2m;�!�[`�낰�y�G\�}���׺w	F�qq�S6�>Hs��ٚ�6�@��ul��籆�8��yܛq�tN��-c��p�l�t�E�q닅������Ba۹vmm�}�}��������Bsk��ɬx�������t�!궳[; ���Ml�>�$�q,!���f]���Y��v��9|)��f
�M��w.ݰ��^�,�C�M��fϮ�I
7$�:ٯ�F���ృ�D����K2��!?z���h��6�9o3�d;�w�;�6}��}�޳dI�g�ݷc��	�k9��_�NYxӊ4�q�`�$�͛.A�p��C�¾�sN�'\8"���"��K��K�k�l�;��J��MQ!r~�n���0N+��QY��ӈe��g&�[�t�������w�j{��XK!?z�h� ����n���D�X�T���T�E�C��0	fh �U�L.�\s�b���G)�]���;#��`/����q��\��Hpn��&�{qM���U�E��dp'y����k��A�a� ���`�6_��!D�bR%O4}a��ZwzG��f��l�ZV*�ni��;��������u�4���8�.��P��d6�lYL���!���|�<������:Mgq�ye8�x�%[9�Z�;;�ޫXl�]\:�[Me7l$����讈��vSY�J+r�+X��pJ�I��.��n��n�ȸ��z��EF-��am��5���يP~�5Y�G<fG��>2�8s�g�a(�`a v�pA�`.�H"�d��oӰ���8�Rβ�,��op*���`.�H&�n�a�h�4����Y��)�KkY�mk�=��t��OEkw-�RI�����>�`��q�X-9�Վbn󢻢��%���T��*�v�euu�َ��`K������]���E��8ס�<��r	�g�)�o���Lb�	��})�t�8턽�=����pLˇ�}ݽ�!��a�c�s��9���=�������o���ʽ	-�A�>#/��;3��J���,��^修oz��߷B���s�}����{ڬ�JN%�__V������N�J;z���J�뾫�$�*�G��fU��̧2�.��;�Zr66�
��ÃX��"��OW�b����1`��)�����)���w[��5n��O2�!	�VRQY�r�Fݻr�ZL1����I��9�vM�{��F�f�x�`���87l�wJ�"Wῢ��8\/Ŗ�@��,m�,��p�#<[�f�s0,���q���&�dQ��ϖ_�ӟ[}�{z����5��6��Nl�e�D[�O1����7��Ǯ�0_-��/i���{P�{�]�,k`��]�و��Ŷ�y�zM���}wn.��|���-�XƦ	�jO1�r#m0��O���J`?[W֛Ne���;���&��{���?�?[n��ݶ��2g�7�7y�Rf� u��th�?k[/]������y5�Ncɋɱ��w����2�An'Ov�o�w��D��k�{���]A�yWd����ݸ�a����#�8%����٨�c�R���׆5�����쿯.�]�"љ~�Y���s7
#��,�5�l�ݞ&�O8-�n1Դ�l{@1�b�f����m�܇�\��,�]��7�WxWj�#D^/��)�^���z�,��]��73_'l����X�{R���Xio�%�.������Ѝ<lO�u�I�v�����R�A�@2+b&�.Ƶ؝�bX�epڗ��v���]����6�S/l�mv���_DFYF�%,���o�n�Lc�b;��)̴�m߭��[�Ǻj�VAz�L�K�a��S.�o���5Y�fʫ{�mf2�"%��ݞ#��j5���/� ��t�HaDS�^�5-|YE���Q�f�����w��C�Z[��g�^X�x�������cj�$*zt֎'5	T.�]\�ف���K��m�]q<Gcr�=��r����z�z�13����{[�k�1W>xu��&H{n���礪(�x�.��N��S�.9M��i+���9붝����x��Z*�j����Kml�5�[�-q����>�>�6<��ͣ^q]Z7	����C�F�k��m���F���A��O��n1��x��y����]��w��Ӻ�����1`٫CڱϷ���ϊ7f;Q�8���vȁ�=i���v�크�
�wQ���3�x��1f4��H	��wov�l{�7���l�젩�x��ظn�}�l�Jq�Ҙ���g�����Q���En?������V�Ύ�&m�r�lf&X���H��M�]����[�]�^s��a�u�������H��̌���/;^����nM9���O�i�-��o�o~�
�_���y�C(��ٖ��fS����Lݿ��:�Gv�������b�!�h��&�i��%Ȝ#7�0�� �i��-�p�k[q��?���.=��=m��I@�̽�̹��5С墟K5n�=Lމږ`uj�.���v��>t�a�l�ZGUcJ>|�I��$�բ�?�!}�=��p��`ڷ��{Lؓ��gn���9i��z\�l^�<k���c�����5'6c�n�}o�������g����'�y��8�.�I����wjη	7�\�����ܳ<F���Ҧ1dl�Mw�)�WxRd��@���H�,�����l]��,{�s[\˚�8��tE��ѵ+q�{������`.���qPnh�yD���y�\S�]����qZ޻`.�x�gc�{���~~�~�v,q���]:F�	��p���$��W���I2I���"Z��������߭8�\l+��3Mw)�WB����<hW�M�wq�wnW�Y�nc���í���j���l�#ׅ�P���.ǻ���0LGݹx�}�㖜������}�F��/�
��_g�hΓ�^���D�R��i gn�޻48���ٮ�,~���7��x�o���Q]��ܘ�([����^�5C�\�x�L�5w���R�^�~i�.�����
�m�{�����pm۳��y ]�h��Wӂf��:S��q��l�˿�~n�����m������"�chwEn��׳ؘ��W�����8�av�4���5���c��bA�D1F6ǒԽk���t;%x�l����mZ6m�?���oL�JoSj����t���Vv�Y3\�R��l�D�[x]ۋ��jmբro3�mg���L�jyWՂ��.6Sq�z��s0�k����j��M�.����]��wo2�ֺ��;]:��Yr���15B�}�L;2�E�
�{�(�L^��eZө�v�1EG7p�"�-%9��:,��XA�iS>�y��W�*$5TPs���3�{l�d���	.SV�:x<�kNo\_z?M3�m�p����t�s���~�&���qv�]���z⾅x�������ZQV��]��L:���m0
]��]����p���138!��Ǣ�\��'�6p];�]�����4��' I�(ʯ��9i�,��]�v�_�~�fݮ�]�F4�R�ݼ;.}뻻���K��w�X��a���oN�ɕs���T��"�v.v����-���Z��q��,��T����]�*R"�l^�����	5ݸmv����D��ԍ�s�����ݸۅڌF��Q�LS�֏\��Xw���]ہv���&u�a���œ���&rF4J����\
M���{�>�/O�������ʗ�:_}lh64B���.���6'��윛��7w���n�����p�2��A����qDv�;�|��泾��%	�j�W����Z��� }�p���K����O��'l>�؃��Ao���{SC�y�/}��0�b�S�3�JޕBFl �{�m>��<Mq��m'��ba�V9�c���<�!�Oo��M�rv�;��qTH|P�{��{�{M�M�����.���8��;������DNqZs��vn�w��S��|�x�x*}۞�_�x��e��t�ǫ��,�Y��H��}���l]٢��{p���@#��Y��hy��]Z���|PG7-���I����n���.�x-,�H��A��/3o-m-���{7�;'����D�S�*t�-�zg���`�_g���%V��m޽8Y������g�F����l���ҕ2�c���vރ�#a��u�Ǔ^�o�|O/���z�d:��)W �b�xn��y�ͤ�����$���Ÿr���{T�s��_m!*]W�0�}�[����^�{��=���f���sf���)��=o[����ӱm;��<��i�qh޶��%㽗�M��n>�}s����J�w{�L�}��1{K�T��f��x�f�GG^8E�&`,ʈw�e�7���Oz�A�f��XV�%������'���dj����ˌx�0�uV/[�����yx��8�h;N�͇o�c�o г��b�q3(bg�O�q�3-�A����d��V}~og�7����Z䬆6F�-��Ĉ�w&������lT~+F�k�ƽLj�7ڽ=9�*�^5��-EE]���x�Z$�Z+���U�F�-\��k��Ux���U�Dk}z��4m��5�\��/�o�����m�+s}*��+�j9sWw��69_��lh��B!"�u j-���I��$�d.P�TA��U]���nk�5����\�U}�x��ޕ��70\�RTWڹ�[snZ+�b��h�U�b�Am˖�65r�7��^5[����<V�~uEx�.V��6�st*%���bo�5��^�ESEQ�^�ܯnL���Қ����X�+/�a�uF��hKt�>oY@�t��ڎ�nX�:�[k�-׉T컋�t����U�W8�������t��;X�^1�9��!�{%��xu�N���+��n��H��x�'�g�W�q+��vGa���1��:�9���ڏ*�Egڊ,�*oWf��^v'd��=%ێ=c:<�\�q�N�_�ی��؞�R��8,���S����}��ca��hC�:9B��-Gm�>��u�z8��m�.A���7\B�y�C���I�vӠ��u箻u�(�=Y�8�{kt����v�r;��؎�b� �kuI<��ٞn�-�\nnm����}����6�Gn��O�o&v�G<wj��e�H��c��K/me��ݻ��sSˣ�R����\�;���b ����+�YOt<q���j�.��`��獮s�����y*��Un�r��v��;>Bݎ�7'F��
s�i�/�Qڻy�W��79�b"ej���]��І�q�َ'�;FlY����ظ����n��y�����hu�y1�h��MQ��q��z8��-�Iؓ/q�OB&8�tb��Y`<�tpb��:)����a�a�-��ۚ�Nݍr@r�緉m�5̳p^^��B{�&6��uȡ._\�zb��3ŧpܭ�^�h�,��1�Dآ�4�s���ɘCX�N���8�&ڄN�ٸ� ����ҲC��>�������1�ג۞�j,�,��#OR�4�I9�C��[8��z�^�L�T�s�H���^n�-��n;y05d��v��v\4��pAэ���ݺnۭ��c\�J��N͔"���.;W��H��<s`7[u����Q��u׍�7:�=��'n*�wn9WMr�V�W�;�;��l�ݴ����E��ۍ�S�h�=��Eٳ��ku�W.F�ݎ9���t]�>��ݻ뮪�kEbժ������ ��}����n�Rj�N]��y�;��SA�P�sؽ����R1���u�"�Y���nZcK��4s��pv�a��tNq���4uj�u!��O4k<a��¶����n]��ˆ3��8Ãڶ���<U���f�R>�+2a]K��*n��\�y^�5\u�n�&ޘSd��Q�0��u�%n�����&�����������?���v�p������۲���t3�T�j�eɆ��݄AA �1� �`+?��v��ۄ���X��j=ï�f���Y�a}��wwv���Ii�YvoMc҅��2L�Z�&m�N�Bo�qw��7c#u5Y��x�m�]��pCKT̶�)Y@�J��=�/궻k���yۥ0!�^�v��
�|�kG[㪾v3vk��Wp�n�-���4�qv��.��qwv�b3�m�n����2�u,z�wS��׽w#�}��(��f��:��m�U����1F1������g��mN�	��v!7X��jo]ۋ��[+��Ig��:v��m�'�SVD��V�c]���vޟ\�w{�y��dc����!��x�\�#�{��?Lݳ��M�)zTv>n�A�.��f�N�>d�f�^/P֘&�v��u���V}��>�n��>��d>��5�mg�z񀵞	*3Ud��k�6�{ 	�p.�]�����Nt��kvnk-�w�����oJ����m�v�v�8�<@.�-��o-k�	ldѝ�'AxQ�s��4/k�w�C<�%^�`;��@�o]�����wC�4����d3����x�֘]ہv��ΰ���=H��wSy��U��	v<�C�;��ծu�����L���ȞJy�Z퇮�����������hP}-��en�`sk�p.�h��3"�[�+<"���xr���7�h��8��Y.*�]�~�[F�ӊ��&G[z���w>n5֢;�5T[�a����B�i���/"�G�a�}��Ċ;wy�ony25Gy��LO�`$�>��&z_�R]�Y����g�m�~�]l�Y���-7�ݸwp��b�[`�$��
�&wX�r�<��p|�sj�Bg�<�o>��ۻ��������<�ڎu�8i�Lg&�,���퀻�L��8��O�]�C���<���ʺ.���j؝���=�LUۋ�nEK�=o��u���~�m��ڶxۤ��.����r����>�sg��}�����n����������]� �֪��]�p/���V�)o�{���ބ0��ϯ�gx������}k�U�|�ֶ0�Ҽ��
x�����Ռ.�]��|p$wm&�v�V'~`;5�c�[:-���u[ܛ��O�����1��_�n�7�~{����oMae�k�bO%��Ow�P��Xt�㝔�::q�>�{�w]��>����v���8�L-5�W������vޫ��`.�\�+�ô镲[�<qU����w8l>���dy�Gs����Xp�Jc1��e�E�Ϭg=v��� ���4�n)�V:[ֿ?��2[خ�E�zd�^]��#97W)�(*�����m���]�ݷ��������\)^��v�x�
����w�-�&��1.Vy���n�ݵ����ҕ�vWM]oO�2�LfU����]�v޻awn�ꎫ,�sU�xl�n8l9`a�q{��Fq\��h.�؟n�ݵ�z��]����v��wBµT��D��k�x{�K���v��q���T��ȟT�<�ŝ'��]��Xz���C��}�'}�۞ؔ��<�s�R������; �g_[�9������X7ۻ�`dNx����w�y�J��5Z���\��&_Yv�ϱW$�a1l����piǒ{W[���;3�;�[�hy�C/G���l+��]n��6B	���y�\j�D�k��h,[���s��\�q�d���ll�sі�Ƭ����5�d�B���Ԯ(�Cn]�Ժq�َz+]��7u����~�>�v�R93%vѷ���Ӝ��}�lp �pGmN��mm�����o�n/+��uu�M7��p�W���М�`%^8w5�y,���%/�ƻ������N�󜘅�ih���cMU8d;���z퀻��ܬ�f2��_P������s;�^#8������"w�ѫ���`+�v�m�Y�ޞ�k�fS6V���w�c{֚���l!��CKgr}���9�50	'��ݻ.��/�-^�`b����"a��p��1������Z��$h���g�v�#l<�͘���w�K�Yw�������מ���^�K�z�9�n�9�z�b�:8�R�W-Cn:��:����+�����fx��]M/�����7nާ���z��mv��݀lߨ��%�P~�.�X�RT�3�y�EF�c(��3�n�ph��^�gT�p�2�c`Ե�F�q�9�=k�ɔ���-ъ�+?�Fu�{;��8��eӷIvYy�Ba��w�Nq��N���%�P��x���]ہvxk|��l̈�/�ə1|s��_�m�v�Xl]�V���yO��x���w�|�	0ͭ4�Fz�TC���aݶ���g�c���(�޻�����~/z:S�s��z��\k��E�D^-m����1ۅ�=u[N����m���p6�q�m�l���ySz��L�aMFA)�����@�������]ۋ�4��Kct�h�9�	m���"{����{�l�v㟮^z��X�n�έ4��n���P���i��wk�L���u��ҵ��o�vsم��ꣲ"CM8|a��yw�jH|���dy�*0U���)��vN/����&{�@9�	���*�M��kh����-)��I�9��>�`6�qv�mwn.��N0*[��k�]�0�٘����	��9����iD����q���[�qwʥ��G>υ�s5�gx�)�Y-����Wwr=w"�4=F�E�C��<��VK���[��[���7�۵�vz�^:˴bGx�C4A�r��Z��������o[�,�vś��W&rp������E��q��I���3��x�Ս�K-���	z�n���8�dlv��+�We���-�v��ڑ�ma���1�,�E�yL��\_w�o+awn�z��]�m6m7��q�յ.�n���cS�����zrpnk���k���=:v��`e5;��y^}�/$b��qx���_/�9�/8*���΃�AKB�x���LӪ׼V>�{�on7�z��.�z�Wd��6�]����ֵ��s,��������z��=�k��p�X�Y�6����YY�y�#v���=�$���1ڧ���4FW� 0x���=�]�醋VzT��R�Wz�Qg�Ms��-v/�j�|.��twfѧ�,y�r��v�m�˜5fv����\1�,�Rݩ��G���|�����O��ǭ�ݸ�ZŴ�;o2
p�4�A���1�"5�v7���.��v��v����mc�ݮ"Gf�s]����.��n����K����zr��V�n�ݗ�]�����ܪ��F�m�;ۛO9�o�cd�Y��S��}�/u�ju�*O��#?�_̟������6k�{iW;�]��t��}���Tw9uOs�6�X3O�sp�V%��1��&�,��CKɝUw�u�gM2I�ۧRuS���[#Z��m����ޝ�uF�@��p�����\�n܌g��������v�\G��,9m�����&X�����].��oU	m��C��u���D#Q//Giu�%���:\3N��ַq�nx�� ]n��鸬KhY�=�m1���N�F����I��m��ǖ�'K��:�V]��s=zޫc�-���;�g�����?t���ppjzM�;t ���c^��sbZ�7�
M��2p�ǅ2����v���2ڲ����\!�d��nv�T�ݬ�����&���ګ���wO����sǝ0�\�*p��������]�t�,��cLi�vT��]��z��h�/0�B�uV�T��(�(9y�)e�Z~����[��9�=�K�<s���֜����n�XL�n��=�o"|krQ/Ы{7|7���.�퀛�d��c檉A���4Wn�Ogj��.��]�����{���.�k�A7����IIg�Ab���>��]C���ps�8x�$�Y�j��=~˸�Kr�Nm�\paR�𤚹6�ޅ�}>m�p�o��U䞼z��m���]��U���(�X��jҏs�<�x痟]�_���Y���C#� S������&�5���W9o1	][�����Ɨ��d�;�¸����%pzy{�3BFBV����W֟��S<ǉ#w�Uzw��u�Ai�EK���O{�mwn �f� I��=�Ƶ���Y��wf�7i򶯭4�Bc+9^����=k�M���t�g7x$��7�����؜z��*xص���K;6����}ಒIq���':����>y9���`\=s��ގ�v��d��R��u��ۊf��� �� Ċ}�n�{��a�����S���O&�M����^[����� ���(��:�j�'97�ݚ��¶.�e;!�K|or��c�̖i�m0x��3e��`.���O�Ky-��{=>�/_��ʋ���o�U��
���6��w���n+��b�9O"�ؾ����b�;�z�t� n��Y��N���H�X&*����3��;��\�.�Z�\��s�O�E��}��	�t�Ǘ��M}�r�eW�Mu�b��xD�	��^\6Y:�G��X� /G�V�m���c>�X
u�Y��!��EL��P��sDlYe[)�޺�|����>����Խ/a:������"��%�{�g��&�z�!�����k8w��a����h]���xo�%���{�����R�Q��z���	�V�{�4�c�]�|���v���SV���f�q�VB\G��:�xRE�t���W;:�����{�y�'�ǂ��r۪VE7��ǵUE��Җ\n�3���)Kk�����x��[���X��J���l�0x,��z�A[��r]��XE>!ۿ�KE���v5�^�@>�|�걋���/b'=n:�/��D�M����{�O���j��p���ҟ�>��1�g������s5�O���k���/]=�,�:}(�0W��(X�u"]����9_ywsm�&c��Ed\d�+nwB��'o�8�Uo���~Z�/L�xv�|�Sf1Ὃ;��
E���������|�K�t��O�ؘ���^�"4mh���ӽ�YgR��ݓ�ɜA�x<���A�Ws�,:�s�����ǇwS�8�������7�Ĳ���}/���?�x����q���n��z�{��<���a����s[�J�n��sUʋo�/<�~w�:7�p5W5sn��;�u��r/�cm�ns��RVwU�Ey�jJ<V�kI_KsW���QwtQ�__��"ޑ[61�Z1cF�5Y6�[�6���\�-_��nm�5rƿW,FЛFш֊���b�E��|^6��p�m����\�"���VѴV#m^��^�VX��Z�K��x�E�QlXŹ��5����E���MQRh�X��k���{Z��+b��ֹ@�>�|;|gu��u3�\��S����ww!�g<>��p7[��9����ъ5����n��^����UqǱ�k�kh��mv�]ہv�m5�峲s�z�z�`���Kd�R�a�]������l�K��v���5��i�����@�	j�s�[sW��[��r�cĊ�L���8�����|~��]�p'.���'ؿ
��Y���]�5�k�{����}O��76�Ս���<,hų�*�7��k�ܼ#}Zv��n7eǮ�]���l4�h�������z��7���֛���v�v�<�w8ީoecݷ�AMW���X��8_�S��4���ښb`S�
P��%]y����qk��e���vF��-l;w�$G��s���\�~7���`��&{��ʈʈ���>��l'�o����`k�w���C��Ĵ�1t�
UC� .�®�����~��w�`O������G8�o�֫��PT�z�v�ѻ;m�����!s�j�n������v�][U��=��b�C]V5.h(����j�%��k��wp�IG�M{����L���|[{��R����8_�R�����j�wG�ۭ�wo�o��Ș�<�F�C�@�S�+&��z�[]ۋ�m�X����_�:�����p��њ��Si��R�*�����o+:*�{5���v޻awjnȝ���D
��Z�9mNgE���K����O�v��O�	4�Hw��c"A�kBy�ofgf��If�!+��XZ&��r�d�.�`�P��������{``s����q������>T<z�c�K�e$�OO��GW:y�+����]�ik��v뫌��Nѷ�4,KV\R19���ஷ�a᧳��cN����X��bf�ɖ�#�.��V�dd��A�P�l=�t6[�r�)ٻ]�wm5�nѱ�9`���xj*Wk#�ƹ������M���v�hJ7��ڷi�{\���ۛ��B�J�6�����r'�9'HlN�uծ�e8��X�9|<���� �9!�h.X@p�_xl7��ǻk�ވx᨞��a�4/��uu��\�g��O�m�p3��bY�����Z�Wk�潽u�Qr+%hm�=wc�Is�UT�5�^��Sv���]�Ɂ�3�l�U(Q0��<�5�(�����w�Wgf������}����xx��l�,2f�.X�<m�J{��6/i�I�[]�ݵ��\��7��+�j;w���]r�\��]�V�z���'iA޹����������)}����q�����ق��W����ݱ���8�r�<� @��=]�ܟ��ww3�15^���j���u7m�;h���`:�-�Ӗ����mw�����:&�X��_ߺN��N�^x;p#�}��k��X�|�-�]/:��߲��*K=��~����۩=K����qV�������8�����oron�2��hl�`���z�����O`mr�6pl0�����.�,cL���{N5���e5���Э�?�e��M�x�_��I&�y&q�z�{1*{�/�B��.3�(�o��ˬ3����u&�P�u���}v�]��]ЬQ!�Zg�1^�h�Q�m�gFCd�]ts�M�[M�~�l��w�n�'�)l��s <6cG#i�\���pA�c�'! aU�ʄ�-������������2kכ�ʸ�yW���f�ͯz;���v��v�gjmÚ�.%K�i�J��l�cз�WKpQO�켗�=޼�l��	�Sy%w"��n4H�]�n���ׇ�r��2��͹��u*)��C�k��ƛL��+�q�X�ȹ����
���;Ǳ\���E�OS˸��K!�c<2L��>M�v~����yrY�V���f_~����z�b3s�}�N��*�$�X�g�>�k6���F0�ݸ��x]�����ή�8,o@�8��3�����t��l.�Ҽݣ��)��0O�m���\�t���Z�[��vX�<E�� �y�����:�^�&IwlN	�Lӣ!��޽��O�^&�}�R��z����������ŁM��]�ڲ�BM�=g�������ԛ�����o��$�$�I�^oS��k�6��v�3�mӥ�8lK�b`.��v��^�{M�vw\jk�����3l��S8;x�v�ͨSa��f{���ح��[������{��}�8��?1���.}�F��┛6�.��Y7�3��r�p|}�{=si[]�U0[�j�3�gH�����������i~����~Nn_hWU���Zw��ԛ�z�퇮�-�4	�9�Y�=>$��x'幷T[���k�����c��]T���gc����;{�
���qn�`�)�gGs�M��UηT�qr�$��V޻�����g��Ю�Or��o^��F�W�]:��;޺j��IY��ؗ�N7�v��r�m��9�/}�G��N��b�^K}o��{��]���P�ۍ���w���ѡ���8��P���q�8!Z\c�ح3m��4�?3����әi��O!�f�%�0zΤ:�*CBt󃷽r��ݽ��	��Ŧ�)�&�ġ�b�B����n�}ܧT������A�7�I�K��V2uw�`2j�A�d���8�'�(���;���������8��������;:y�θn�>YzN-�0�n�����r�t��W��F9���\�:}�뎴qݴc.n��2�3	<�3��ܫ�>׭�v2���@sYN�E�7G���϶�vVQ�Ku9Ŷ�b]-�^��Rط�kv�Lr��9*q�1�ݴù��_���;m�]>*ٺ��q�Oh�lXn:�`yq�z�l'r�����ȕvmk���?C�����q<gu��n���,�Q�=�-qql�9v$���`� ������q��wp���˾z�L�7}b�kFd1����k������\N�N�L�����淸vJ{�Ơ�it7xlS�]�n��B��;jR��rڭ���zO��}��tݯnOt�hL�0v��v�����yJ����'e���wp�����_uB��l����{ܙ��w��^6՟Z~��eE�h�~��v�ޱ���7��:jYV�Cp��?�&�oz��{�v��m�h���~�8_�'s��ۮ��PM�/��Uԛ�z2$�t�s�`�Z�-y�{׸�]�m�����M�(e;xqMXڅeŦ�]w>T���]��������Zu=TͻH�f�����6���c�-�5�� 1���Kڧ�ef�>=���m�i�"����dȨ��P4hSt�Ա�w�9v�Ah�� ˆ�����m��SQӿ��.�&���|	�f^/�z��g7�v����g����v5��}O�WL�e;�G>�W+�8lE�{��^[R�-P�9�O��o��Vz�����t�R�pv��[S��}zu�SoN��v�.���]�IىF�P;N-,��٦�����.���ˮ�n�ԃ���~�|�w $��HH&1�Y�/�a�s��C�LSsb6�b+m",���O���`�?j�/��v��ѝۘ���y��\�މ�n�Ws����!k��S��qv޻͎��l�z����S{����d�-�
YNp��,.��w��UsW�;{Sjǟ���z�͡P㱲ɇ��=5�XM�]4�\�F(s
�7 �������f���/������r�_[Ս��kL0�/�{�)豹���:�e��Y��\�[FG=kÎ�]��}���.�]���ٍ������E7���7�s
�g�|��4p}�8"�m9�+�Z�m�v�]�xE�\�к�b�!�ߥ�s;j[)hgJd���趻����?#%�q�����L���ǌ3�,NN�k��7�^G����©�\�O�N+�H\��o���[]�܉ڍh��[�\"c�V���
r����}��WS�i�j�ә@�d���ޙ�/k_5f�-9p��n�5��}�&��� �ñ�eM�F���]�ݷ��fMV3;\ƾ2��Δɹ��ދa��տ���m�Ff�b�^ǀ�ojl�!$<��v`^�=�u ��M�A��o�����o��d*���;O�td�;� ��"�;x{�eb�p�x�@�{�=��p���w&{������^Q�$P�$�π��������ػk��?8S���h�3�T3=�F��\��ا�����[%��4
a�C0NZ��y�2ݬ�-��ㅢcOi�4���/=<u�
Y�X�`;ݵ�
���M;��L���)�ڬWN��	��-�20u�v����'�-�ܖr�d7��ầ�x���u� τ��o{��]�kn���-<0ݗ����]ۏ��-^�����d)$��w����K���8�]����@�cÎ��+j^��v�}��V�h�U-�pk;�w3ʵW~��
��<p�%w����Yo�1��Gg\K��D�6껑w���?�:�~�TV��W�<�������������]i��$��[E�E1X�cE�1X�Qc ���P�E�U0X�c�E����`���� +JX�c �Q0X�b(��QcE�V1DX�Qcz�i�Qc�E1X�cE�E0X�EcE��R�����"�
,b(����

,b(���ƵM�+�,b����� �
,b(��Q�(�,n"��,`�����"�`,b�`,b,b,j��X�X�101F0107�AVKg�� Q��}ȃ$�*�Ȫ(�H
����z
���3�{C����_��q�AS������}��{J�>�ou��o�z�>�
���@����ϴ �s�Ђ �������T��~@�ޜC�AE����}a>?G�Hz�}���������Xzl�J�4�
�REYQdX�Q`EaE� E�E��Qb,V+E�E�E$,�T$ _�@_�(�!E=����
)����(+ �H �!-O`��ߏ����E=�P<����xS�?��ϰQOR��(���>��ۭ	� q�a��&q��*
+a�C��m��" �+ǰ�߱�����tt� DW�h|F���������%��o��%��i<R�Gn���EAEg��?��ݠTW��C���|���{������a��a���PQ^~�}��H�.J�,��m��&ժL�"("��� � 	�j�m��mU&�T�թ*�I�U&��m�%�T��Rj�Im�ɭ��VXDa !�l�mT�[l��RU��Z�MkT���6��6����ɵ�mU�Z�%m`�EVXDDUHA*�j�%m�MY6��5��ڪ�ڵ&�l�j��mI����m�Rm�i5����[%T�l��5�Z�jMI�&���-d�d��[&���5Rm����A����בE(,>���_�}��_ 4�t�e������`r�t3ߧ�TV�	>�D��8�������7�qb "+�0(5` ����}����o�R���PVI��{%�|@����@���y�d���>��w   @             � �� *��(�((*�((U QY�     ��   � ��p�8   (��y�M�NB�Yu����d�ҽk�z��^�<�ˡ�h�ET��Dk۹�#�a�P(}4����H:���>��@ @�h
�``�������`ס��{�z�P��::t6�ph�(�T^   E>}�Ap0P5�2A���Q�'���=4��H$��ֲ@IF��"O�}�   >)������F����a] ��K��A����Alҏ0u����R�T�/    }���t���u��gEi�ҽ���h-�Q��:]�K�^%J'��>����k��Z��}��+ё�{ԥ�d�R�Ɔ���     ��@RT�'�4��L�h�4hE?&R��  �     �5@QU4 2h     =��M2�ڑ�1 d @���D��@ h     R"&BhFF"a��j1��Q�����?i���Q~�=�N�y㟣�<�DAw�t�> � �����b���T�&��"�K?���L?����?��S�Ob�aS�Y�:�<Q�i%6���2@�D�}_s;o^��������k~�TPAz�<󣥽��4��5��o���3Y���Ԗ����S��)�� n������O�*�'^,�{�xl�D��^�Yjy[���;&J�rGo`�\�z�<���Ò�ݕ��`rTs�dU,nu��Tӣ�����wD=����$��H���9��1�l�k�,7(ӊ�[كj��v.��$K�c��bf�����i
��*�u��Dn�ia'q�o :�Y��.F�v˦� �Q?\�zc��`o���h��o�.cK� H&M�s7���^Mx�'���>i7�P�ăM�κ �e��7�7��.��@�A�vn2
{�E�F^� ��.���n:�ߓK�R
@�A���Z0�m��;fT�z%T�<F�Xǌg-R�8������_�;�E�����l���I�XF�c��R��9�I�W�vJ�il!Y;ٺ�S骡����.�f�{{.ݪ�i��]ۮ�o��y)�(��/�R�N�m�K�v�y2�)����9#����12�ѧ-Ʈ���晓�Vs�(�V�L�a��$�^��`�&��'g{6�U�C�p1�o`
n*�9wo��s��t�Z3NcCٷx���ZIoV΃���i��4"�v�>;���X�M2o=�SZ�ka���
f�C#Z#4����
3�}Cs��y�vt��4�D+�8-�-��^��)��_�F��:���%�!91t`�P�Z�w]+��"E[1s�t�ma��m�\��m������x����N�gf�*����o^��Jʧ�9�w+Y1�L����ܯ���5�n�LSi]�v��f��,��H��:�+f�0n=�c��ߔ͹9wW�7�}a���eWS�{���JD�[�u��í��l���[�l|L�ެ��:f鰡�k]�X��2jwn�b�eדKvK1=�6�8�w_dV�ާvT��Ů��Ė���v=]5`[� �7����ga���/�{���e�����rA�ug$j�#j^����I��\=�i
�OrI���!�f�ja�6�X�8g��Ǯ��qW8�˳T���L��:�t��Zg)����q��wc�\I9��7"�;���I����s[%1k���v(����Z�p���-Gr���yR,Fuj5���ۢI]W/b��8��Ǳ&2�ڡ�ǰM��ˤ9q�:����5���"��[ѩ���>���x�:�-�F�i�Hi8޸q-�3Gm� �7��y�VST9�&����I�N��5��SC�.�ԧ��9�V6v�1�O6�7p�5�y�w�<�@��n���M}���G�{��������W�Yŗ1����4Zq�Ƚ�[�ٰ(R�d�;4Ł��s�Q�3�!�X+����زdȺ�OG�Wc��4�då��c+r�o�M�T����v�8��f��
^ۛ\���l��`C% �o�^�]�>n�T�Ϋ6�{k�F���0-ם/
c��7cp��rj��0GZ4&���k���0x���!�m�'�'ϩ��9��`+[�]�2m�!fuF#��֍8@κ�1W}:��d;�8� ��	N�L�`��9�'A|���s���%����m���CXr]A�^�9��s$�h̓�w/G��l�}�e�sS:J8���۴��f˷{m݀�&��8@�YZ͗f1.S�:�j��ǚ�]#sH`۱ݰB@�f��L��!��ϳ�,�K��n��װ�1�Yb4�)l�{���bB���s����rG����l���S�}.���Wqa��I�Gn��"Z�2�4#R��]�����S���]�ʸ�S<3R���7��U�zشq�E���Wc��&q���ݸ�F(D�eO��w��]���ڸ
������=�qG:��0���wf��#�&�^��;����c�D$2�I�F�v�}γ����0e��u��SY�7m�����L�h0�8T���9��`'��|^�VRv�1M�vθ�^Ō�5�*��6����w�u�رW�r�6�{�	�z�q��]��Ks^2C�3N�����o>��.�׏��b�+���ۯ;@)���@}bA+!6�I:�V<0�;��?,���^�)�
p����'�
9��b�V���+�ҵw�@;H��J�j=:���
���N9�Ʀw��a�!9F��̽�ue��]��$S�t\��v<�:�u�fv�g��� �܂i�����h�(o9�=���*o.9{�o7SZ�3� n��\}rh&ؘ�xE\��.�f��n��>��F�(��M�&�|��Gn
gN�Z~\�m�U�G1��O! wfZ��c������ �L���N@eN&ɫO'X�/Fnɑ0XM���`4��RY�A�	[�>/�7i����0�p���3��W]�fƃ.b�1���bޯ���+*��Fr���I�eK����{���.:@��{OW��Y��t��>����rr�>�^c��Q�D,ѵ�Y$B�n�t��YF���Ê�GN��w;э'[��q�|�;�IY%��<����<� ��OE��+�+ώ�,@Q��h��pܡeד��w+���T�˼�яhg���w���ךu��:�b��\�]_4�G�%��fCQ�7K��c�
�n�<�q��
Fj]*��!�D��j���<�2ۖY�p��Y2̕�6�ρ#wI���$6H���9���w*������ȱ��5'wn��wXop�G����ɶ��l���M�{���[;�F�����n���+���u�Ա{��'�]���N��0��)���vR�E�x����өq�\���G��6�4N��9<n�\5%M!{Wo��vv����f����u�0Ѵ���9Bp��&��f��<���^�v)n��������pK�l���R�8��N^��c�^�8$=۱r}X�xL�%��\��uO��{o]�A폶X����O��g	���%U�>/77�tv��@Mw�.  wl�{�z4���Z�&���&�[��w�b0e�n�̫�Mg������<��h=42s'�4f��i���ɷg"���io�Y7�;� |c��!��;���٪Ͼ������s����G,$h<|�;u�[����q��<�\Cb��%�T�BKH�"�"P�PB
�(�* P��!@�Ҩ+H�J��B"P�R���@ �"P	B��
P�ҀR��"J� R��+@!@R(Ҁ4��B�Р�%(	B�PR ��������{�;4x��/o�;<|�!@D;�qƹ�D|��Q������zϒ'ET_i��y����z�[<����q��}:x]zt���gto}cUP~���c��X�i��I֗�ᮾ{��xt���DZ&Sw���|3a��8�S͕B85K����B>�a�_�]����E4�~�Z{�fm���Ş��Е�C=��Ύr�0��^�%�20�˼�N�w�4��s��D�n�s������{�IN��*�B� 4L�&h�N9�Mg�g/%�e^��5f<��qܳ�����zM�K� H+�)ۭ.s�)��Y�^icK-�oڡ�WI�0�*�-���w+
�Z(�~ԇi:=�	Gcb�C���j�`�PI9�.��6�z���;�_  ;t�c�r�Ѵqǣ7�B)�3u���M��-m����p�O���ޣ�ⱯIf���z�ۡ��m�r��fP��RǦ�8S{H��a�}�ǣlS=�����U=<�LЫ�h{$��gzN<��ۏ(K����(�1�;��{�S�5�;�NC�����v Oy1=�p��_��0���Q��9�ێ�H��ϑ���^ʦ�}6Ω���6�pu|��ְ���x{{�#a�1��Q�&ul���n+�]2M��\�����4�3�t��,���J>���3�xuM���Έ��r��o�nv�=�=Շ��G�C��Q��L�=��=��5����$za�ׇ���Nb	��y�W ����W'������.�s}k+���)�b�ly���=>�'�m�3�{=:y��A�0n{}���#7b���=����^���s,� '{�G�kM8����2i�U�ݸ�K�ǖ����j�Y=��k��m'��J^he�gU ���]��K���|7�T|��@,8��Ӻ��������s=���ΔKaٜ�<�vOW3�t�}y�Fm/����Ei2d>�+��\����yX��`��GQ�&�|.�����0�o�%�O�e�p����I�'��~֐nd	U$Yku�����[�e�1U��1��Ś_A��nyp�&��$]��x�nHW{B��Û�h֐_�(MgC���/K�㋶��n����I��a�sybE�n��g	�������]�
�F�T�v�U�����T��{�t{|�������;��_�y'�<e�>�G{�u�6A���������ǯ�������w(6��*�°���v�쇺�<�s�>�<)�c`�	u���ܟl�kD��R+D��$�g������f�N/��m�����m;糗������q#�|/n�l¥�x���c����ks)>a/@&��������䏁�y-�@Ҫ`�Z���Π�S��^�r�7@�C�{�ǫ*���W�����;�Q�a�lh�/�	;��>��=�Bw�A�vV�ˡaXE�%�N����gǷ|�?<H���a�d,2�~��*}����=>�y<��fsKV�h ������R�������^���!@�R*ͦ��ic1M���a���@���Ĩz��#�}ڏ�W���3NFW��cdg�᫇yY��(���q�9g����$��hI����t?�U޸�Kס�LP�&<��z_o�)^�{%�2��=�^�ֿE�x��^t�{��/59�%����j]�[>���0{�=�ҟ�/#����7�W�9v?Uײ�gvG�sC%iHs9�t.���z��\�G�3��+|y�T�^&��:�֩�gjMȄV��D���!T$���6m���i�9
��M���L����5\o���)O6�'������uU�Nn��[�v��4����*Vq�w|����./������9�z�殼�;Nzޘ�z�A�� S�T�������������6j��&�v���	�o�x$��lk0�C�u�
-Ojk��g:��u�[��r�o����L�t�Z���`��R�S��,8�y��VnR��:�XdI"T=��>G��e���s�U��w���r�d�K�
w��^�V�x3M��P�K׫�,�����Z�H�nV����zŞ����iͼL
�0�aBH�t�	�;ueF	���Sd��ƈ��")����5��Ƈ%��{ݲE�	z��MK��ٚ��هwc�}˱����L"���<e��<
�y�].������w�K$r����Dzo��L�B�P{K�.�<�G�\���tT���\�ٵLb�KY�D��JU�P��R��јm9bnLhZ�T�ӛt�c�5��ٸ�(xr�Q�b��Iz}˔)�{�9�rS�K �ɾ�����E5\.`᭎:2<���^�*T�M�բ��Ϋ�u�hNh��[��2YV�������<<O���eh�m����8��sg��Ī�nA���m�t�5�}�P���Y��Aw���=d�Te�Ħ����i����,���b�uO?M]R��t��ǻ��|�[��]�º���gQq��*�y,�'s�	��`�] �`�֔I���?oz�0�ZyA����mn>��~����'���E�p���OT�"g�G/C9��N�]�F\���a��Y0u��m�@��65҇	B�B��ce��]}
�(�2ග��s;��l%�KC�U��]�Y�`�%��J�p�c�+M�u�=� H����ZwnK��|��ϔ�-^�zvw.��7!��ِ.e\�~S�
D����&3v��^�ʅ����ј^�Յo(k��t=τ�k����){&>W����8�i�3ޝ��NG�������������n��=�W; M���4VL%�����lȅ�=��9����i�gb���ʁ���v4���i���[Ow�x��]��מi����U�:Ju5��^�љYq$Һ���;LΈ�A�a���l�����-�w��vq�^N��FA8�x\����xMx�ԡ5%aλ���,�3W��T�/V��������2�;�|s}��x�)�ˉ=��8�b���齁/3�IҨ[y����U��ۗs}8a^�-���>�=V���URy���}�/'ݵ�-�e{M}玽���W��b��}���b��7�����֠eV$s�+���HX�ܻvI�����T'��/,�5b<���-�W�g�7l�|��n��I4a���C�W�.`2��G���b\R���w�����pR���ɍ۱{�A[le�"��B�K�v�JS�Y?vw�OoB�=P|�'_G[������υ�b( �E)W�uW�hJ���xw�$��3���n��^��(�$]��+۬��Պ�E�]
�nJ��݋ ދ�{�WM����H�K��.ׇ�v�cc��6[b�C���{]��=�'�M��Sͱ��ʍ�cN�7)����pc�zpn�>�m�la��r����]{W\͑�q8 ֛s�HλW��mk��8x2��<�uϧ�,�"�`\��x�n��Ѝj��6.�W1�=���X�R����e��X�w�����+�oR�n�C���8!��B�e�s�������;g�b�woB�)�7h��o")`�֫n��hCT�E�.��v���ç�<���zڭù��s;d�Q&:�.�v��I�<뺮��=�=m;m�UG�9m�xc�R�jFX��Ocvy���S�:��]���]xi�l޲ݪ����ǉ��[�=���I��n��Cc���\���ܝ�E���ki������Kn�\���I9���ݎx"B�M���>}�=y�A�������������gc��/�j4�r�5�g�E��t�+˒���p��N݋#��9N�k���zI�Wv=�Whg����OG8�#�Ll:�p3�c��W�^ۅ5u�c�dm�Gb���� ��z=a�qۊ-����"��G����`�@u��]93�j ��6R��e��ٷn.�F��M΋ugr�仢��]�wl�uq�*}�����VK�Jj�zŝ�w&켵�	��m[����'y��]a���h\i:ݹ�c��x�H�n������:�.�-�6�n�a��:׬9d�sojPN��l콫���O�GQ�h2��SE����q�x烹.�v�+]c���r��q���6#U0-�`��;V�r��1�g��v�|R�F�m��n0�����ڣO7��]��f��v���V��y���9sjn����ّ��kw9ܰe<�G!��v�v��\�a�wd�kV6�l;F������ T�:�n�u�=tz1ɽqo\i �cy0.;"&(�5��xn�8����sm��������nܳ�n��R+)ju̕dVdbj`(ʷb=�Iݒ�m��:�=v�ۉ�m��Zyӹ�\�FV�	���l�:��I۵�IڷM��/n�l�
<Sփ�X0���s�ݺ{��t�U7;	��sp�tmf�r�!��`�,��oGH;M����xrHu�Lr�v��i2 u�\�u�U����v;t:6[S�^(7.Z:�^�ݎw@z��[����^8+�y�8:��ֶn���5]l\f��1g���®�.C/^sƊ���E���uǰ�9�,!�n����϶���W��\�X��WQM7f�/c���P�1�����s$�l$j���q�gPX��8��n��/Z��/\oGN��[>SeL�sB�`�k-/	�7[��x�담k�:D{tk�xط�8�K��r��$�<� i��3sګ#筢�n��["5[��탇��Q��^.n�qk[�9�+�n*q;�]<)bܖvP�;�ٮ�=mQ��U׌�ӎr��ڜ�=ROg�k�ղ&�ש�<����C�ێx�Rg\�����&{���.;70��ݖ*28�vD�\���'���-�7���OKö�i�g���[�Y�<-�[�ț�9dtv}H�v��b��m�ռ����dwS�7'6B��T�v�om���;���|y����1Fknx���X� ��::8)�tm{Fy�bnS��x�Nؗ���T�&6��zC�)]��s�gu�cOm�FsӸGc&�v��!|:��"n��6��v�GXo3Z�N�y�9�sѳܛ=�4��Vc�X<���	2,��e:T@����E,DP ���v��\)����6f�=��k�A��s�ьr�봽4�<]X���@w\����9��AoQ۶�8c�ݦɬ��ܽ���E��0�=�ޓ]c�ɧ<[�Tl�C�+]6��X�1ȇ/=v�
�8��'v'�f���=i0�v�����\��{%��v�*�9���\2܃{��vJ�K�����
�{sΏ��ԅ����ͧk���8N^C�q���70�� �5�&$���>e��m֗��d9\=n<�����j}�4�n�4{s�E [����Gku��qT�ڹ��t�i�۳F�묉2���n�� B9ێЛA�L՜Ƴ\̰�n�l�u���vd�]]-�ٮ .���SM�+E4V�            UUUT��i�U�V��qD6㋯��ӫ����=[D�\s�m�aW��]:��OM��SV�8���K��.�v�gj�$�8�kf�Xy�Ɓ+!p�:��59�g��vsTu6��v5P���m�����a򈎒��j׆
Pqn7�L�$un˒8�R.��%;�II�f����u[�w�4�b%$Jd�j�D�H7-��j�(�@nU��S ��2p���9���.HP�&�KT�����,��-��%�
�\!V܊[�����l������9�y8�iE���q˫]�K�� �;s=t�t���U�j��Ou���g��m�2�D�`��[���6g�N����[�t\;���(g]N�5���:N�6�i1�n������p�����6ۮk�����Ύ��q�b� �v<�V�m��>��F{Y�mس����m�F����u�v[�cV�ݓ7e�۶G]G5>�L�}��v�o>r�9��� ��V{\�v��;lr�d5�ݗ�8�Ν�<g���ƅ,��h��5�XC��G\t�!�������V,nՎXg�\#)�M�]�ŵ_h�w�w=�����`�݅�8r��.;�a�인�m�|�d3�]�{lf��/&�����۞5���7c�\�.Οm�m���=�͙����ۮ���t&�8�'q̠]V���Թ"�4��լ�![Zu$�UUB�غ㳛v�pF�D�ӹ:��o{���ZO;�y���Sl�n{��99��aL���.���,HH7WV]F"Ҷ)t���=���o�a6�x�p�7v��Á��]�����ku���v[�xx��Mw�v픉�T�_'�����;�+$�;k�ā��Af��(�I(�A4a���O{���2V>���k��N����3���2 *��o.��or�<A8`���|�0C!�t5� Y��!��v��W�s�����d���]8�%ӎ瑼�g����i�e�����ע�|�Ƅ:�.%Cr(Y"�Z7X�*�GƸ�h��(h�=��X}[vDe'��>fqd4�p���[�"�O[���#����
b�H[v�b��^�Q*��x�!�Tm�g�^1����*'��E�bG�o&��z��:@�>� 2��Dv5�Y	3��w�}~u?&�3�6�x�\�Bd#��y�|{��� V�����z=g�������8;w�7	�����B8���b�a�dy�S�����F��c$q|� �� �}��QC>��󳾿:���G�:ao����H��68�n5Oh���1�j�O��'ǁ4�r�o�Q��l���Wwej��ۍۼӃH�g̅����Ϙ�H�j=EK.���z���#�|/�WeyYdAfdQI���"0D�]�ܫ�>8�^�+�5�.sH�SK��qV�1U+T�'C*��>4��,��t�foF"���Q�y��>gю�H��QwՕ�ۓO��!�8Ϲ�|���"d�8�2�$�O�|�'yS����{|���X��#�G��.�:��D��"<t����|�3z0o@&��b�m�1��*������8����x-��f7��4��<�}f]�f_���ܼ���=�=���;Ϸ˽5�)��.B�#��卅�"*�"�bi����Q�ᐡ����W�Ԭ!Q��A�����dAk�E���\��v�u�r���}Z�G!���(Ɩ�MH~;k��.���@g̲p#�3Mt�>�h��)�����}�ӝ~��� ��k�AƱ�L�Jq����u<�;�Z���X��>D|��7gLV*ǵd��`Vc`C��X�"<���M"2C���ST*����p�	a"��p&MsM�6�αc���5c�\kczn� î�q��q3�4{iܜ痉�z}ƻRW�Wm��nM�g&�#�#c���qD;���'X8�
��E�Q�Th���-;��Ϭ�Y�,�ڜ���z�����Z'!b9��6#|�'�0"����<A8}�̸l��W����0:�"�&V������~���%�BSY8�9����z׭i���wr�i��:`��I����x�D��n�oȌ��W��ka�<z(�����E���KSnYv7%h$�"X�#j:�删��Z�\b>��C�{O3�loG�V+�7�����.`���#!{�z��B�-�]��Gw���:�L�*r)�Sm��hq�Fޛ����=�@ �!sf>�;�x�Z뉉$�Ng�o�����X}����`�
���32ҹ{��cO����x�O��8�\k��4uw�s�{k`o"!ǙD3䞞
���`�z׌�r�kW���D�<ȁ���q�=�;�j4�<�|CLk��}������f�6�gt�ޏQ�j����&�������'/o��|\��}Ց�{����E�3���ٮc���ܹy��}��a߈#�Dă�F��]&$�-�D��,��^ow��������;~��8|�E�!Ǚ�
�W-��}�ӃO��G�8 �\҈�N�9��	h{)�n�v�n9k�����B�Q�]��հ3��7���6�4��k�l��6m(�H��������������lG��!� ��p2�`9;v��k�z����8�(�c;>���,������#�@��Yò��$��t۫��3OU[q���aQ����Q
(��M�,m�rq��"cX����������=�Gk_gn���A8}�̳�jX���,��X�m�.��^�z�j�y��� EǙ�!RW��{0o��M�����%bG���'&>5g;w�k`ad�<�$%lI�� �C>�����2�s�p�g�|���&%�g<�n��;��r˾s=��w��k[ǹ�#�iƱ,q���5�7Lv����י���3�zHy� �N��:g72%0���7�F#�L���}�4F��=U��/܉���C1�GF�uOls�'b����u�u����Y�l^�kuwcPl��7e0nՠ�y�ɺ�W4��m%�\��k��>�^�n�۫XD2��L	h
�����RI\wɨV�p��@�-||x�H101L�gr�>��Qqh� �|�y�	�5D�ϑ
R�}{��O���)�>�(Y�2g�YJ���uٝ:�28�D��T�4bD�+e�y�{�۾�"��<�3o�G�ָ�$�C�~�����!�J��f�`�8��p#��;<��A��&��ݵ�.N#�q��rZy�tn@d��ovl��<�dԐ$d{���K>�����K��E�{vDT�08�O����]�onj*N����ޭ��I�\9=��:@�����{��<NI\H�B8�'c����ۧ.�0il��!�@q�Q��Ǥ�N$x���;��{�����H%!ق���ɏrϙ� *H���ȮW���3��,�VUš�(X�NR�k.kLv=���t߃��fk���Q.c���(��e�]�]��ݽә�gȬ�ܻ2�%?�,�~#��߳���˸��F/���Y-г!�F����V��5���}ft-v{ԯ�<��x\K���=���M���ٞ���k�+;��De�ß]�_�92�;�pt əS(W��k�$���jw\�-
���˛Ѷ���zwFs}�2b�Z*v0^�H�{̠�yb�7
�sH�(�VĴ}�A3Ԏ��׷,ˠa����Iv���b�/nT	۪�w�8��K�6��yuz���n���/����c��tgKf��jߦ�O?\�E[���/���ބԣ��Y���N�Ć���I���UqjҼ;�܇d�#5�ͣ�4-f��>��w@ze4n�J��h��eȭݭW7�/6of˶��.ͥ�6죾���=�k���<��j�X���P�TMPj(�kQ--�й�1TDd�faIC@P4�`QF�
��#&���XaEU2�Q�sY�D�i^¢5�l��a��KE��܈��#�hZ-"* 
�ZR1�Ƣ�0Q�r+322�(*�bh,��i�F�H�)���&�
���Q�ED�ͩUTn2)MOE���}xw�۷n{ v�ő"�G$H��]A�	r~����BD� t��"D�3z�y���| |��Y�|<>�Y�_�:Hu�):��ԋ�@܀b9��A\h���{�߳�PC��U�H��2GpH����}>~?C�q���g���ʳ8w���� ��h:�V Kk��������C��G���đ��$A�$��.�]5v9��`2D��@�oϽ����������Jh� ƃ���Ǆ�7 t�$^�9"n���| ����~���g�>����@�o�jD�܀nH�3[�]wƎP� "n�����C�U{�}[�����V�K&*%N�Y=��36�1�?aTB!h�&ml������!��i�B�Bm7Y��ƘH���&�ȭ�����Yz��v?�e��#�|����}�V�* ��u1D%)����l�nmpE�/����{�����̍����Y��V�/v��<�����4�T��x!��*�22���9���4 ')H;\Jfĺ�n����dn��rͳ�y����>��z�sٻGA����'�*{q�l�mq� �Lm���;:��+�]��0rۊ�9{��{�>����t���|��)e���(B�}�߯�#���Jݷa�-�WW��������Wf\�vo\VZ�簥�p�UI��Nt���w,��(����QRW�2\������u�:RH��#��]�DK+�f�ozH��$	(�����������y'v��֚�E+�h����A�Q6Y(b��-$��_w^��UG/�P�ETU���{&�@�B�D}r��*g/��DT�ʵ�[����߇.��}�}��QP���(�d��V�nm�s��B(��z������$�M�p�]0����.��>����W0�Y�z!Gh�4�v8��x��(a��>��Y���m���aĒ1E����\�Y
��7�xe-w�@� "��*�M�;�I�85R��ӫ,�97=*% �l�M�߽ᓷ���ׯ�!%wDwf^r&��7�.���w2N"�"�;2�����ᦴ��=k��\�֢��R����!Bi�d4�|��������ەVک��.�ٚ���x�J>Ho�!�W.V��[ݻ��F��Eٹ�UfU������O���ݩ�1�(J���{<ԖU���T����v�4�������C
>E����ϿE���;���C���z9!�)�j-�@�jYSc���ny����yͺ��("vu0(�;�s�����YglefG���%�5[)^V�k��'�$���U	;����ޛn&m�����ڸtM�x�mn�<�$"
�H����<�A�������mS��M�Wau�}XJ��U��U�%��*5h����n���j��kl��!�n��Q�m=kq�;rٌ�<�FK�]�����͝j���'��u��
�j��)�rpy��T� �;>V��(�'%MAY�m�0p�n?xY� #ۏ�s��ve��1�D%7��ز-U�egu�	>���x������۸ޜ���!RR��E������>ݭ�wa�B)OC܋7�]��կ�B-]G	����!�0�M&�ۑʭ����qL	������s�7�vp� ܈"�	/ٓ���q��/�>u��-��.��`�r"�3:�����}��w��_�uLu�"m�A9*LpW��7����Wvf�I���8f��;���I��Q�!$7��{V�s�|�=�Xy[���kVF����@��XI6J(@f!��a��B+n�o;�xq�q+n�{���X��R��	����}$"�4GH��d"
�����n7�sy�U%\�^��AJ�1�<7���/߇���o3ﾥ���"�
��v"��>�Q3W�}ռ&�(^��䦫3�4܉ۻ��]$B!I��ñ�R�Q�rD7��Di@�E�ZwaJٽ����P$��Pg��j��_VoV���-�f���y)ٍÒ�f��%�=�3sj;��ٝԣ����������Le7"��V��%襄ؿ��Fs����OeD�Q��=��iD"��~�N��ϯ7�{�EY��s�m�Ohҹ�\�֊����q���()�]�Z�]\���{�z���݃��P���]�&k�7/��t�$'n�P�F�"
܂n7�ݻ[�}*P�v�(�
�e�f��$('z���ȄU����3�73s�>E��\e�;�tS���x�۽��΍�v��㳻܊�T�4<��z���0�خpQJ�`��Æ�J|�f���gkn�<�^S�雧}v�w��kge�{]�15{���H/�e����C�cM��%��o�� �!�x[��#��8�ӽ�!�Y�t�=�Ĺ�>;x��x~D6��.�k�<�p®�Z��t0�)R1IF�
PD&"��V�:�L;�'��g������仹*��[�{�AEٮ�g(=��\3���;��D��x.J�_�`D���FҺwޅFN��<j[�l�S|�]E�{�W���ڬ׻<o���Nw���^孃�[�r�b��їQ�4�k�ٖoM��H�l/��/h���Ŷr
�����Nc�sk�T�
������U1P�T:�)��h�톣Dd��YI1$BIT�Tb��UD7I��������)J���4CTSUc�eQP��E0L�[��	�32O-J�Dd�*��"l��.H�0H�Ji�FHU�m[���Ti�+Y�,ka-�?O��8�60pC;�n9��'��d�m=���ڄ�/W/9컭�xγb���/눶�b�cl�ƪՠ�M�����˗v۶��� �\�ڧ��vg���&v�[Xq2����TY�Y%l`��u)>u��G]<O�p��mBq�c�ŭ9���O�n�N���НG�9�`|:�j��Y�wm�]�QE��ٹvy���I�sˎ�yB��v�3��%������A�wf����9<\���;���q�۞̸Ǜ�.e����ޙ���F�X�8�N:K�h��U^^ɬ��cs�h�]���$�Re��Y5g�<w�+�vgX�^�MS���ʺ��6�b�C��������2�u�v��N�/C�n��e�%�:Nnⴻ�=�g݁;q�� �J�<�\���A�<�(���l{!]�z^^z�g{[r��j�:a��u����j��Z�k��C��-Obs��s��f���J,��VU06�·1���d�A�-�[q�p�����_$�^F���h�� ��Z�Y��Q�۠��#v�Y�����B��[�=�F��nk���55~��~�m���nݥ��ox�֣/b� �C����߫\Q�غ��J+s�Yݷ�{���n����RIm6]i����*_/2�m�wٟN���4���QGȠ�E<�6�!�����y��[L�JgrD(�I�%����Id��"*�	�-�Y}��޽�Q��Y�B�P�\�iQ��M�g�I7��s$�yS�3n'�v\I+c*&c��
*'#�� {�?����s���R�x������tkbY*EWoot>gȥL�T
T�����Ɏü��Y���7W��y�ӯ������6���rRZF;kv+A�S�8^%ۋ��E(�����ޅ��8�M�� )���TUV�owd���B�Q�Y�"ϑEQ|��5���D་��İ��zb`j��S�1V�IP
�� <<��vw};�� �T��ve����۹�	w���RQ�o:.;q���ʟ`j�s�zgo�w1������&`�0���dD7�,��D"�j�;zv�}��QG�^�(� N`���ޅ�d%�\�)��`ɇ�ȢÞ����v���G"�Gg���E>�����9��5{u0{;�E�CU��m��U��p6'Ɲu���'V��#���<=��$Y�P��A��<J4���Y����E�A����8�XX��.*r�J҈ii�#�E"�{;�*oTj�M��ꂣ��,�u}��;¦kr��!��BKz��k��sR��JT33!:�{�ݕ<����YQ�UM?:ͭ���*a����k������&�^�/PH@�!V�тVeн|�z=������0��uf��XP��\R�.'ܮ��Pk���ѝ��ͭ��x�kZ,c���ώ8��h�,wF�����v�N�4s��ᱢ2��c��������2�}~w�}��v	1E���7 Y��COx��������݊���qqYBE�u���ܹ��BgfI�������E#���k3�Q��^m�r\���Q�!-�U��8��vwe�y��͚�P�g��i$B`&^:�q8��<\kQ�n���,����z:�)2�(����ጺiq��!ɝ<]]0x�{:IC��/�ܷ�)eE�<<����tv����vnì�P���SqV��K����ϒ����f�{}�{�xQ�o'M���:8R���+7oz#���Y�p�w%ŢCnB3�[��T�n�yh����A�]{�ٔ�ELt�]5�i@D	3[��,!�1f��_s�E+F8����ѳl��jD�hc����I"'���ڽ�*���^���������U��%(�����ly��}��u�잺h�fI����7;7������P�}�����*ti��UN����(�Kj�7��b;&��me3��\TB3��J����QrL��GĲ$�(S�Fc���{޲(	3<&�$�Ewtv�wDw� ��X�\Үݎ���i��F����$��D��b���������#~��P��굳_}�U�R�(�;��#��0�YnP���a7Y��>E=���碪/�I#�L��S2�B��q����$��Wc������:M�ķ�{�w�RH"&��.�Bk@E[۫��4����x�X��SR$��{o��pE(U�]�}<u��X�v0\F�lQ0$�6E90��OxMerV�N|�XKD�\!ZB���uͭC(&AS�y+�s˛l�m/��@���u���mn]�r�q�`FN�nfpr�q�W7s��nX3F=����12��k���S��:�F����a�@j0�O~D"�[[۽W}=���QED����*�M��-��N�]]��Hq�ڥ#v��of���IƞS���s�����>Ii�I
[���[�u$f�E_�$��(�U�]=uV��}|��"���[��:+�h�(�N���%WN����&�Og�<[G��PS	a��U5~ �x/�$|~ŕ���U�
(��y�!$�t�)|�o��o{N�%"�dL��׼�v�����t�ڄR�����ޫ��������N�Z�8\ntkn��RN�Ļ^"�� E.j���i��s\�p���B!���6��[�]�Q�E�	%
�q��G��DJc.����Y�(X�œ9$b����F{�~>gڗ����*�;�$�N��-vQ�<���lS�4^���&��xD�/t=����׾��0��N�O{��)r�`g��������˹�	��Y��vHG��:1�^&5�4#ڒb��B7EVr�nݣ��ԉ��MC�kf[���j�2�]���X�t~SsK��k{���ѬG�;q{׈��E΍r۞�A%��~�~{w�6�ˈ!��D���@e�����%W�ww��6wdYw���wC���K�|<Z�x������mէ���t�6jr4�J��Q)a�0Ƥ�q���*Œv&���!�[�Y�9���Y�Ͻ�q?4�%4���YQE1-Dwѽ�MPTTAJQ�1�5UMM7��f�"j��E�PEZF��5ʗ&��]��F�6]HTETF���d��^���J��;���kctM��)�i$k$����iH��K�o )2�� ��~��}�W��G�G�\j(�[��f���
��.�J�V�c��Y۱��� (����s��p�!��M��d�Ӻ-k�>~��εUfgO]��a#.DL�!ۊ�bAZ)S���;�}��P��p��P��L��;ڻ�W"�Q��DM�WT����������f���Qo$��0wr��R�c&edi���܁��o�{���_g%�BUlL�w_�o�{�BQVr�������jK���vM�3�h����r��\�(T�i�P�N]���c*�z�.�ᙇ�G�,�a�c޽��ǔ%v��K�B�7z7�W�m�tBP�(�eb�+9��mu�>JJ���j.�8�Q>]N±B0n\۶gZʗF2���x��Yט��\q��x90\<�����y�ӻn�N�\�%�c���n�복���.�vq4Z�;�[u��9�q������=c<���<��t�6��W3�_}��߀�~��ԴN'F����)Ϙ��U�m9�{�[z�j�f�H��6:;x{{ur)|s��,#ȄB]�5;��"�r��gȢq��Þ��RY�ټ7��j�A��̄�	���������D-�[�}�zn�f"�V�i�X�-=�P���[}��}��Fqc���JFO	P��R%I-C׭T���<�/lo�����������|7��26��"�
"zҌٸ����E�WS��������Wy�}0p��� ��O�N4��gp����f�b �JXIK��	�7\�0F���k�*�E�gdf��WO#��pJ'��,����ɭ������o����W;�%�[3A�0^�r9y�r�'K�`���n���mh����{]���7���]\r��tF �23�e��*>�I <�bxD�\�l�M����:㶳d�@@��ն���t���}J�����YO��6�U�5��-z�Mv�gv�������D%0��[w��7޲��oH�����W���t�bn�cMS�]�s��M}p[��뇍�O&��++�����5��BK�DC�{>��ݳޢ�yj�S׻��W�t!�J�q��%#��R�(Ny����5�Otے{h�j����"r=�F�^��#��iF�� IJ���3�s[�{g�BJ�eݽ����˚�����dZ�B+3��;ݽ�wy�ƅ&�%�i�9�n�!j9?R�����,,k���(�2F8�j�6H�VR�����ݳ�$ͺ��S����^x�Ҟ�����Z� t/U����ݍ����;���`�a�9�1.x9_C`bFc�����ﯳGm���z��Vcu��l�U]B!���[�0�ҍ&!�% "��ι��鮲�59���"��Yt���Ν��;��x��T�e�Q�9ady�7�#{g�DD�1R�"�Ft[w]{{{;θYD%La�6!2LD�U�1XJ()HX��7�5��K;{7��F���]f�FCi
8���x���R�p%T�u�h�]L��U�nꐙ����M|�U�ّ��<�E�Q��Z9<ʹ�U��P�!�P�sN� �����;�m���2�Ȅ�ι"����̍힤���`�Ypp�(n�u�t�2����P�:o��)B����;rg$+7��(G�;�B)'5��w�C)g^��=*<4�B(�\���3zK�1��=�u+ڃ����Le�v/|��J�!x.Q߼=�<�s5wl�JEu�.����,����e�	(��[��nV�oo����;��p�ў��.������WM�{�V��7Wݙ϶p��2B(�EI{R�Ss֯7��P.fJS��7]N�q�}�"\D6�"j�3_l�$��
㉧,���\Pz�9�3}B	�w4�:��o&> y��$��j3sOrH��WK��WP��vU��;�wo���X���3���B�� �P�I�b������%
�
�B�;3u��	JjxTU@J.�Hk#a��һ�@J�=}wqE,����;H��вIC���Xb�]��|�W ���=�JPGL����B��&�0��1�Fw�X����͓>\��Oe0��[�c5f�8�9�/a�n�\jd:~_��w=�m�g�o�^�ו;k��Wc4i*'ui�1%Oj+����^�ԃ��=	���{�������u+w�]����w{�cH���K���'r���8J��ywX}�����^�W���Vo��WڲY������./ՖsY��jv�QJ`�L�KP��}������r$�Y�ZJ�a�{cƽ��v-�`#�3�h|�s�����-^f�):���Ӎ�Ǽ�uH^��^#���z����^�{=�2e�|r�s��ɜ�E���6鳻Ӟ<�.����߽���� ��7���<#�:T�]��ݑU��D�^J�-�i~n͹KBԻ�Ta)j7vX���
�Jl�FdCQPDD15KŒAB�.P-�l����D*�������(oL���#�Ȩ���j���(*��svP�UB���*]H�N�ˀ�(�ӹ'�N$��ۜ�ӰH�u�F>���x8��%ۍҷ)��=q[�`�g.�&�f�����̳6K�}& �ӵ���Ū�;��U������n������mb	cpW=��n1�����u���g��,�����s�7o۶^"բ�d�z96���&�s��lGX)Iw<W�=�' n�$[v��SW<�m����.H�s����[<R'�7]��.�v8�ϝ[�y�$��v�v��&�ŁE�;v�R�Sz=':�,�Ƹ��zɣl�.�n5��$.��v0r"�j�@ݬF�c�nۜɼ���ƨm�u����nGF9񚇠���5�-s���x�a�m<����7�q9�qb��<v4p�S�;�0����sս�v'�_�z�����b�u�<��u����׃�pn�f��5�(@X�m>�x��͓�t2��UT�������\�4��%g�k��K��T��"��M;%�1UQ	L�v�OG]	�!��G��܍a�C�'�c=Q�Ş]tkf<1�y�Py�箭ړY���R��kr9 �;FN�{E`bFci���[��6��\�!�Ã��Y�F�=�?_~*�ʜ�ͮ�η!�;q!Q�M̗!6�op���"�ԑ$2�Ed�0���޼�ݯ��R���v�,21<��Y���v=]��T"�ԏ]��*r{9���櫪^*{���T�Ăe#,@!2B)� �%7T�9�������Z�efG��W�J���խ.�ΘW�D��~��{��7I��w3\�}�jy۳�����{�ﳲ���E9*=)G�a:w�����9(Sx�]ڐ����ս���j�E�T"�EC�u��r�+�o��׊g]���\z�rIw`�St�48l&��6�);��֡�{p�b�iEQGK��	��ڷ����$u��,�r�S.ѧ�u�ӹʢ����H��}U�Kʺ�C��G��w��:�'�1%�l:�\�	�A+�՛�8n�
�]�������[���}���Z��uե$U�V;cU�0�����Zv��~߽��M�;|&2jE�!$WB��̵��;z�6�\��E'�T�B����Mgv�JJ*��Q��c����3�u����&c8��gz�mУt����8�M���M����aFmE�����>E�πwB'��ۣ8<Q��̈�R��3b���v�j`2��]x��U�w;�@U�d���ڝ�����gx�D:<�b�tB!Qo�͖��wf���Mm�E5�Q�ݫ���*ڪ��(HFrc�.*{{{�8�v��[�ݽpnrlɹ��C��*���wff��\���j����g���=��PX�o�mOsѹQͧ!�ig�ܞ)Aؒ2�][ث�M���o@%v�g�����g��k�8�:�8��Q�)[��n�X\�m7_�����ga��(�M�/���6������dG>��O̧�V]󌨲i��voj�\򹨋�V�a���4��ݮ�;��C�D�U�^W��q���ys�&#��E�� 6��#n�yQ���-pe�AQ���D�ٹ��l�ƺ�)%=��M[,ʪ����TQ�ʛm�S�ʦ��'z�t!��X)��SOy�պqs��b��'�j�����_x��\O���}����;��1k"�TK��;�ѥ�F�Oczz����`�n.������sW�=¯����^��lNvVdFe`�����k~�H+�H���d0�!�%��Y���cV���g��|�"�b�bm���9����K�qm�#t��g�P�-�E�j#�錙Fo��
=����-Ş��=����:>�J�Vwp����6�A�H�h�{������q�gC!��)On7�w����}��|�y����jJ�DTb��Q�D�t%N�<���D��-��鼊̀aھ��g�9�I�b_p����o7%oD6;c{�p��T������٣'�!��g����M�-����H�b63Vt�UB�9�kw��V�j���[%�Y���_��i�"L��BD\ؼ��g��l7n�'`�@w㔻Iԍ�˔��lj�I�=�{�2��_^�V1�,��n��ݲ������sQ}7��Qe�p�r��ۚ�wݳ�p�g��dW5j��]�mþ�ǽ�+�ؐ�HI�-ǙXP�v��Uv����W6�����]��gD��q�Y'O���y���G����3�zg�~�~aA6�D$W�-ym�[=Wb�1ۥ܏!� ���^�9����C�������9_cvv緺��[�e�X-�i��n<�Y�ud�2:�I�呝���RWW�蜄-h�E�6����~�Y�d��gݳW���$��3��i}v����[�2{��!�S0�7�^i�۞Y�s��.�ۨ����̔ɭ������Q��wmx6ӎ%�MT�u��я��nN�]���p�8��^�+���mN�>*�ը2pwB�{�p�][�.`Q���m���>�v�����I�D�a5#hn;ȝ�m:Oyf}�{��>�j�s�;Rj���u\*Z�t�^��Cmy���닯]������T�2@n<�����ٚ������e�%�d�|���%ۭ����],6�(�U�Y�[�os��:q���̊Edy�[�fTEQ-D
����5r󈮎[��k@�Y���
�ݯ�>�<�~��^	�:5�>d��٠��z.��g�R�aN�x�J��x��qSq�"$�QF��މ�4Pc.�^i����O{���#��ڻ�	}Pwp��!��%<��������M��ۣ}�I��Zj�>~=�o���'��FE���<��U��vY�J7^=��S�H����
�g,����.�\;��ӧ��w�Н�~��_���^6tޜ
��tQ�G�����K a�������12wa�ѹE5�<�e�K&�e�[�z��֚��
���Mv7dѩ�
�=ʀg`^ �v�I��u]���d��LhK��\an}�u�p�w��=��S<� ��b�'�g����̝��������
j���D�0P�Pt�$�9�\�h""F',��(�5c̥��IMq4�nL�W#*��	(hL� ��8�tEY4��RjV�
8��
�NFdI��SU�w)hA��l��.@U ����QQ*:�E�R���"Er�Ơԭ?�y���{�]|�����l��m1.I������*�wF�Y��:�ps�=�c&L�	��{ڹ7s�w�y�l��Z���#LL\jT�C"AMں��OvY���S1�������V�fd����+�8l�*�biT7��s.
��{�4m��b\;v��wm��j}����*7g�2�m��1�ɖޜs��.�T�9{�ub:��%4,�t|3!��p�t!�}���cm��{��Ne�^M��]�""�#���[e����-ǃl�����4+g��m5˲����Y����!�p���*ʆ}'��>n)u�<��޴�m]vVjȒ�-]�����̺{V�v�M�CnUp9h ��;����q��7����r)���&s.�6�e�G74aOPDiC��jv	���P��)ǚ�a;������=:���:�7h]�9�;��᭶�����T��=C��j7� V�;
��pn�t	��Q��v8y��7��_90��R�h�w�y���݅�\����m�a�-9�#������ĺ�ca	��p�y�=5q7v�'<{w�xi�]3��Xʼ����,�omF����7���J��7���o{�lE�f=.pt���R��_m�w^���>�y�Ϟj���%B���(��MKc�-�A99���Y�w��{��̏1���3��.���N������έ��ۆTS�����L���7>��>����Ym����K�ɳ2�Po%�*QJk67��9sA��]\�ݶ���[�UH�Gp�����L�6�ef��J�pq>%�s>Ҝ*jA�jn�(��֡,D0v�l]hxA0Jg~���fV
��.�,��O�&ݱ~ݻ�[��ِ߮�;����m��ܹ�z�R<���~�+���<�1=�Ǒ�硜٘��/V�wmv���C!�ߪ�������Ä泣������N�RF�2ۮ�:�0��)_l�q�!�N*���O.HER�qEm�	me�M�z�cl���gWl�C"6����n�r�*�
��ݾ���|C��f�,�[�5�"WU^.�u]�ʹ�W:�1�Rd�ۼ��u޳y[%[ZoU����'�iV�����微wk���N_�J�������4܋J����y��u�6�|���LQQ�D��	B�Sq��[hA�ɫ[��7���2�>H�$c����`w�[ߧ�)��C�k�)J$o%�
������m���U&��5k��U�`u�k̆|���%�<�sw��j����"�D�(>�a��;��&�gEVjZ��Ųr�|�`��Dp��-s��z���\:y��[�BG�up���ۯ\�^��n0n:����qn��*�!Y�x�ۡ޿o������^��rW&���A����d��m7*����%eu�ʁKL�����x��V
(�\�O�(֣��u�/���s�ԩ��w����b5E���׵�U\k͖��2$��j���V�Nn�-�#�-�<�f$�=�W�7�]�a�V.��㛉�Rb��p�F�j�(�!�8���&��3_mR2EuSA��cc���R�]�\��ה]�-J���鎪ݨyWM�*g������a�}�>�������n�-���1�1v\v�l�>q�m���!�l�8�3y�������O��I���r�UF��h��+�2=�zs����{�
�Ij�u�8�Jn!��GHn5���{�u�;ɕW��v n��7��f#�{;35��p�o0��Ȼ�e���Z�����8sU�I2�g�rV�e
�ڗ7<`�TE�S&�N��χ�����߇�<�n6,^�x��wW���VB�cb��*�z���ӎ���1��;WmWe�D��o�΅��ya�!�eL�LJ�2���@�틭]��]�����I����4N�y�><�*���V�uH���'�GHm�VEu*��[|�g^��(u��Y�h9�y{��|Y�S2��&��o,�ܢ"�dUȠq����]à�}�����nm���ׄ�V^�]�/Wx6v�EvM@��7���q��tb5uۮ��������lv�p��D�&�L7�4��C50N��o^�r��7=;�qE�����:s}}9Ϸy2�B����{��ܫ�;�5ޗ��T�,��z��M]wc77������>�W�Z�옋7�h���[7/(=�n�֬U�3e;	���[��� �K��ٍb"�N���( d��go���q���,<����5K���]���2狓��!~�/��~8�\���(���¢�eg�U;7��UY�a;��RL�bol�!dm�u6��n��F�t)�k̙Lɛ����i���;X*s�=�N�=rf�]ܜ���4/zz�^��P�2��Gkc�K���B~Pi�D�3U�'��l���$�ʆ�bSIL��Ö����r,iP�APr�cV�!��)�ni��A�=�|�<&�^�sȎ���.���U�}���{g�H��}(��b�zC�
O	�R����A����Һ�%������&���5&��T%!����QMqd�0�(i�ʠ�Z
���������&�(��
Z8���F`�p��V��7� 79�F��j K���.�p)r@R1�iB1(P��T#DB$EPR�@�D�ډ��VW7��f`�����kF��Q�-r9���*vV��b��;dF7���]K<��ugv���K̴9���]cYɳ�y��-�ɖ�l:[Z7<�ˍe͗$�ɞ#��C�S��;up#������jM�ϩ;�Oht�qv*xN����Ls��Pۄ��M�7/[��`"�gu]��ʛ>�$�����;;��nr�{`������g�į�ڎ��#�ܹ��F��X�ngx;0�ct�:���{!vG�c�]�@�y�{m΢,[���s��iZ��8�Pxq�?]Żpptnv�wŘ���%�5f�8�����Crq�u����hٰu�s�!����n�����^}�ݺ���x��k�Z�(7R�w�U냩��.�{f��Ka�4WG ]��U�mh<6;9�s!�-vŎq�h��i�A��]��rMm�8q-ʝu���=[�<��c�FXv�T�n=��kV�2����UUT�Z5וst�n[�2�h���-#v�_�{ܻ����C�y��KKy��N�a����dU�!���e;�5����k���ݫ�b�u�FA�P�NQ��rME���чW���M�}*(�T���P���I��븸��e��ȝ�[n
��������Q]���x��aQ޼��Yv.Ys�s$H��ӽ�]$2��ڥu�2�x�vq�����I��ޛ�t�
_]��>���H��qg�1�Y�Ǧ
�l(�up��s���&�Kw=��m�0Ԛ1
����S%@�Nql�`p�x��vWrݑg̶ѕ�P5��"9������w(^���*"3�v��0��-���x��J��{�|�n�;�5OL"1�p�;;���0cP|�0l�鱛ټ��X�my��q*��F�Ὥ��}���+4h��u��Z�e0����Z$�7�(V4�w۱��/��ˑs�p#f��Si�]m�v�oq�ƨS)y��p�{��"#������-��3'lC���[�1�V�p��mܴDmZ�� �������͎p�VA�3r*�����ܗ���qg{~�n<�UOd����9{ٻ�SAዋ��%jQD�E�0�4&���P�h'x��AK��~���ǽ>��lӬ�/��g��uv�p�ڔZ)ϙe�e�1<Y�6�{w��ʛm���b��J�&9�^mt���7�L�r%�.�dWs���[�ܱ\�wf���7)����/�2m7�zj����͏�k�N��9v\zɹ]��ƚn�GS. � M�V-�e��k��Զ���8�e�� ��b9�gmt�jO;1\?VC8@m�./koc�k�-��vAww~��=��y���H�5w�S���m�$����o8qm�EF8Z�[�%�P�D7�H�y��y��j2q��
.~�ĝظ�4�����Ss<m�/�֮�f�;�s�<����y6�cuHq�x�]��y�:�ݎ����ݎ��I㌑.���M�8c��L�ڡ�(P�{�uV�q0*q� �b�m�N������nѽ�*S�<0�C!�O�M���Qyux�w��*�U��f��d6����s�}[={ s��F6�w@����wUw�{v�Yv���!����D�F^����{��t���^6�Uu�r�aj0��bBn��6��]5����N��-�n-���#�tg%�sg^lD䉛6��d°�[��R^�t�d�π O���ӽ}�n�s!�3Y�6�����Cz��I�M�n�O�6��"/��lʚ����^�Y�Ȭ�ɜk�e����t�v�f�n�pm����Ψ�\f�E�m��`�	�:1�tp��}6�b:w/'7�x�U��t�k�ξFF,P0������Y����Q��ܒn���n]B���F1�i��G;��4��M��Z%���'~ z�sw�73�p�3�}��\��[�ٙݾ����2K�m�����t&S����װ8���x��>N+�8��)[v��TĒ��!��ۀ����ލٰ̝c�]Ǚ��X\�UL&rr.�{3EN��4�����p*sn���V��m�rc�`Ic�f�=��Y�Fk*E@���ʡT�ʃ�*��$郠�Q�ی�U����	��nn�`K�����gv�
T�r�ۉ��&��#X0!�&��`D�vڡB� ��kaE9�kٵ�4'��oq�m��*Q�ȒU��������[j����3�[�Rx��UWݹ6�W#j�ҖWN^�)��݉Y��d���LP����緼4������;$�J��o?D܇Y^�LCeW:iS��/"f�Qd0b�LR����2�y�ѱ8���5k���v���v���E;qdw��L/nch��<k�gv���p�m��9t�8��˧�؎;rZ�� �]��P(��|$Q:�S��B&�i�IUE������	3�r��������̷��0��+;o6yp���36OOf+�o��OxM�E���׷��!��g"ir�����]����Q�N挶�-�3���w�ˀ���m�ا�kNk���%�LQ)S�a$$(�C7gՍ2�&n�y��{uH�ғ��%B�n�7����NI���`K]��[�ua@S���_
صu���s��T�C���!��y��YoE��ܝ\'#�i�.�Fn�my�3���/{۱k9�9��,��x;�c'�S�[��۝j][�^c]i��,�l�,���%s͈Q	�X-������Q.��b&�9��2�(%[��*2f�{�^���v8P�n��Ym���	�������%b�J���e�A��3��V,mړ{�4�5�-�K�<&�[ùF�⤅��U���O�y�ڟ{����ݝ�R8����u��o)诏�ĺ׮����N���3����ov�����X��}�v3��֎xȣ��C���yi����ڶ�����o�sޜ���#5{N=�<�g�/$�o���{�����r���mF��'�����NL^�f7��a�O��A��ɂH��e��J<���ي�{d�&�҂���ǅ^�8R �;�~��O�m�/-G�|��
}@}��������N���ZV������67��Ze�3�*������O���{(�� IbM�8�i��g��]L���
�U$P�Q�-�X4[��R˲ꅪ�h�C�]AN✜��D4�E�5.��56�ܹd�C��8��SM�
 ��MHd@d����j��5	�T�!��)h�@#A�-j22WV��Ԯ�J�b����ѭkQƱCv\Kę�P��-,h�� ߼��������,�0m��U6�Wם<��YF���m�8�.H�1�;}������;�������b�'m��)Fن��W�-�+������40.-�ms�+/h5�*J���|����0\r��f,-�e����ʙ���癸���{MT���]W۽��kC��B�3Q�I퉤x�4^������++3����?u�a���8�U;�����d �����|�;�����!b��6Q!B,�H��Z;m�R����o�}��6�܍qvmĮ�]����T�fd�LKm�D��}��ӑ���fH��IeC{y��3{�S����eF�nsk֟n�[K3;{k��h;���iL�Z���x��+՗�� ����tG��������1q�h�+��F��C�[Y�z���W;u�b�Kq�������m��]�ӎ��^	^�s=�a	�C]�ô;���̼��<H�5P��J	�B�t(�y��}�w5�ܱ�A����n3๶��ٱ��{:�Bp�C$n�Wwl�o3�zs7����t�]ښ��߳!UF�M<����R�m�zU4�T9\��:9����Sp�^v��	�0��t���f���[��l+̎�qJ+%��M6�j��QT�Bzo�71�Ow���1�֭%`4s�aq��L�0�[#P�t36n��X��J��r�-�nd�oܱfM��GϽ;i�阒���33{��ٛ|�m;Nm�uE���O{w��i�l�5�"�A���{���=���ӑe�7�V��\�$�Q)d,�����hN��2]O]��n�7���2m��ӆ���T�;s9K���߳)Y�r������U�U�k��5q��%���a�)��h�K2�O�1�^}?	Ȳ��ю������UV^�v�\\��UI�mOTu�6�]k�������m���Q��(�-��dc+u%�r�$�^gO�~j�M�Z�{���������n{$���u%:���Z�:�#��Y���;9m�v��o�v��`�����_��'ej��GZ��͂�0����߷��� ��d�& �h�ɂETzH~�>��ߣ��}Yvt��_C��Ƒ�ꈛ7�<rJ���^���{x�R+�l	T{~>y�L@ �3+�z��\����s{>��~z���u������~�7R]ZF��QX�L��J��v��L^Le���U�;����fu�#���>�r� ��C1���2Az����ߣ���|�;��߿��nW����ݲ�ֵ.�Q�ͯ����nG��D� ���f>y��Q�#�>���5��{�χ|#�$Gv{�/��z���X��ag����;����>�?Ml A���#3�PK2�|�
=�&���-T���Ԍ�8�F��:?M(�5��3C ��:S�5���:�햎���Yqa<m���e�԰�[�m��'mkn:�V������g���A�λ�;Yz����*�**Z�����!�u� ����kE>/<V���W��R{��϶���n@�*x���\ �z���ID3X}�(Q��qt����p�>?����̱*�/Q�$�2פ�߲�jy�������aG�������ˈ�� e��D�/o{v���m���}�s�쮦���Z���������&^;Ǜ��p�>?�d�&w�Ν_+Z��REl�ێ4VH����8I�o�>��L��"뫫����_�~�x�}�:#�����܂��]p���9�3%}�4͵�R�(X�:��u��9��4����<�j\��.�>��Y:�s+�xm�'f �n^�~�P ��}%L�l��vr^��3��w�G���-�9�'ʠA)zH���~ޏ�O��kcɩ��6�V���!�u���ӷ�ӦA�}���ﷆ��I�����5B5�+I"�.̃J*^]�̐W��G�ۄFO���Ur��ϻ� ^�?y�">���L!q�������8�^"�@ں���_}���lzO���;:��]H�����7�'�{�Oo��$��i��65��;q��F�ͶF֙�3�j�+?�k�3+{~����@��9�O�����a���A30���y�w���~"��s��}��03�H&`A=����f9�i}Y���}�	���`@2@���ޯ�]��31��<�9x�F"�:zx�_at{��A�^��0��n�}�7>o}�ia���8i��>����{��2��p�&������χ�������ϺƋ�VǴ�$�3�fiu�s�j����?Ml�SCvV�~��wS���\q5=����}�7#�~"oI��)�FG}�Ɛb�U&�E�r����޿��O�Ε���� ɂ31�!�;o�>�}�gϭ�w�w��ҿ!�C)�#�盼�>��A>���������_]�~y��d2פ�����ޏ����Ϡȏ�|��%zջ��	Z�6w�?�|��^1A���'��xv|��3 L���߳̎<@ކD�L阨�VR�>��{�	�Yn�a��ͳ�}����S�oe^�����~���ձ�DL,������&H�A�A?}�ٙ_,A����ﷇgʽjl"n��Юi���>����Nww��mC+�+�:�1]�=+>ͺ��ª��!���=�˼krx�xz�?��֬�y��"�Wy�g���Eh��b�cH�K5�ðsov�n3��^[R�RsO�K�o�i4'��>.�j�(���'׷�>���svw�Vs��)�>԰t�-f�읖�����X>�w�i�K�.�m ���x���ox��.���d
ܓ�ׂ���b��/U�vm�=�3wq����N,����]KVn�Ƈ�����i�YxR������p��o���=yy��fx�CIv���sׁ\T�C'c�پ��,�x2�C5h84��1��ּ�*�b����'�ieҷn������rZ�\[ũ�w%��3���3y�y9�v��{r��9��ls�v����U�D��T��F�ZT�Bd:��+�� ��oB�)�9f�u4P���C!ܮ��r�CPHJe�w��5	�=%�:��7)�	Z!2@7� ��&�1iP�.�`�I�rC�Cq�S#%2CR�)h*ե(��a<�2�b���e���v�b��%8�. c��ƍ�7b;p�y�k\[��^N�Ƨ;YÎ˯Mvjջ��sa�}u-��;�cQ=n1Ӑ���m������U���Y��ۯ�����۷]��͇a�;up�cz��gnvw��[��ݯSl̻���#q��ܻ\\(9��-V�nq���6Q�u�w<�4�t�˻Z�-��/����0Y�E���C��2��-co+�\�.s#�q��u9��u�؝�ڃ����z�u��Zu부�b�ܻ�j�i`�3�|E��e��S��*1�m�q����շj�m�����q�n���I
��|5���v����N{sV�v��!"�p�\=�pV.ޮ������z�Ls�x�=��u���s-�W����Uִm��:��u�;^�ݒ$��)��nX�K9�q0�UUUU�\l�N�����l丶�p�a�8-�k�э�;gA���ҝ����s��/��nz���b��nLd�h���B���VjnR�X/�3�l+�&�������zk�čX�&���Tn��q�q�J�eQ��i�Q?��>}�� 7�igݿ_�@��!n�� ]����&`#'�a|r��v0�Y��������7��O;?a����T����X���>֥��\�ۼ; |t�`	��c�Q�t��1� �f&���ݿ_>��glڡ�af2} L���{��g^w���>��F2@����{i!Qqa��ù�st�]v��a]�<��#22`f���'��xv�N�<>�@�3#�c�|��"+��E��:��~�B��_X���r���f^�A�aM
�G�_��&��e������q��>t�2V\�]����#H�K�}�e�It0oc�k�;�~Yr=$	�� �V͐.��hf���w�ö��k=�hM���m��Zֻ��~�J�u�x����G���zO�LD�ݾ5�/���W�Q	ᲶH���Z�N|��}�|D�yL�����a��qi��q��Af='�@w�;����x�#����g���;�|p�`	��C����Y�n='�} ����.X�K�7k�ZP���Y���;�]�G1)�����UT���Wz�wk��@'��At�'�`@"e;�J�$Yv�����o}���*�g�M5�G�J܂�A��4��v�!�߷{�߇o�t��ݕ�}��߽��U�H�nܒ
4�
��d�TP�zM7�b�(�\L3
koq��}?�@�{S�Yj�3�H'�=�}^ˏ�A�zH���}ֿS�e�u�|�p���-5����d�H��'(d��+;��v@���	�&]�l ���ɨ��ݖo}�{�}�Oþ�q��i����S�8�;���}�"Vb���u�ǥ@��#�R&��<�^=OR	�v#�MCt���r���7������A�<�0}3��x��u�ۮ�9��-�&���v�7��}$��]������|�{���"w��aCvb~�����Ț��}��<8��x�!�zO��Kdf��7c�}$I(/INa�_?���g��@���vu�n��g����̅�b�5G���xv@��G|�;$���zJ>��D�I�����p���Vw}��q 9�I���c�����S��T`���>�W\�yc�hS5A��Lަ,R��}��:���I���j������{u>�Mg�x�v6�����Q��bW��ͣn��/8I�Q�;t�\����^�qԺ��<��\t���o>OUp1#1�n���Ѷ�������lq=���)·)���O��3�0 oOfn���>������$�����@�"� ���W}��9��D���9�߿{��a�}b;v�_ïow��O��ǔǤ�Af*o��H4�����È� 9�I��"e �rB������`@���w��}G����HR,zƻ��d�&���=��n��������"H1�&���~�F<8��c,dq&�u3e�ߟ���K�����&bg��5�}��q�v%2G��F��`A)��o�����W�oAǞ�������/p�{@�UԳ�C�}p5�ٛ���?@7Ј7����?~홽1�e|�ɨ��n�C02��������vG��D�L��'�P#�?t� ������3^wܸwҽII�y�ӎ�q�Z���b�Z�������y@�������~ ��DYd��9��"=�^5~ziQ�����&6VYvdnᗞ��R�	��Z֣�W_�}�; o�զH>���)�IG�1�C̯a�쨚߳r{�|;� 9��x[�>����������S`n�֣��<�E��bɈ�m�-T��4~�7{Y"���֖R�5E>�Q���Uf����=�X�k[Eݕ����7����J�ї��}�������]���z��0}3�&/q�\�_�ٟO�}?�=�00u����Ν�a0�}�����b**cV�Ӥiq]Ŷ8�Z���=$;swݿ|~��"��/�������0D�I��qT;�`��g��e���ù���Sav���-�y��GPݛ����;9�O>���FLf2�i����&; n5�">sw��|>�� ���;զ}/����h�mb�����Tl�U��_m1ѷ�k��=��x�.=$0d�(#%T�LYpެ߻xuǨ��ܺv/6�~��}�"����8�e��x�����>��D��M�2k>����xq�f#�E�{��ܠL�gI�x}��G��5>����u���"�:��g%�$����Q-�Uc�~Ϸxu��0A�D�yLzO��Oe�A� ������;�OÈ�O���'����|�v�f2����󺭼���@͏Y� 7]�Gl�d��*���e�h̅?Yc`d-�VE���,#Tb{?L8ҁXJh@ ��j:۷%u��v�k�t�u�iT�mݸ�^c�0^M��97D]��<a��j��P����wtu҇	��˷4]:;!��.
$f;M׼�������Tu2�lb"7�"? @�^��0�����xu�W�ݷG�@��/I�A��O<���~d
�}_]��t��� |�zO|�"B�{�L�1�0>�V��U��7���"5�#�GvZl�zp�����}��R��^��3 ��;��xu��F����v=���fc�c�s��n¿�n�����G�H���n���]�=c�)[b�˷/c!��<��7��|�qۨ�">y?g�4�1}1[Q$� �L�zO��Ho����*����ڊ��ʠ�\^�ۑu���ob]{M��:���G�Ay�����P>4c�L2�WT�暴p��l"$�O��Ξ�W'�w_Wt�;��P��N�67a�}[���9�Y0ӓ{���?oмF�f����H����"f='+� ����ﷇT�ԉ�wI��;�Տb�w��EI�ʙa� �����_S�َ4<��b{>������}V���1�F���D�d�3�+,Yix��f��$�WZ�gܹ���V��ԉ�+Z�at����tr��&W°�)�h�X�n˧&�+����]'��E���G�E�#����)�ֵ}�^�ޙ7C{����y�/_44{��|�z{5�����7�h<�.��e(�����_�f�{�bħ�c���㝸Y���&�8ٍ̣^D\���n��j�����.�>�qz��H�ej��T��"gu�҆F�-5������o�Gi�.�,|���N�m"L=^�.�]�g���^k�^kwq����`9�Rt��h�L�!vF�/oړ����8���ݹ��.`R,�k/�H����{��@{�W�}٩#b�s� �5��z9�ŗm��v
E�ɭXo."mab�Tk,f�G�MN��TA�[{{�xA �O�����
�a�x���]�Q���)�ud�J�C@;�B��2 5 h�0�!%ܩĮB��J\���܍EpHGIEE#HP'�08�8т�:�Z��ɧ�Cƫ1��@P)E�}�q��w�TzO�1�!�0D��6�����	���7���;��(��o��z��l"f2}`@"f����^{��y;��Ù���Ј��(�f-��ځ�dji���xˠ�m=���)�}w��,� �/I�"w~����~p>���&LG�7���V���x�?yǧ*�k;�g^o_���@'������8���8̏Q��$L��"6�}��ןh��|ߥ�>�:Ʒe��g�����W=���A �}�������l�x|:2���}���$)s�=[�T�W\�\� ����q��fO��Ǥ��[��������|;�����>���]Tu�	�%��uH�K��'�VՈ)q]>�� �����vo|>g�>��?Wc���'!�kvZl�����6��q D�q���~q�?��&[�!א��}sS�� ���Y�q��V|�q�Ǚ��"<D�.W�ڼ>� L��0!���;�����=Cn~E�C����zH`�f2e�"�Ő�WX�����u��f3�Ax����J~�|�*�&�Ւ~ق�LA(�5⩋6��&+8����X����0#
��	nH�8�v��+��0�D���lc�n�7[h��	ޓ��k�7m����G�E`��b+$���,���2�U��%n&^!���1#1�Ds��s�;]��xh���i��M�������#3MV��W|����⫷&�>����Ag�B"f=%��?Od��`����ӹ�}���;���5��{�4Fd��\B�ۭq5>�犝�k�w׻�:��~"H1�1�(��z���b�� 0}3�����>��|H#�>��<�Mۺ�R;t�ｓ��#>�߸�?��G��d�3�|���彦'"� (27*d"�uB	�
o� @�#'�0&3,���g�5g���v͐z x׌��d���#��n�g���t<��� ��(͊��]��=�kV�&k =Y�~����?V��e}�p�~"������u
 e�ӧ�0 ���D�,��r�=;�|y�|~�-�CvV�?wsw�YͲ�b;	���w~�>��?�]��zn$	�`�0 .��3�1W�?v�}��q��3�,u�K���u���lI�3�ݶ Gm�B�k��i��,�`jC�7�������}��/���"O���@��G��#g�,S�6F�7������Դ���8<�T�G��6V��f`�T�����}�Pܡ��;5N�*���o;��įr`���U�[�g������DL�u�#���~��ǽ_Q�&��D��Vg����|~�D)b�w�, eǦDzH1�6��o�@�ݞ{�}\>��1���Hl8O~|�;����9$ttU�hCE;aNy���y�L阞U�ӟ}8�u��" ~���C3l]b{��=�ӽ�}��ޭ���� ����zIJ>��]ǭ�&��D��D��V {~ߞ�mp��<`��7l.��m=��O���Й��U��[���@ ���P����%�V]TM|���Ո;n�툁�̞��k�?B	�+\G`n���'*'.��Ϸ���}���}%x�f%�3��;�0����m��D%�V���ʽ7���Y�; #&3v�y���p��!w�L�F@�/��� fLy]Wr�3D��Wou����|x�x�ё,"%kr5������y߿z���G��a`�113�~���!�׬LL���U��χ| gו�L��.���" 2�.�v�>�}�_}�}��w�	� �|ϓ�Te�����;2M���S��gۚf)���}���n�z���.�>9�c��8��Tn�=����Oy��FևVzW�Y#X;�s���7B�pdT��E�&�m6�<r$��x2g�W�٨ovκ9([aE�6����]�M�]B�D�RB������Q�D/�w�߾?3����Ț,eY>2��&$q"o;�����^1=L�߿,���þ�M� �}n2.y���A�3�@f������}��>��A��#��11F�;���θ��nV%���ϻ���}��GjI�����2 �|�[{ʅ��_�{>�8wހM�!�NC����9�|����٘��%��@�Z��i��}�+�s�f����w�ɺ��A�Y��f�3G����������Ш�4�C�8�Z�'t�싼,�;�b9[���x����o�G���~>��_Ń8��g�B� 8�>N��F�O]�Ǉ}���)2T��Ƨs��F��8�7��}￹����??�'a�M�Ӽ6�j��+2ѹ�!�ݫ��:������(��˺�gu�H�K0#�Bh�0�BjK�S��_�&��i�(ǈDkܟ���?'|��ݍ��"d���>�ٙ�_�]w����*f��þ�O�AB8����é��P^11k��pU�ˡT%����=j���Α�E�#��dF���*��ʵ8��^�}��}j~�q�c��]��$u�K3�������q�����u7eAf.<��>��]�M���ﻇ�?2 �S!ϝ=��DH�}w�iże�l��L������ߚk�"�=�滛�Ga���/O���@,��27A�?wh�#�w����xqg��G�w�Y��dQ��4}<��r��S�O�����#�	��1��19����}���0G)G��U�}��?8`���\g�ҩ��_}'F�u2f�3%�*��)W�qn��W�oᥘ�|�Yg��!����߿o�	�� ϓ�n�߷	T�ه�5Ud`Fݪ�A�R��a��>��2+^���8w��n!�����fJ�	�w��<��jl��[����?a�� Uů�dAd|�����Z���w݇�� �,�� ���/�m�Kk���g�6{�þ�~"��;+�}c @!��2��>�����v�q�&Փ��?Q�>���T}e�ST}i���k0��E_���E��Њ�{�.���9�8���>g�Ϟ�9w�;��� ����Tk$���K��q0���'HQGQ������|I���;�����T��PA}�5�t���<�K�-�~��'S��٧��L����dh� K���؝���S�&�x�[aχzΉ��Ѡ;�x�t��׺�/���>���x_�@���@ �/��A_��	b������|�ف�� ��A�D�8p�~::�Ѡ>���/�y/���}�( �O�'�?�����(�����N�iP��!�������������jD�������ʒ�������⓬y>���c�|	y��riE����f�V��|��E\�Sk��߰� ��"(�qT!���,�+�4|�N��8˸~{;�b�/�r'3@g�����>�}����Q��6��"/�����~P��C��;�@��S�_2���l����������*/ ��hX~����'����S����ه�#���4��1z(~_V|���Ϸ��Wz)���}���>��׊�#��{����C�|W�!DPOR{�%�=��ұ/�~'��z���G��nD�I�b�b� �-��(�����ʄu#��bQ�zh]�þ��S�0D�8S�'�Q�9V�����t^�X��Q<����.�'@�=g�9N���5��$s��p`����M)�&jA�C0|��������PA|��>����_`�-��{�?5�#��~j{I��?�#���������<��M������/�}��� }�{��I��ރ�������/@7�?�`�/����z�K�P��L� ����/��./�p�Kutc����~�>�d<��}��?g��NN�/(1�����Ȉ�݇����O��u�?<	~��믿�~Ӯ����7�^_P\(�����P�!�!Ǽ{=�h�3ݳ��G��0�3�|�����_:}<篩���C�O����V ���>f���A:�'���a�=O_o�� "��{��$!�������x�\C�!�M|��k��<�"P���O���G��ܑN$3��� 