BZh91AY&SYu��U��_�`pc����ߠ����bC~�      �J�	D}Q��j�UTQ�-`٪زՠ�h�l��)�SZ����([em��ZQ-�TP����j؛4 >�[�T�XR�P�[kkfd�� �YU%�ѓTѬ���Z�1�JQF�%�UH٭�VjkZ���m��*��6��Sa��P�wym�,�Y���[�Ѳ��1���8�Ͷ�V�bw�y�)lm5����W�Ql�kYf��ѭ��ZڬZ���,��%UR�Y�m��m�fMmf-f�Wn�ƍUmX3� 2���`�QWN������õ�:+Kf�5�j��Zuv��4QFژ�nu���Alnm�ؠ��5��&Twc�DͲ�a  �Q��� ����^���{�P�z�]�݋۠��{��hVZN]���=�o�����}��j�JR�:�9/xC�����{޽)B����Z�h�U; �l���(�  ;3���졥>j_p�(;{/x�O����o�w�>]�����|�@��Ҷ۾����|���_m�����z4Ӿw��}���@��@>��핚��m���gbHTX�>  ;����J>���wʂ�T�f�W�/{a�N�}�A�5l<��}�B�^�SN�O����w�ﯣ�+OC��r��v��;ӽ �=z�ކ��R�B���Q���Rjڙ4n �y�t }U����Mw`�C�4�;�:i@n��0��R��uJ�f�����*��z�n��JX� ��n�%liN�U-3)�2YB�V[-��� o�� 5/�ծ�t��)[.�=i��*�mΔ�=����S������;g^Sm����^��o{[�@7�@=�m�*��W�M�ښW�h:�-X����E����� 7���}Js�۝(ٚj�t���4��]=(4���xo�Қ}�[��B�5^�84 �\u@']pt ��@����kYl���l�j@i� ^ zVN�Q�4vk0 :-�ܪ}Ay�� ;��tcGC]Q�@:��(	�( ��u�� n�3EZ�2��w��K-�Zj�7  3��44�ӟ@�y����s���$��  ��{p�Z,㵭 ��࣠�5ej�r%�Kf(([4(֭�j�� �����	r �s�C@Ww-��� 
;�k�G�z��@����] �u\(g��ڽs�R�|  �          �*J�F       �{M�)*��&� �44��2)��ꪧ� �    *�	*��0!� �0�i��*����oI4ɠт2b�S#��jH��4�Rz�jz��i�d����O�G��A_'�_*������n�����s��2�����q���;���6m�����f6m�c6���6m���6m�ý�������������������?��mo�9U��l���m��e��n�����oo���;C��hv�X�gkgi�[;[;ZY�A��n#&õ�n�f�c�����`�m��f��ݭ�;F۴ͻF����h�a��c��gkm�km�k6ݭ���n��8��l�3�ͻY����;X�;[�Xgk�����v��h�v���kf�6%�۵�v�;F�;X�h�a��ݢL�;[1�l;F�h�v�;M��6�;[gn�a�a�[m�Y�k�1�m�k`�c8��чkm�K6ݬ�ͻX�c��v����n�ݬ4�Ѷ�m��`v�;[m���6�6���,Ѷ�l���v�m��;F۴�v��7hô���cn�6�l�c���@v�c���;M��m����;[f��F۴�v��hgh�6ݬõ�n�۴�n�a�ٷhm�`�m�km�ht�7hm��f�f۵�v��i��6۴�v�:M���ql۴a�َ�1�`�3�����c7hٝ,�v�7i��;M���t���v�ݦ�i�;Y��6ݣ��n�aŰv��v�;Y��l�h���f;Cn� ;F�h��;M���;X����1-���n�l�1�Xn��v���ͳ��;M�[gkv��n'hݦ'Ni������iv��m��i�M��i���%���m���ݡ���gkn�sn�v��m��i�Y�۵�h�v������v��v��v��v��I����;Y���ݡ���v���;p�۵�k��C����Gi�C���GI�M�n�v����6�gh�K;X�6v�n;sgi�[v��7j[v���kn�v�k;[v��i���v�i�[v���kI�u�������w����|�o?������l~���W�N��8n�į.��v�t���F���]2�5��a����9!(0*R�p�ٖ�i�� ���lO�t�wBũ���GG �e���[w6)�M��sq�̼�����(�b�F&(��5
��ka���D�c�6aԕ�`'t�n	�+*%�����-��5m��n�'F���!�;��f"�B1lu��(R��j�
�sd�l�mV�+���ek͢+���v�"�H�4��k.��t��jl�����)���Rr���)5�Զl;g~�ng�f����VC��PU������sX��}5�VRT����r�M*�s6��-J��t�j�(K�(�`V�J�"�m��@V��f�Ch�.��YvsUٌ�cϦ��w(!�#0�3�J�1�3�?�Zj�
����D�yl+́��]��zm�aPhJ��s�`Z�Q֫6к�������@��׹���e�&�������TǸ���]��@Ӳ���ۑ�o�pN��7�<�Ʊ�c���:	��[�tN7cD�^:#B:��)�v�v���0	V���e�<���ڷ�]�9i>۬%C\�Gmy�j�!�xۏv<H쫇/.j�����b�uQ��X\�,�Ӯ�6,*ӌKӺ�4���a�M���d�n�%��׍T��j�Ǥ̨enIo"�捄���K``[�Y�˭�\���w[J�,m��64�G�5R�՝�]�n�ض+yV��4V�" �6d(B�;h�{�;{�=�3`�%C���9.|�Em��BY�����ܖ#u6�5R���n�]�*��Ύ��ˋ�)���i;Gl����"�Qi��b���	�n�d"�
�h&d���Z�i��C&�̃
l�S497uͲ����!�vf��W��ٳs6՚ʓF?�"vr8F��+n؎al,�em3���`��������̳.#��S`�Y�	a6J�p�&q��l��un�	1�^pH�RR���α�<u2<��U&2�1�r�ƞ��,th����^�01M�v�úX@\��NL6���Te��Ӗq��34�]9�)K!X�n$�b♑��F�AL�B���axMo��B1��R�p�,b���;daJhX��J˧1��9��f���`��Ւ��T����t��;W*��jb$�
��(�X��Ci�n��ҭf�M��/M�{�VDK	G�5U�P5YI�!Y���-���ن(�^"�i��A���-�h �5��V"��r�����ڴ�W���N!�6VA�6j�Kך� �7dj3f�w�Z�{�c!���)@A�&���+���(-�EM�P�ޭY���f�Ų��i���������43N^��G#G!Nj (E M���h���!�]�͡+bxC�6)��I3*��7[�wA�4�Ch�p�wWK�Z*�13�yJ���X�t:�nsx�/Z��Vp	��\ذ�`c��d�â�93%Y�9�����35*Ajݵ��Ś&T�e�m# z�%�����.�0��'��_e�iVE��Z�ףgڲ�2b���W�����7P��0\򖁂y�c#�GQ*�y[��ջ��ï6(`/l����ƒ��@<���-��pi1n�5a3��yJЫel�J3K�P�^���70�L�Ӗ�T��x����d�[*˗M�v5^nn�"*eK? ٹP[�{�1���͚���LܔF�ڹ�N9�����픾Iv�,���M[v�/�0�u�38"oi7�Eh�D��Q��݁ASZ�Ld�Y��enY�f"�JML�co mG[�a���Vj�6�&����ֶ��4�N� �Z��bЙ�U�ke*D-RQP�PU���m��C%;?`�+-U��c�x�~f�i���X��Xh��|lu�a�Z�M�����+b���7s�ɻ���e;ZB&����ř4.�����!��N�9oo$�V"�y;�x�hM�	���g�an��[�h-*j&�ٵ�d5��){%���(e����f+[j�`�-��.(��! ��@�.X�c���Ej�;ZQ붆���,�GF��	58n�K�S3 O]^ڲB�F�7y]݀*��˯Z���|n��u��u��9c%�RP��7�������ʳch�C@�=��+u1�cV3]��e��� �S�71�a��zJM��r�����feH�U�˔f�E�T�Y���Mڷ���ʱ&̼m���5m���卧��1�y��6�E�	˴����*��5�kFV�Z[�V4EvrhS�ydh�Fļf�tJE�r�qd���sF����S1�j	��li�v�"�5�fb)�Y�j�f�S0�yKu��/.A��tr�2FwM�Ў��c���S�h�8�1��f�41��i%Z��o]S2���$E�2�dc��f%�6lhH�r������m1�cv/Vj��
d�F�,�)�2��*�lfh��G�e�Bn� �-4�1��.�]^n<�5��:P�Abjw䚙.�P�`�S*�����-�a�1G[�(� ����op^L�N=}��;\4�b��:d�<<)=��!¡b�T���j��0[)�RUCb�F�j���"���A���e��̸�jc.�n�E ��1���=v�0�
:�M��UIfL�a��{}�Y��&m�I4Z�%�3*�-�e�;Gkr� ��#`dݦ�{D,�V=�ٴ��2*�st[�96$��6�ҥ ������U�Ԭ��iM�,Y�6s���t���\Y}}ԗ
�U�u�݀^.Ԡ�7M�;�L����sf�z���>9�Fh�8]�q~h��øj�`�XY���nՈB�����n�ɗ��pG{e%�i����1X�yJ�
��E����i�wкڕ��X��κ�mQ�ll��6]�V������ �y�V�0���B�+h�/.�-��׺1��N�͍.A+F�N�M�U��oPʾ]aR����bΣ5�6`T�b�е�J	��Q�2�!^m��D���4�k!����ts&<��}��'Z/*e;��D�7,f�t	xŸ��V�s�v�l0#�Cq���񱺲����c2Q��ec*`������=�T��pU�9J���[�]�1T��]�%l4)��䣷oZz�^��^�	�t�2]ֳRP8+PFh��v����a	͒�#{.,[���uCT���2����*c6��L�Q�YdXPR�+D�t�Je��Y(�6]���7wE���U��M��V~c6%!�E9,	"0ҝR�=Ԃ����5&h��vڻ�0�)�B�3Yiطh2h�3M6aٰl��+G�!ulpg�]�m[o[m�6�#j�	2�mK@��^PM���jS���bSTm<U��'0mCg)�
�NRTUgtb���N�-8�E	�5j֝M�����@�M2o�G��W3ɹcu����SEP4n�5b���%fm��I�8�)֓Z��^m�d#0�8�0�Қ��Oܫ�`b.�;��j3��{��Z����Ʈ���ua��m=	�u�*��*�K�PS����)*րj,��������W�x�P{���� �kf�+.�/!X�bZ�����f	�T2�h�F�e�X���m^H2�1h܌m�u�.md��.����i�-� �M�Zϕ@~��3�7F�'g)G4�6[O�xS@AO\u��1a��jR�lK���֖L_c�Q���B��V0v��NDӲ�ܸE�#B�b�p�
�"��E����<?^˰�ۆ���ӽ��5��, jeޱ����c*Er�Y4����w"[JG%81+�+�����,�d��]��*Ԧ����I���̮��#cT����Wa�9M#�m��j5lP����N�!ڸ��/.<�A����K�<��Ղ!����#AIpi3B f�?h�(A*m����)�P8�i�Ǒ`i���K��cǜ��+���vo�8Ef�XAG�[��;�U&��&V��eVԷ�C�L��O��T �����ܶʍT�4��z�`��r��Q8h�;5�Q�N�&�f%9wh[�k�Uէu��b.�%��(�`;��]Xya�NV]�Z�3u����j�Vm*k^�n,�H�,Y�:a�9�Y&	*f���+5"4ky�4(lĥ������R�f�32�e�ܛ��6�I��" �͔�V#0�]�b΢�F����\�9G%`
�l�jZx�hTRԭ[����ts�]@�Ws� �7 ���Y
�i!�P��@󐵮�]�Q*���{�Z�ꁣ�?)b<DuN�����ʲ���u���Y	��0f���f����:"�U)�We4�L6-�*<ҕL��^T���ڼ�q���sw ��(\���R��J�0��b�����h:�*��X��f�2X�`A�hV��Ԇt����!`�ŜYN��U��_.�m�z���h�=�
�sF�E���d�m�ma6�Z�	݅P�Pf�tPF�2̺J��յ��e� 5-��M���Q�@�_b�r�	�&|c\�5*��O���Jt^ṍ3�T��-5��Q�����sr�@b�.�)g퀋65�;c%Un�Үē�n�t*���ķ`t�;-��퇌��H�(�B�l
����P�уp5�̣���ٳ#���Z���k��R����j���53e�%��+��2��2�e����Y,n�V�S-�RS��Ǫ^ �ٔ�
bh���hVXwON�ʶn�4'����R�;2�`yЪA����|�M�t�w�@�[4�b^i:��ѽ�M�2�T��8\�0�i�fM�G�4k�ƵԬ��;�6�ɩ-ɐ7F���JX�)�6���ܥ��d�̺J���դ��Ee)a��*��j���-nE@�t�鬤Յ	m���՜D�yG#�ڦM�@K3m�����RS� �l��ٛEj��a5�Ḟ�[Gt�3T,*���6>�	j�0�J44�S(	�'t��3�.)/"l�v��#$�T/4��Զm
,�G���J�45�̼��X'C������1�� f�1����.&6�H�f���-D|BSd�C^U�oi�i[9���,u���$�2��P���<�;��گ:�S�P`Si �����<"���.BN�5�\�?=X.E�
�d�)�4�Ө���T��o-�E�t�ܰ�zsy����\�7�q	�c��sR���٧/7��c�A9t�K�S鵁 *C�Fk�1=�@�&��m�*F�v��	ӵxÍ��&�*E��Ii<csVX �t�ǄV]������d;�J���f��M���� �2�?�^�ɭٌ�$p4r�?\̒,L
��v���Das.�ӶSy�:�V��/i�\X׸�5��a7�pm�Rơ7e�6���C+K��.I�#�j��Yv�I���
���c�A�hQkn�á��Tڒ�kh`j:wH-p��6m͊��h�85M�e\��5F�
p�XT��d9PVb���L�ZH��n6^�KOݵ{rܼ�S�NH�U��i��j���юEc)���;�h:*��A�oJM�gp�����@7��`��c���Mk(��yW��ة����h����l�v��[��n�z 	�*V���Tۆ��ɹ�&��&�vso���C+ڛ�+M�xpa��͊m���-bkV��#A	B�#���̬�5=�F�����P[V�sD���q�� �b��Uj�T@m2嘭rU ��R����9M�focl�[�D� vCyt��R��v��%ї��AV�%0�vQi�Ό�8�^��Ԥ&�:�U����P�u��Q�P��Q��k�32x2c��4��-]�nAu���vf���C`mƆ��t�%,��Vs`Z.�sr����yE5&�'34���v�6��S���� H@YF��2-���^^U��Vf�/�/;�XF��l�%*�j��0l�rE��%ϮcE�Բ��B�M�u)d3 �u�r���ɣwv�Abh�09$&Ć��j�J��)2�2f�ܩ�f���n�N�5J�ʢ�v�@m��p`����KR!��C5
V-�4[�ݸ�ˬo�*�Ձ�W������>M��jU�uv�޴�a@
J��Z�Ŕա��;SZsf�kY��i'e��۔Du�:ͫ�E�1yLc<y�N��U����ۊT�Q,ؐ���8�V�&��5ٽ
�jǲ��mU��ұ];E$f���Ĩb��W�:@Q�e9iiʺ:,�(�CgR8cà�$`S��ywl���KU��`��i?����вa����`녴�Кm�=�(��(�{e��R\m.�G�t���h�kr��AA�08w�o�Y�X���K9`�Nk�ݯ�S�W0�2��km�&�`Q
�6�x��sd�+x	���lwwCRv+m�@ �\`�	 Z�7K�ګ�2I�^˂J�t]ۛ��w�d��x-c����2em1SXe(�c���:8h�.lT6���bd�,����,�4�h�-���Uѩ_O�����OGN���㷷N��#�ӷ$�'n��;{v���=8���;{=�N8�Ǣzvzq�v��;q;q�N�;q����������N8��I�qۧ���;q����Ogo�g�O���{}zHt��N$����$�I$�G��ۧn:t�q����7n8v��Ӊ�N�#�n�����v���&�v�t��8�8�Ӊ۷gGGN��ӧn:go�=&�����;;}q��ѢD�#�$X�?�j����/�7���H���W�+`/��qf\��X�Z�<-��7EQۤ�q@�=4�a�!(W�������K�N]�b���h�F��:&Jl���g(D5+C+$ّn��A(Z
�9w����&
�f�Xӹ[P��(˱�����d�?�!FX���B�̭ɠZ.�! �>T��~�ߑy�����{9�OUE��~��/G!I�9���������L���E����e�
�ޅ��sQl��c8�ew#kDP�lm:����Fv�J<^�����u�*켃].m�Tb�Kn�r�l=7�,��}z6���r��؝���L��e%�U��`|_pH��bڧ�,^љ-�*ʂ���:y�4�2��	g;u7G��mު��e�gEʱ=���8�)M6v��o7vM����[�j���i�)�u�2ḋ�����@e!n ��řnK �a�|���1�����ǳ+޸LIL��计��oz��j�Md�o-�n7j#(\,ջ����s�,��*��3���.J�2��2��=fKT��%ڝ���	��}-�s��_�;�d囶��SN�Փlj�`Ѹ)�V*�Y���0wgV�ԅٝAD���9RM�Pe7Z�db}#�3�ρ[.j�H�^	��W�1����\J�K
��N��+��\�d�lgB]N;�V� ���^��S��&ު�[�mf���#A"���Ma$�{��wy���joj��ρiӖ�k_XlbKA(�ʔ��,��}���\7)i�K:i�]]{�Ep3�a����˷2�5Z�i��v(]�����x��6u_F.�_s��-^4��F��u+�Y�!�;���u�{v�n������k��Z�v����6�sP�v	��>VUĬ��|{s�����45_rU�(���V�k��r �_}J�d)�-�m�
�P#{�t3��	1�$�y[1���\1R�JGMŉL����M�U���AF,�Ƒ���d$�}"���5�b��
=z���8*E��:�f��K/�P�:�ʓ0�ks[��K����F>�l�e�ʒ<&������q�33-I�X-��;�1Cu�]C���2I�L��R�B@�5�����wtOS���e䘶�s��5ΰ.����i����ڳO�tYOz����^Υbh;���-ǹJ��g$��=j�r�ꥸhb��(}����:�$��s��g
�-S��h�~}r���G��F�,�F��h"�m�%�X��J��6VN.�n��ؒ�:{WX�ŉNa	�8ζFv<�Q1-���W��ƏB+����õ��bڳ,̅��K/�h������Eu��9�ӡ�����+,�,vr���m�hƣ��W��u��6軻9��v��t��s�`wf��+�|�.��E|���	�ǘ�	Yxaݼ���WӺX�>��c/R������/��\+��O�v��Uқ�����[8�+1�c-:ܹ���Lלt��Z�Nΰ��ܬ�q�s����L�����͛u HAc(',wN)��~���j1j��̸/{���tܭ�;/��+������b��M��;-���j��_a��A���?m\�C���nv�H�Ć�+�E����r,�u�G4j<Ct�$��V��ϯoӀ�R=�D�Q�@j���V��Uuf�h��ZΗ�ho��Ge0Y�N�ز�-1�^L�8�H�\���3��o)eu���Z',6B�:�<��g4��2���x�{�n��L ��@ST�Q�u}�[QuC��n�ˊ�ӠƸ��r-�-��s��m2�ܼ��(��t���"V �l��eM�r�9v�+p;����\�&��c_q娄���f[�V��C6t�J�[�Mz_t[rF�8��h7b쎗�e�����K ���m�j�u�޸�U�ܠ��X�����[mҘ����P���>J|�7�j�]����)/��<���Wֻ��2"ե�6t�t���8	[���&��ϯ���� �E�:��J�S���C�f�#7�\�2&�Ή��X>;xN�|�\�PMڱ��N^q:�3�A%�6��;���4��N�:�3E�y]Y�9GG]�(ܷJ�[�v�ѕ�,ӵ�t��ڗ��c�^�6*�a���0��v�M;\��itQ��	����CׁXۼ�O$ZçP��.^�*Ѩڑ�Fӄ]]�N�h]8>��3�}e�87a똷��*#-R��.��OmHi�`8�ˁ��+qYg�X��.�[&��/.D�U�o�1�nW(�v
�Ͷ0�oK��mt�#�Ψi�h�sK��7;�,������z�nε��F���x|�ݢt����K���j�ڈ7f��P��y>�� vG�ͧX�)������}Ҵ��/i��{��W��]f'T�qnh��*�fVu�Cg\;���p�{M^��\�i܎�Y��j���%�(+�L˭Yz�k$�}z��9'w@�I�JO�$70	�i/;��A�;(>����0z�ۏ:��Ѯ��3e�\��|M����1`�i�An_�a���;�C0CRD��VnH�wn[.��ܑ��Ļ�#Ȥ�r!��V��C��) V��k�TԅZ�7jȢ�fg*/��%�-e�(��D*,�A�xw�� ��ٛ����\�C����L�#�o-a�3!�3h�p�]6�y���]�!�<E2��n-c���ϩR}f�f��R�P\T�#2������|~�����[.7k)L�}D\OFֈm�l����ra�V_K���*�}i�6��󨽚�[DK��b�a����"���������EBW��"�Z\Ǒ��J��j�I�C��B�k��7En]8���Tz˗q�B���ύaO��]G�PqJ�����G �N�tH�BAH:���ܭ|Ƽ鯠7m>EV(�qW ��OJ�W҂�������Z �ب8ArI����`��.�q�]'�q�7­9:�NEwV��B,�եn 3�	(�.L��y-4A�Vbz g#�DKf��� ��c����\ȋ2`9O��H�hzt;�ڂ�K,6���v���yr@ᳺ�q�g4�+2�]�2�z��M�r�Yo{(���S�y϶�m��iH�E$��M)�	;�Y��t���º���f�����|�т�!<���|���y�P�ܔ����޽jU���fk/ �y]|�x�]�3�R�gԁ���ɸF��4V��oͩC��Pۥ,�oF
��1F�����Q����T�rUս�b.ˣ�R��%��R�2�,�`V �i���
��S��ZKq�V Z�މ����0e�;�`��R�����Fm7���ʕ���x��T��s��s�fU��æ���[�\�J���d��GKλ�ٮm���bJ8=!�@�4Z�$4n&v�5}i�`u���װ�l�O��w�����\+q�2�^���{��6eac&��.���G�3z�f]Iv���bn;X#�R�Y+Ȳ}� kF��
�z3njK*1���X��nU�zˮl�
p|_}�o�B-�xq�f�9g���ɍ���E���=�������N�e� d��<vQ�Aw��������V9Әt�J�榵R�N%7�P�nĈgL�A����7�q)˝����Gt�j��X��8����\�&V��+ul����(8]�/d���J����΃�U�����rNP�D���8�")-���@�C��9�I�f����::t{]V���#V���u��\-̄��J�w�5Jz��dtr��³-��̹������\��]�J�M�W-,��с�34I��%h�vŽ��[Y��|�a���U<!���p��GRǢfQvX�Cz˥��܂��d;��uu^;�H�y�X�,�
E����gf�9R�Pl���Ʋ��Jf�iZ�2��E�V�h
E���u2��B�	H���݃�G�
p	�~�&�c )�Hn]%�wK/GZh��[y�w��Iy��>4�3+ҨP�*�/�m)��zM�+���C�7X���ʍ�O`�A,�f	�v�4�{������V���1�ZMqriO��uڮ�l���G%[�5�,���ӥ�M����A��[�ln[y�.л��mA�k���U��M��2� �FGZpδ2�P�d��V?�٤�Q��h˾���wS�Nc`N���ӓ�A�(]�%�a7z0��AZ��5bi��V�qD��:5}�è�M����=}�l���:{lS�j�r�ǵ��wt�M=)�4K��ز��by�u�%_O�I+�*�Ǉzb
��b����+Z�h�8��Fk�{;f�@���In�ˣ�i��s�{7�Y�i Sq�W��]��Y��͸��'j�ST�˥�
�T�R\��ѷ�:��jH�f�(��n����U�5�e)�d��n���<�K�.���30i]�!'���y����Һ�d�!h��KP드�/�ne�>ݡ�FZ�ںV�X3�Wrx�\N��oSb*Y����S��G�[�x����7{�}Iu�s\�[����m����<-�� ;CH��n�ݹ(�{��*t���ܗ$��R�xNe�Պ�,��'ݓ*=n���ټ��y�O=:�y��ǂV1�V�Vݒ��mX�2&±��蛉�7l;η�K��X3�:E�݊m�YK��Jjt��
JW�]�o#"���h�sxЖ�x���J��3��XUن�N��I��rZy�K�� �/Fe-W^����+�9(T}��j�H�nz[)泙������n�t�y6><OB,qfoM3�iKc��b]c���v�P�/(GL�;�� ��3��0p��"���l���ڮ4�&ro,V#]��� N�JI�F���w\�{gmthX�ƙ�(s�9 �䌕۴����[��e�ٖ�+)��Zs���6�od�, (`�hkuÚ�U�1�a�$:Z�md��6��"��fl�4��v��<i���0��n��e0�(���s��Ԭ�2� �'���vR䕲u)��X�)�������S{z��T��[���h��yP��m�չ�0؏$w������tt�"{"�i��&E���[�/�N(�zF�;�����̭�����R�)˞�&�
�]�k�i��D��5��\ٚ�1����vm7l��r�M{p�46�8oR�ҹZ����@��n�i�٩ݛ��F�]v���xq��kD"JRӻ�*�4������S&4X����5� s*��k�NwNw�;)tt�S�R�e�|��(��WH�k�*�^��X�g�VnɐPꏝ��Ú�b��]ٽ���3t����2M����.��F�]��j��DVi����m���M�1�oKwAM���%&0��V*ۚjk�Q�k9Y��.��$U;6X�{v�=#c��U�mL��ɫ�������q���k5�tl�5�JC��â�3��NWou�˂�_U�n �s�AZi�M�X1	Y���E���᎗&��Ph��\�X	d���mSh���5d���N�ȹ�]\���`�"�+*���WʘyFcB�!�'�w+��_p�:T��d�*N���P	��SngL��!�"xl9\�\��-��z\��PNCoC/��Y��L�o��͗6:|VA�	����WZ�y�-5�P�T�d��:Q�D�x��V묬�(l��B�ľ���?g=��|�%Ssh�}����t3;���n��V��_	b�7W���F����iW �˰�5�%ݗ���Đ;���v�BU �z��]ձ���{) F���#դk�d���,lӁ��#em���fC՟��.�d�	�i8�2Q�����|�s�+UW03ӫ9��&���%ɴ�EQi+3�󿈃�y�����υ���ιZ��p�nc���.�N�ݸ�R�Y	���K���]Kt����xp�w��syb%�>L��J�P�"�/Q{����("�L��)viy�)�1���ygy�ڗb0n�q�y�D�6�T-t�'�$����.�������N��C�ДXz-\(�K��WZuַ��%+�F�V:���N]�F��a<o 3J{��\8��ܛ/B��j	�3�3�Z�=n�p��sOY@�5������j�����m庎��h�� �J�`��;�X9�<��;����j�Ř�&�*J*�:�R����5��������س^ۧJ������N�<��,[>K���nu�����7����c�`�Ҷ_��W�mᙈ��פ�9Y:i�Y,�@沉�q�uK#42ap&v�`ޏ,K����\_�hmt���Du��.Q��ձA��lڰx����:��K�r�6I����E1�օ,�؛�n&���Vt��E�0d֮մ��"b"H-�N�� ym=��1��ڽs�7�6f1�p�t�Ή������$ȫ��Sa=|����ֳ[ύe;y�K%���$�Rݦ��uk8�����"W;�<c{ze�j�gM�7M�곈X}}�l/)�v��ǂ���%�����B����'%[2�[2qڻ����@�'j�������VN����|�Df�Wu87o%+��&!��N�u��y��,�ߍ3;xZ�Y�H��T�g#z�cʵ4M�:�e�m�u��U���RL�$��v�%��Q�l�%l�${񓤝Eɵ$�d�t�4L�I'(�I8څN�WQ�gMNb�g3s7JIz��cy���Q�Xt�q�܊��]��Z��d�W ����e�;�I$�I$�I$�I$�I$�I!�� �
f�)lݑ_il+L��΀Գw�nc�D�Ђ@N��K`\2�(�!�a���t��n��)�UL��m�)T��H�	���?9O��2r�N����A&�BH��Ji5
֨�f�F��<s����aP(���F�%�|��}ﾾu�xٙ�/�Ͷ��;����}�����,��fm����������@�U��}�TYsR<$1^�{�ޏ�J�O.�J�>��0<R�B�m��W�B����}5�t��u8Ct�V9���c�^ɺz� Gp��y`L]�H%�wm�׸����Yנ]|�Ħr�4q�4�b�H+�jC�{�uu䖯�δ-o8��P-fa��,�(��>�a�r��uh�D�
��uZCd�����HXx�: ��8Y[��D�+}�gs���r'��ұ��l̮��_S�G�9��s��Q�+��;.��ب��O+P�����NW�ү{��Q����j��ܙZs�VaR�p����m�6{����NӾ��Λs(
ꋑ��k�7L w s��!��ߦ�;�&���a`s�}�̾���KuS�f[��\�ۘ�P6�7"� �ze��E��_Q�
;5��a<��6:��%̽�Y��!��0��5��r7��ռ�Ʊ�*��c��J��5
��G�6R�$l��Q׼(f�\M��.�.+���J�� 8�YO:�^�Ǖ��o�Y�j�Qƒ2����*��I؈�x+K�S�Yѽsl�5��!ᆂɂ���.;�289�Gn�&U����v$��Cr��ݣ{S�3��-�kJx���6^�������8U�!d���8�7R沶Y-:�h��ʩU��+iWWW(p�Ä8p���p�Çx���x��Ǐ<x�<x���ǧ�8H�Ç8p�Å8p�Ç[E�ӍrMO��E���E�x�p%�R����
�w|w�U������H(PЋ�q�l��fIa;:�N̡����u��Rm˙ ��F�"m�2m5K���
��m����2Q��Z����u�j�\��kg�̺����\�9�:�0�>d�v<��}������mС�VQ���6D��^'��3o-��%8�*|ԇ7s]��PC�Ƥ���K)��=C��ˮ�8V�u�jXpj�Ǥ���9s+ve�{g���BG+C+�]�uIz+[i�O{�|�F����g\W���aԣ0�/%=p���}+��y$˖v�'���0S�1;����]v�TT��3J��հ}}>�6����70�=�4>w�"(k�)�խ5k����Bb{�fQ�,�R�-�76(�+�}pI��$*����$�Ct�4�1���L-�"4F�nu� s���ZK�c�-���˓��eh�	�v%^�P������C�vz�s�����M"�;j��Ӷ;'����f��d�u�XZ%��>�j�Z�\v����k�:�	'�EN��7�b1��3t�x�W�ej8-g&Ρ0T�|�1+r�ҰS���5���}6���Q���:�>߯���@�����:����,�;P���I������Ƿ�:x��Ǐ�8H�Ç8p�Å8p�Çx������Ǐ<}x�Ǐ<x���J�+*T�U*T�]R�u;�f1����kOcThN�Lk�.n��7���*J�;1f'Ԓ,�G�]�(�ܢS�T�7�����3I��z�զ�oo�5�%m��᧍!f'ӱ��j'�!�)f�x�o�g��.�{
�X�ak���;�����tuL?�㽥��S҂�.�<Z훇��U�7�ʚOPK���T�͕qa�id��(�ھ8�e�8"T�j�ҡW��o,gse>7`���C5��͊7��۩D�8��GMN��oh���.t��o��uֆ��B,�X��%�]��Ul]�qiE�@y���Z(�K_�;딅O�e�ۋ9�o��N	��Vm�ۼ#���:�J|��ʾ�'��xӐ�N��v��֪ݱ�Sv5]�F�(r���͝ѧ�)!��rw[ק�@��S���vV3YW*`l���Z(w&��`g٧`��M��VH�Js��jQu�J���cx;R��Z�z��[�i�,5[-򮺺m��DE�嚱=�`�ivQYD�T�%�E���a1]��\\�=NdAۖ�������.h,����u�@�t:�#m��콮\���W+�%}����޺�,�V�1ڑ��n���mޙ �F^LO��z@.�"��2���� �:VY��m���`h����G������
��v]A�擛�$���4!��R������+kǏ<}x�<x��Ǐ<q�Ǐ8p�Ç8p��G8p�Ç8x��Ǐo<x��Ǐ<<x��ǎ�����c�)3Z���� ����q0����a�U0P�Q�Y4D�ܧ�#ʛJ�Rx4�� 2E�F��왝��/�'O����m+��U:�r�K�Qo`e��կ��)�NP����I�%����q�u���ke;h�d�E�$^SWP�Kt�LA�ʣϑ��w��.��R��b�fm"v辬G�x㝜��+B;�/CO��{�+�+@ؓ���D&�c�J�� �Wd
h�r����B_d����v��9cSX�Zz]�cu�`2�|�vrK� �-UJ�z¦y�m6�����r���i�����H� �˂�F�fsw�
�c�W`R4�H�AO��R22j7��ox<�)q*R�v��W���.8U.�5(�;�6S���!y[�5WZ�v��ʰ�T��7���@�7������nغU��X�"�͙�si ��y�}�P�W`�T�
�B�I����7�U�.�)����T�[�_��VM��S�뒘�[5,����R�W;�ԂȨ�u�����F�F�OrC�8ޚ�3��r�O�����M{�@C��X��b��b�D�409(|�8�3��}�� �[N-o��#ұ�;1��W'�]�2�Eɨ!{|�`�ڲ�yJ^�¶�,I �޵�� �XG������g#ܶ���ޱPX4��@<thUJ�R�
�*T�R���Ǐ<x��Ǐ<x��Ǐ<�8p�c�8p�Ä�8p�Cǉ�Ǐ<x������Ǐ<z�>�%Ք3�s��tQUdaM-���w�>�7'm83���S��u>܃h �8��W˖v,���<XT1�ۥ�T��\�n��7����]ԟl;�4����V6.�jw�J�RLģ��˥b���/��P�����5`<�q�A�*���*
o�f��  �E�S�/�1�#���'��Y�	�D��%K`�4��ݏEP_4�o&��^�e3e��M��7pئ9��ZCU\���VQBk_�-n�����!��<�#!��U�:����J�mt����k����}����Ca�K�W��R;�� ɹ
V:�C;�ͣ�*���jc �n��Br�r[,b�םL�\7)�1�EYÅЭ�:/6c��Cm��9���gR�AK=m�S!r(�dF�����+�f�J�"�0��*�+qb��w�^l��Y>��b5�������i��r}բu��Qi�Ύt�C4��{^��o6]*�N-��:�;�T�u*�f'Yvwtt�N�n�s�ݹ��wdӈ�i��u���U��K�m]������V�ۺp_\��PΥ�m��VF�
�4aC�$��ɋ�p�Eh�j�ioǲ`�*kg��66�cBZ#$�R�8L���ڂ�J�:�����F5ȭN�X�F'ݻ�o�{u�+*�
���Fb`��1�[q]WW����l�B�d(q�T�bV(�1~-G('�N�ѽ�R=
�:2QfnMѫVuG9WP��%T�Um5P�A^�6�v�>�]nm<��Rvɨt��5r֐eW5�H5���VZd.Ү�[�3oHڄdV��7Q�.C��xL��v2R��/��#Ȕ:�T)v�Y2�a1�fu�t!�;5m�N���G�[�7��nVeaK%��V%���h�2���_h���ê9J����R��C�\�{�'v�r�c��sSw��[����p��@���a�.�����C� HŻ��[�Sx�=y\.�q������I��������� �C���8���L_�i�YKx,\�U�Ÿ7��wTsGe��@��j��SM3/���4˰bT��ݙ&a MGr�m������c*�Q7���.BA�Cc����W/�.lPqb��.m��od��m��&G��>�R���t��ȹκl�2�r��{�Z*|7'N�b�!����:�5��2�b�k2�u⇲�Ntt��_od��z�3�e�*Ķ�����ð�D��2���W�c���dKV��h^�K�p�ka̜���(=$#�eӽ3�8����S��Vj�Zg�jÏj��@�A@�5dS�co�v�>�Xy8��^�4��p>F�cJ7Z)�y���+K7&t�=B£��
���׬�z�c��(I��0+��*�4�%勔�W`N�1�
��a��TnN�"�D-9�[[N]K:����1A"�Iz(~�PC8n.����� �
�R�P�nV�����\�Mgϻ�%� n��.� M�Jn��3�;s�ї�[�k��v@Q��U�o;����4��2�w����q8�	k+t�	�Hw����u"��E^QI�
�y��fZ@1�\T�!�L5o1�^��)7byw�[/o��y�ΊN�i�]��Uӻ��6&1�]l��,\WC����.Kͺ�K(�XNb��E터~��a��( ��?�r��R~V�����f0�ѻ���κ�v�Q�e?��,P���j�ݷ�{r�1'�]IN�$��ͭck��Ћ�,��S�;<yM��wC��M�3��^�	kA�.�=2��[�' iˣ�36�8��oj'H���76����]��|�d��i��(�	[x[�`o[��7����0T�Y���� �� bed�v��s�s3-�n+��ʐN/���Zw^l�S�85���	��5cn�̣�ل�KPo�����=�O+P3u�K�ѩ�I�Ȳ�
�A��+���%6��>�5k�V�MF�L4+�jt�h<�+2��@2;GaO�'N�����0��oz�u�o(#B�.���V�&��qN���yl%5`k#��hq�33q,����5sK�M�\�{M7b*�2�e��;YHΑ�����i�K׻7ha����&���9)X-J%�����ΥvѰ��Z0"屁r��-����v�
�U���bEkeF�d��/�{�l�)U�j��~H�Нx8��Ӵ�v`*8t0(0�IRw3m���J�Q�R�Z�C��\�6`�SY�&PNB[��Z��=w܆�b���ˢB8#ש��]7�\��l�^�000�`��VQ�['oh����8�n	���͖q/ U��4Iq���.��5�ۢ���Ng-\;�Ղ�ua�eЮ��s�&�|��.�u�+�������"'`�o��~������E�އ����n�c//���h��m*b�X�E���
�W�Wm�FPFr�
�XN�mR��^>p̎�Y�P��j1u��e�B �**�
q�i�a/j[��v�䯳�OJ�3(	̆&F/2�r�XZ��� ����fl�@���WX�AIJ�HG��+�r����7�h��}�]��J�^�����'7�:�;��9��=]tK<H���7�δ�����+�E0]� ���h3����6�L2�ӭ�O�EhQ濟*{]�E�o��.�;���j�!>�w�ց��ٽ;KH�t�v�r�����J�t^�r:�2���a���ҹt�z%�q%��n7;9:s6��5YP��zZN��t�Ww=o��3�u���6��\�lJ�2���nQa�zc�6��Mq�J��h0�K.�T�o!���$����ܣXai��[��w̱օ�Ƕ�b��[�vs
�Ъ
{�&6�?8���A�f���ڛ��	H��v�.�su);�v�5ݧ�Yv[ǂՑM0�Ie'F�y��_�T�i\�q"�9o�N9�	n�`n+x 
�L��X�t��݃>Ќm:vq���P��s�V'[�sh�nh�U8�r�j� S��gاv����.�b�Y�*r��H��d���Ҿ����(A-,ك���K4�;�&ô �a�0d
�%X�$̙{K^������y��qn���+a�i�{
�n�S�7O8�͜�����uڞ8bj陋$Yl#Yq�ٗ�����+,���S&Қ6�c�K��fv�e����us��f���ƃ��*q�ٷ�U�<��LEA��%ξݷ�m��	޾���"���0a"	u��9�CN�U�J�+��닻�*퀤v��<��eG�e�ʺ5aқ��-���+�2j���wwt.�텃��O	D�3*�漭���8J!�Z���O-�-.kw��΁z��lT�mY�5����go�#V�
�U�y�[4�uR�ү�N�-	���]���͝tc�8��ӮϳEN4 y]E��߷~�s]���7��<z.��E�B���l:7�uS�Kn���}Ub�rO�^�0� ޭ��2����u�y�u�)\����fd���c��IΊm'��nRca�IZߝ��$�Gj�鮭+��S��Q���f�T>�S*��m2�O)Cn0��$���Z�a�G`�k��:d	&�W\q��$��T�͊�{an4��8�Y�51n�"�s^병ifW]΋$�(#�8m�​��Мk/i@�J����_pT��.�Y����V#qŗ�l���y-�{*q4�n�7�׋��X��pҹ����V�m�ؒ����LQu3tL�S��*�i4,��3F]Ek{��B�:,7�z�[� �3/�	N�.��[���×�2��yf��$�<���p �%�<x�q��q��+\h��Ս�U�h[C_Xm˭q*�:4�wS��:��E�}x	cފ��ެU�C%�mBSHJ���슺]N�(+­APc�<9S��Bh������Z��j�ktM����L��p��ݩ��Y�p�9N`�[��ª⬸w��T��[m��b;NF]c��*�55Vf�Y��3�'��VSN�7�zwi�9W]��o�V*������,�f:0�ӛٽ�6�Q�u�x�[����_��m�-����?��������o�=�����#��N'G��Nݓ�N�N��ӳ�$t��=;zq�t��4������v��:q�t�t����J�P�B���S���C�w���M�O����t#���Y��:�oS�p����;�S�����]]�Rx�V�r��
�f`�Xc˄�2�7W�E5��"�V��D�g�좷��a�"qJ�I4�*��j�;�5�ϲ�Y�j:[}ʦa�ܝ�@j�Y+��I`<�m��Nf̌�謆X�8Óe>�ޑd:������K�}����e� t�fF0��d�gSƯU� ��s��d�b��)�$M�ig����4z���ŷid�+t�oT�|8�G6��y�N�B��z�.bmvĬ�֊����̩ �D�y4=���>�1��5�pX�
�!���`5T�����J�.�c��.��QJ3���,̫�:�ɛ�Pv_:p�6v��5$�<�:��;� �y����Fh�z�6,[t�IY�v�91��GC���Hn�ʺ��Ѱ�\���.t��&�L�`�}�/�v�k[�Ô��vS,�(	��HL�&f�ع�)a�&ݔ:�iGm�e��PV��&%,Bz��Æ��Kk�\�:ͺz�i�N�٘6�'A�b%k����R��.�5N1����J樽��p��yFb�j<:����9jQ�<��� ��;��f��ی�Yp]H�%t=>�t�̊k�'�t��{�@ �&:lR�F�L�M�IHeD�H�T��b��?�)�ʶ�Z�8Z���w�5e
�T���7��N����}zϓ̾�*��Ws�oW-[��E(|�)y�L���Q*t���Ƿ�=g�U��)E�jR��\�^����j��qI[�N��>�����YZ=[���e^�ʊ�ܒ�"�i�3��YjUy�ӎ:x�����ovQ��9��U��T���){�"�.\(�9+J�R���ĕ�*�
SJ��9K%V���իQUZJ.�r�\�Z����T������[V�q��Sz�����}�)j�-[�qYW�̝��J��R����7)R�V��:�h���ԩJR���{�Uj�����9J��̦�j�s�Nu^��}T�;xN#�8�t��w�]O7�_���r�)SG_jٕ���T�YY9��1�=�=(J��?o��e���c��Ǻ��,T�]$���P�uJ�M�E�uq����9�OwT�У��!Wt
�U���W	4(�n�����(�{������2c�^4���71GNi����h�,ی�o�9=��-���x�������{;#c�Խ^K���{*{f��}�ŽP��Q�r x�����*����ץ{�N�&7�����i�W`�7��_Ez:|��z7��W�M��U҆�hz?Q�Vי�L�1��`G�->�{Q���tӖ6�v:�=�+�h�o/ju9�7צ��汮�\������q��۔8����gs1��K7L	��j�iڞs��6a��A��U�yZ� �'���Ǭ���͠5���N�l����<��V�6�}�g�NzqrRk^�?{���y�.�d򼺤�fmLU��
,���;�k��j��.8k1x��=�Oޏ��#����y��;X��d������"h^�`r�����iڽ���{�m�Z��)�"� `�nĻS[�/�n�T"��:1�Bg-ۃ4D�|Jy��B��Ҽ�cX�:�#W���l��Mj�s���IՑ�͜�,\�^uj}m,��)^J��� Q��ZC����r<[3=�{l���r�zue>�y<���^��%���l�-eG�oR�v�2�m~)�
C�L�.�+�WW{��a(oZ�q�S�`�z�����5���[U�a�c�_`z)	B������ws�z<ƭZ���t�z�U�g(���`p�}Y^������嬱�[,��z�ON���ژ�>Oq�~�J���|�������/�w�=�t����v�Rm�\��d�������;��W�)>���+��M���U����	�\f�o/Ԧ����ݪ�Ѷ?Fw�~�s��ۋ�*�^E��ݳkkyI��z+��6%��ї�_^IU�x���<�H#�¶�׽=��l..(�������2	���;����{�dH�m�fٖ��-��=^a֊�8c��pq�����bkA4t߰��7�8�t������;O���Y}X��:c0�����糕u��#�~K2?V�~ڑTJ�i�n�Ɖ#�+T�bP�S{��ڝ6�be�fV��\�x���uHN�����S��@_ݕ�.=�r�ESsg\���w\ܷJJ�b8��Y�U�w9�:�R>��N�������'rsޛ�{��n{�0�.�nK�uB�Y��1�������h�n�s�/�����}��]7�c�QfШ��ޱ����3F���^:S��y������U]3��K�gv��-�b;Zz�Tv=�[�`}y|~}v�*\x<����<ÓM���Wv�`Zݤ���j1�C�q�%+��|�Y�����ܯ~�V���>�;CC���{�X@�{Ns-�.H0v����z>^��{�Ý9�&�>j��
��b�P����
�~�d�^!Z~S�'����ܟx5׵�&�A��jV��������QfJܣ]w�����0�	η��s6���oQ�6����tfGv�!z�T/�R�TT�Gu�d����}����fũ�Oq�}��k�: �!׵���Btt��U���_�{��Ҷ�'+��oE�d*��6�B��:��io,�l�,���*���/Fit������̨�<[��di��ѫf�I�Ea��n;Ս��Վ|�ߒYy/ a�g�GR�T�0u(�GY��rV;t��*���Uٴ�m�Չ˯��xszw��Q���JA�d[~�1��~.x�����m���+���P�J]��]r{/��&w���W��i��y��˛�;��4�s�="�����7��j�I�9'h;zj��z��<�8�}5��3��|�_���B�|!�4����~�����N���#ղm���Y�<���^}+��B�z=c'��'�dƱD��oy8/�}�[��Í7���}�Jo����S��dT���N���{�ߢ�sw~�q497��^Z<~��3�p���w�;��^�ҺM�G[aļѣ��#�`�Kf�5��;�= �0Se�r!n�u?T���^0V�=�=�zֺ��7��ו�W��5AR�s�>�֛7xx<W=��Ȉ�b��U9�Od�y��g9�ŋ`��q7�W��K�����8gSr��Z���1��:e�x䭧�Z������wVZ�&ܲ�pHw���H��w�B�(U
��J���Wzery��ẗ́f�
Ҍ}fΗZ2��҆�f�[ce-�:0��r���Ԗ����X
�z����pr�Uq��j�PV>��F�P�P��������� �b��7��Y5�C!���������q[��u3��Yc���;9�3���N��H\�.��7v�r���/��]��l�Љ��]/\�ޝ�8m���A����D�j�����}�~�F�O/�^p��:Uq.�� �f�T�[��z;���k�/-x�YW�(t��'��ڨ���άj�"�#�y�ݚ	!���^|/=5�:DhȲ�����Ӏ���y�s�KNq�8_Og/���;�#��\�~[�Y�}�}�z�0�"Q�-P�|�q��}��<a��v�����x�myrx����m�܇��̮��^b�ƝT����a�,]S�o�_�(}�p�����-�O{��^N�U�<��6wM�����ޞ��޳�8}Jm����F�`��_�e:����t'4�����3y�&�|�mW0��D�d?����o��;�w���r��,'-��3��3�Ķ5WGYop�8ρ�O]]H�:�g�
����4y��ݠ�R44ydbՕ�r�=9B�_vU��hvˮ�h"��Rn7�ʶ;�ˌ�A֖�b�FIu��ްQ�)Ԯ�2��KI�n{��w{�?q~����F���s�+-�W��e^'Ť�9GeB�������}&'���ON�4k�W[ߤ�~�����@xzb�K�k��!�솆0ݛ"c#�g���&}�C�y�.�dպ*ڛ^��T���g':�OJ�G(��v�;��$g5���<�z_}��3�����.��+Θ�W�=M�~n��j|�|9g�^�)�5����j����uJ�-�2��^��g�ˬ�o��J�͡�O�0R�C��x��t��v� �`ַ�c�3�Y���{�Uq9����Q���޵B��ǝ�ܛ����^����k��X���43\V���]K��Ͽ{}p`�S�ZY�����>��zQ�>���gFk{t񇅞N^/��������c4����&�\|Nr��J�z�M�XU��_�a{f�u�w�K�^�=�O�;9@�W�W�]⢾�t�]FJ�5��X<�8��7r���'�;�ۥ�e>���7Z&����\>�<Aj��LKf�p�2��������Q���q����y!!��d!����n^�Щ�]؎�mumN����\�:E�Zu��;.>3�}���7"C��>�z!�h/WP�˞�8�hs�j��=���,�-c���=��Ue�6���99\o*�Î��Ue\޷�v���g!�������4���Pn���ߎ���u��M�9�"�H՜�
�����>rz���j���z�������O.�{|�|���܍9�TG��^
�_�z�T��Ix˞��
_n�;�j�Qx�b7n�� 
�m�N��^�ZNf����4Ϋc�����|��l��v;pF�%�ZrsL�q�%��>t.y)�0���y	����W� �>����3�`|{w� �=|	�9�Y��rEѵ�D	�<w;?�4�O�Y�1}�~s�1zoı��q5����M��k{�什�܇��zj�5��?���*����s����kR�ww��!b�W���>�/#=;��g76�S��1f�r�*&�t8K;i�dz"5��!�����x��j�����h��,m	��礞��q&�j~�q���lY|@�*6�'X���l!*�K�r9I�ژ�i��\��c���r��tq	���V{^�}ngRԹ˕ȵe�m�E�lA���Z�K�_|;OsqZ����+Zk��tΩu�9>�;l���a��^����\�y~�jy8g��S��M������V'҃ڃ)�r�ʢ�dW��b�{;6�^���r�Vp/��\��Q����u�/���H�ܿWu�����Dd�ї	��ͦm2�j��b�:5~�N��'p��i�}G}t㵲�C�z���%#��q��E�?h
���Q^�s�������~��_�{�ۧT]6$�W�׸�=��r��I���c7�o���F�J���=�Ԋ���b���ﭴ��rN�̬� ^U{<��l�,d5��$��h�ղY�Ɩy�':�#v����;�U��8%2���nh�7�+�.ת�:�kp��j�_	�k�g�t��/�$�p�?W鸶,s��G������T_j����.��V��p�<��{��N�Q{�*�y^�<�mY��;[�z�w��7�o+i*� ��t��D��%c��cE�;<Y��b�E���(P00��뫚'�Co�WbL\��v�6�Y��pL��i��������4*C���i	U��.r�憈
�}�[V�S�qGO���� }=�y��Sӏ�'����3��y��{S��o������k^�w|�zo�R?t<��t�����/���c\��b����z�\�S}��ߏS��[��?o���yY�>NL�@���6�����W�*�T9�DO�~Q��o������K�.Y6��ӐjZ^�դ8�ť�ǃ�����#NϬ6����{n�^�Q���e��͔R�]��.���y�C�U,�j���ɞ]���nn�{��.�|�M�o�Ly٧:�������j�Z�!W�t�==f��x=�6��o ��e��ߩ��%q�/k�5��z���^?U�/�+�Q+J�����ħ���Kٯ�{{��z��&ߜ���U�����1�N��Ʀs��_d���X�5�Ǭ	3�|g(np1>�y�=����h��U��5�����J��
��G�W0�*�{/�z�~��u׼���uN��P�����C8vg]������`���Z;:c@�2��X�2�/��	�{�L'��"v^��{�W�\�Z���r=�w�yTW�Q�b�CS�nfL4��U�l�1��zD'ь�%�g����;��v4��`�fݘ����۫ݍ��WUm�q�������:�V��&� ��vKoi�ZY㯴����	4I�6n$�>>�r�����H{�*�T�u������n��yjWsW����2r~�}�k�'��{!ͱ���mL~�k7�<"�{��d����]Vyͨ�kW�{ޛ�����U�3�5+.�Y$[��꙯!� Q���k�f�^�`ߧ���q�LuH��'��I�B�[>��^��򭰲�~U�9��O:�ޛ�{�<��<�y�$粥�f)�o��&/-��_�}uN���Yx��1�<sv��͠��Цr�O,�wJ��}^�A�.���}&}Ar�z�}q�/�}ts�*y�_�p������{��G}�2��9=����kf�9���|���c��o`��R5P+�c8�c�\з�W�f�6�m[�����d0���*FW �`��R�\��'Nޔ��V��T��^�ݫ�`N��b��ۼ��fl�����#A-�a
Oj�;�~9ڣ�6�`T�c���f��j���(f�P�ԥqҬ3z�d�Ի7Vӂou�X�BN�k�:j�5*bȝ�W�JTz����Q=J��
Lλ�I�k�xb'#SU����T����Wɑ�(���}���۰o��ʈ�\�X�WR���v�͙�]�cwz42�����͂�3�͐�ը���K�A0�8�P�W��)*"oh���o���|�f�	�+���N`諝JBԗ]�]��6F��v5�t��ݚjBK��1ԭ�����7ݕ���G�/�;�;M'd�uz��Â��J�����)��������3�:�̏�®.����/`��a�8���;�*��@ܕ��+� �w��*н.�^���GE�ޛ�&����2�9�U���/牪�/n�ߎ?s#x@���0�u������	�NÇtc�V-���Hؕ^gV�ܮ�m���N�}au�Z���f��Y�33�,��
}ўC��%�f��PB�������nP+YS��\zM�7ƌ�����&�RfоN���8q���܎��N�\��#���R�̽4����]p�S^�Lf�n����A�����*^���R�L)��7�:����֠������ku�/]�Spg��U���
(pt���m�����י�L6�����LU��]���9yR�ܧP�ܦ9-mm:g��i�M8�*uF7f���]u��V!��:̓VYI��)���NzZ�h4�W	��i�v�O���+櫧#�mp�/;�� I�=z6i�*Z��:Tk%�fʹ���ܖ�ͼ��ӻ/D���d�l�2���4���f� �`[���$��f���ض���7�$Z�<��m��W ,"�,�IV,�r��]���Z3g�bnCd��H9/0ܺ4"6��DuW2��CoMѮ�I��e�-]�!k�aQ�u�}kPX��O ē��+M\/��0�c��b*IC�J��̭�m��o����`�j�Z�N�)	���Z6��W6�\�,;u�j�6W�Η���/�����ҁ�o�i)��pv��]c�-��I��#'��K�e\;��&r�)��^Gx,�)�C��"-(�,8��v�7u�[ٰj�XyB�f!�S�J��3O&��(�����8��m;vp2�8��}�՛��5�9���ċ'R�u�9b�I�1f�^�Z���Y0�b�s�ْ�ic�%{�f>s{���c�0*u�c��Ǚn(��g�����-k�o�\M��0��1��"����̺je��q�T����'Q#���ʰ���9w.�7à������ӈ
 v[wE�}vXs!���:n"��͙�͑�&qS��^�)�VԪ��4�$��+S���]s�R�Z�z~8������������V�H�Gە�;�e��r��H���S�ʿ:{z{x���|���h�%RRMZRUV���W�r_9�)VIn��;v�����ӫ߮9-JTZ�8�jU[�ܤ��T���*��9��/|�׎�=>=��x��H�J֯VⲕJW��պ�Ns���=\����$����W��j��Ô�RKUr9Z���[NZ-*�V����Z�Mjy7\�5V���̔���}�R)Z�%+�橪IUZ�J��*���V��Ui^-�\��q�뜔խI*ժ��r�j�i����^��I^s�Z��%�yq*V�I�QZ��*ժ�뛕|�U&�ս}��=�U���q���[@ů���g	�	S�]���5��a[�  �Oh��ÅB���mB���CtޟQW�U�s��x��'b�t��C�125��9�.g{�eJ��<'���S����7�w��04l̐��o�����/��Z���I2Zc{�}�س��0�v���ǁl�KH�?)����T?�N��La3�b+V�~`(���̓��I� ��ܣ���=����y��ij�*���A�v�]�m9�7ЪV���ixz�Z��ǡ�N��(�;Ta���~�w]���u�g���F��Aܴ�fy�e�deegA�!׽��h;w��*�v#u_����J���U�f>*E�d��08����0��,c4��k��p�;6� Ũ,�M���^e�ڧa��2��@cr2�:����`���qo��j���z����LP�!H׎��yN��tRr�����!�ٰ쪚<�5�,�0�廼Y���/T>;�Rz]���CY}ao�O8�+�TZ~9�T/hZ�ojrr�R�}���[����g ��D$���h\s4_O3���J���
\��9</(z�n��6en�=ΜYf��"jdlmH�^���#(g���X�������o��F�.r|��b/ע�L��'��	zw\�z���6�n�1,,�g)ö4uY�ي�S��$4�p����'�0�G]�2Ｔ��!��c�;���yd'1N`�c˶�^M�X3 J�wˏ����u�N͡�㯨V�5ё��E����Ph��|�[;��Y�C0z���p�cz�aR�ltLwx�Ø	�A�x�xhO�EH�y��A�n|Z0��-��L�Gb���-��2���c�<��%��V�+J �墏��Ai���G¯+��Zݻ����ւ��R�&kg�ʿ���>�'�j8��F�i`
���ى�An�G��^�5��/K��3bˁB8��m&�qڌ�i��ГbUV�1b��v��i{g�wbͲ�LЙ��C�Ij�Ĵ���&��g��[�1�3A���Ի��iY��W�o}��nz��IY�����T4� ���:b�d�c��c�����F0��� �����Y������:?fc�1(���GD�QU��ۤQ�������FdM��'z Ƞ{D�Y]�Ư�1 ��h;@\L�[�>MF3H*�����Sp~���ߓE�f���玫��� z�V%�%��ic뉁i)�z�v�aq�}v;T�+��Ҭ��02]R�gv�T	�*�\Ib*żի�U�4�k_dUo �M��{ҵ�e�m�m
��ߞ];y�D�a�F�smt�}�|�eB�e�/�Jsz�������g�`ka'��{U��u	���˹�R��Ӯ��Q�]]B�VS��o�v¦ԕ�M��V�867ep�p=6���i4+���\����Q�(����aG8l�p.Rڥ�r��z���F���d�nw�:ɏ��+�4����(�{<��%���2祑I��;��{iVk����$ʫ�ɈG��FD0B��SE��j��j�3���fR.q�N�W_6�I�ҟ.]ۭo���I��{�ղգ3��N�^P6 ��׿;�8��� �|{�!�VH!�_@f��'����2%3��-D�4�F�t#�;�
x^�<�ڟi�T6�ͳd)Ś��x'{0q�)���*/�h���(�⮺�B(�t4�L(���>(�L�{�y��R�ç�|�f��67``�lPnCF�{B�E��ByO"��EU�FU�U�1~.�z�y��l<D�D���__?{n�g����}{`-zb1����������2��5oL+#��x��ü��_]w=�']7����ܝy�t*f�@���7<�ڜ�E2��-�����R^�G5���!+η����
j��C^�'a� [�薶@a�h.Y����?5�xX��9���2c��C�7�\[fw0�p<[������i�~�?����')M��@o�L?y�t�猦G�E:��c�\3g�F
��1t��vK�8i��i������b���Զa}˶�:t!49��������|xR�&�?�:��̯�ubw�G�cQ�^'����aL��-��Mv4l�L�:^�W�Ev��/�$�ɐ�x+Ss�{.T�tߵ�UK����{T��#�F��|d��g6���~.1�t�P��Ss�V�k;`�p��Z�[$�z���g-G{���u�p�Č��0�H�S���A�KH�!)�<���>Dh�%^�����s�Z�'������w8~�c�_�H��gB���¿�7�r�7#�ˤ�6o�it��y.��v��ի�*�n���ûo3���L��Ѕ8-w,uOU67q�&��&5⮅!h�:S�?��36P��W�U8�E��ŋ?|�\����X�����o(d�1���.��keo1�u���z_����?Lt�Oc$(0�uDf@;��9.֠�x�A<������b_/��[��3��σ��e6�TĹ��m��m���!��y�4ܻe	�˞�7:s���S�Q[�󣖷^��vUw>�L�t��ڒ��M6pY'_�I���<j��V7��<:�|o&}�}ñ�U;Ŕ؄�C �`>�R�G.�Ϭ���T7��7J�a�"74	�3[�(:{km�n�K����S���Y�&�m~��,��S��	�����A.�y']���A��t�<�/f�pvv~F(k6�2�C��R���J�W�H&��őt5�MAX��]�RY1�  !�6v5O�[+�}���G(a ��V�jhz�K3��prK�o-�	,�ި:�+�mMÓgD���ö�..7�kZ�R tx�t�I���R��} �5���h�u(��ޟ4�V���cg�)�X�}��^�K�I�FU���OP���n�%0ZN�K�рͫƢG����b��L�?�u�zX�~�'��Ӆ��{/�6-I|I�K>XS�i�3�h��mC,�Df*�t_eۗ�Sڵ��.�d[�IEۧw�5*�PT���:��=��<�;#����O��-\���3l ��n��l�s��^l-����@����ʇ���U�	���A�_+�Ҳ����+�P"��uH.c��dW+�L����<!M)�1���CJ8c�e���r�K����� ��p�|]�!�(�#��,'#M�k�(/�� ��4������e���~������m��ѕJ�gv,��x��SN����߫}-P_Vlg�y�_�Ϟ�`,ч�=��߱�aR����i�!k� ������W��6c��+*�z�n|�$�q�ߌG0��_WS�X�j��@�9[�
�V���ܐV�����d�,�e}+&Z��ƣ�S������&�gUS��s|�{���L�ao�t6��0�n���:�H4���<;GJ�ǹF�4�GM����� ���ױ��xw=�'Y�U���ܡU�e�Ny��G&��0�Ȱr�UwJI� �b��N��f�sF#n���n�Σ\�����^�WϾ��w��~ɥ!-�U`0����Oh�ۇv���>kށ�q�^o�u�)�d	kA)�{*1�_Fl=:zb��"g��ҳ3��Ȥ%����L���.ۏ��>0�>�<��~*-?�B���˭����b�$���姐�F�/�
������ �]�j<�%��]�q�۹)-��T'yO�{q�X��k٫�tY��S�ݔɺ���/�������S>��Ք>����Fԇ���&"��n��~F��?��()�l�rY`ߦ;�}a��`-�M	��缚����U�)�֟���V�SA{(�e�b}X�.�C�ݶb �̟�P����.��	CV5C���n/����Q��l��B{[z�#5�Ga��W ��'@���h��L��z��x�t���%��1�<����n��Χ�Գ�FP�U�C�Xh.鸳�rw�S����*����wf�ڝْ������a��`�1�#�?K�,0��r {N��o/q�-���S�1B\CtsBW�����k�E������{ �;��o�����3Jv^����H����r��bV�hS��s2�DK5�� �w��8�jF��c����r����&L���+�Uѫ�]J�B�e`��_g�-�#�>�{�A�9�RY� e麒c��cf�s�œ����Bj��
43�]j�r��1@z�Q9����W��|�si0�c����}w������*�o��6��w�Ӳ큉�-�"��@�e-{�W�����u�õV}�`��EK$��zCnR�%��v۸�gs�4���LozQP���]8�o����� ��ٽ_!<�M����1N1���d��}�!����`C^�p�<��᧪����1�ʻEnv����R�Fm��o>��a'eR��G��]U�%d���5�)��C�ҵ�FP�-t�Lm��2��u�Bς���a��y2j� SϲcX��%��wBe�kb�׋h^���}ih��KmU@��7_��<B�q�wmC�v<��i�ۄ��'�X�e���C�����K��UX�,7S���LJ�MvЫt,�Vy����5�ޘK��R���2����`3]j��F!Y.�#��a\0�ݣn�����x�Z�����#v6��d�75���cL:e�^�!���g1�O��3_2��笵��L�΢á�qu�):�s�6��^ʡO�>#�|�7�8@O\��dO����՛�Zi�8��u�)ϫ(���B�J��.Q4Y��zg�������x���ψ������9]�4����j�a+e��qe�ru`T�x3g�s���ej���P9�"��V޷|)U��6�/S�c��ݤ"K��4wa7*$*p�m+*�(-\��!>yr��ts1i7)��V�g�R�*�T]��\�V�?U����a�� ��o0�K	c9�����������������k�M��6zf9:��tz����
T8�Y��,��`�,Esri�g���ſZ�'ş�U�C<�R��P<(D�s��jsu�o�����T2ʞ|�6څ����긇APZ�"��g���dȜ
�|�]2Uw�CW����	���\�;sA6^��\��[��m�~ʵ\�b�kz�\ϯBMIj(Mz\ߺ�t��>�J=uY��襾����U���Y}��q�a�|��ҩ5?@����,��P1�|�R`(�KC��M�~���˧���=<0�*A�oL4�'Z� ^d�f�'~~16P%�`���4�SM	�]E��b5�����u���ۤ~a|-`�����Q����^�f�{���Ͼ^�����Ϻb4[��:}�E:�9����T'`�aۍɦv�nw��so9��-�~Ԫ�Z��D��Peܼ<(!6��}�o`6$��?O��c���E��9�pw}�P�={X�:��8�o-úUcm5Yw�[x�!V��-O��^ｯ/���<�k$(0p`f�"á��ʽB|�-���S�|�����6(|J;)��o ʹ��(��[�P�U?�V��H�7�ٮ���e�\�F�}:��N������}w�a�mm˨�P}@���l�A�� eI�r�3ۙ`J�8y��\e����C�9o9�?��ze^ӈ�UW��4�r��lr�~�����:���]~?_�U��q)�2YnTȹ�$gՍ�1�la>*,��y���ϭ��]�{y��$!�8�ksupآ!��r=gd<��.{�.��%��SM��N>��m��\M��]�g9���zz�x��[��g΄�˷5I��d�d�y�4�� �*)�s6_[p9�AR������;i�ިlxx��V� xm��z9�~S�\7��NP�%W'��	~Q|ێ"�t�V
32�v��&��x�2]Qm�E۝��y��0��6"o]L���TZ���*���sz"T<b˜Kso��d��P�8�n������u����^T�*����;�A��%�5��ֽN���v����f�y��Y�T���*�y���V�Ů]���o�3C��]��7-=r]�O�8��{�^�#���4���x.1�}L��1>����-C�����m����U]�u�\q��ys>���
0�3c���c[�����C�P�\$� ~%՛������͹�fyI|�>0x��@��j������3Y� 3۝�I�{3u���@���w�B��V�AO\�/YP^aƍ�E�opk
���{L�ZG_5��2+�$����;a��;���z�K媍+���0C���R����wUJ�o�e2�VX��ɮ�A�۾�Ϊ�fLа�y���9����{�@Kl����)�Mϯ7�N�z?�UW�%�-�Lqf��V������Kj�ȥ<�� �Tc���?6��l����9N,˙+���f���~�0�jm
&�����?:�йK��ަ�����u\��4�*i�0��i���T�H�c�#�l!6�|��;}�z<�D�/uny���������pv����!%~	���~�0Ҽ�u��kԭ<��2.�����P8΅���:�9�dҮ%�+�[T�t
qZת2E�oq��3i�g &��Λ�߳YSՠr�l�w�A\<z�I�&Q�)�u��֔Qy�a�v�N��}��m
бw	�oP4ӋZ�4y������;wd�v�s�.qC�M"�aQi���B���P#|_���Wy�>7]~�{���1��h��{ �@�4YڇaTZø\�yi]滨��Y'g�S�ҼUOZ�5^����]{%+o���+�@��ni��M>��v!��9잳I�����_�ow��څ�m�����J��0�],*�cFu��+1Br��=z�S����p�*��"��~�F^�Bh/^=�����n��*��Hݢ�XA`7���)���pp,b�I�]��&%�f�4լ�(�;��*oU���r�U���3b�;7�9F�]NDX�:�B�w�Y*�ƪ� ����GO]{��>��C�=:.S;㷡�d�[�jJ��t�+]�4��wFn]e]n�ΥM��ʎIX����'{[������zp�!�9��WB�Z�w��%��*��vY��N�8f�h���V�V��؝ZƉs!c�?w��sE��^N�uא=R@TRM1�.�����z�m=�uY�V]s̷�i���}�%����7��ѡn��Ϋ����k�[Ǥj�O���}eĔ�bRbt8�1�$��ڷq�:23��	Î���;7���fH�M��eb��jr�r) �ιiQv��e���������M���:B๢�_:�}̵[2��ʹG��ݽ\B��,�v$�c����莥�J;kIJm#w�݂
���A�fB�2��><m�SW�,��Ԝ|y�=h��� W�p*����k�X�ȱz�2��J8���N�Äa���t=;����ݫ��E;5�2�R���3Zf�\�Z2gR��+M��E��J�l����������<f��n�d%���=�G$�QS5d��W��*ɳ��d�Rx�/m����F�ɪ���)p�r_����4M�}g�;��4�:A�$+]>���t��Wc3n$�p�3C�u7�P��^98��O;v��zG;zq:zvv�I�";v�ӧn�^|\.�%I.e�]p��N}��]��f��ס6�L̈́g��Y�5��Nt}��{)fm��&�Wh����|Ǝ��q��w��a�5Co֌VC|��%[ouY�ۆ: �8]��`�=�Nr��C	�z�p�U\-Vzά��q䚻�+}� 5�\�q�������T�l���y�̗���!U���υ�3��]֊���W�ӕ��	η��X�#5�ͨyoCD]���ެl�d�'�xؤ15ݛ �F{��F�?�sn��U.���9����Yx�wx�Ų�ψ�\6'j}EDQzY��u��(:*����
W`k"�/�mլI�7�J���f.���L�N$H���#��^ʰ�5����ƅ�%�)Z�p#2�F�c���T���E��4r��i� 3Z�jGFp�7pcۨw��]Y�ܫn�.2+1%I[ז�D+��7�� ��y�>Mk���J�j��W�!�	�:F�uጾz�+�u>���$_E�X��V�z�Bxp�D)�2N�^���;f��#��WG�t�kl�n8ڋ2���|i\���%<�X;zj�Χ\�ʜdi�t��//����0�s@�b[*�r�-�pΰ�yԶA�(��vMD˕�x.M�bB	tb�O
��zc�y�խ/)�v��3xgG�Jp�| t3e�7[}���8Ӗ�I�6�@*�<_P�!��1F��c����^Ύ$l�����v_h$^�w�{�����)�w�j�չKEMRS��Z��k��UR�iUjIi�ӎ�_�_^��&�J���Z��L�J���J��ۑR�j*���ӷ���ׯ{]�9��RIe*�KV���R�d��W8��r/W��㎟�<z�ҹ��\)�,��lⵕ{�nB��s��<�����OOo�>on�2��bU�)ݛ���s��ܵ�9	JZҲ��ұZ�S9����5*���Ք��)��U�wa՟g��[�qj���ÑJ�Z��nURܳ���̕((�rj�nm���劖z��U��W-T�
ԓ�NJ�*��QQ�9�Y*R����ݷ"�w+�D��8��ϫn[SV�wg-�U�N\��8����9n}�sZwÕ���:~?�I۷T�R�J��o�N��`��k���jKa�V4ġ�3�l_v�,ެr&C-�Z�\��Z]/(lN����3{��Ӿ|�ϟ>y{�������v��c~�f�%�%���C:q���篾�s�Y�$G�������-%��0��4'������������ �hb�>�^]lCB�D�K�9�[#�;0��t	pp�4���#O/���8�(��Y�"�Ҫ�������;��\t�u.�4c�@l�T���:��=dB�WI���V9�97�;<^2��Sgp�/����̭U�?K��8�
z]#��@�o���'�D%���G��00y�l�ˡ��^��͍��%�W<_;�2큤%r���B~hw���N��F˼��D�k��nF|�G�ѹ����G�H�N�&����8��3c�-�>*���r��U���:��"�d�DUDN�s��I�$nj�t�s�j���^lԵ{p�X1��Q������P��*MC�*ql�=��8`���e{��j������ϘQt�j��}��)z:l�,��F��4�>�|��C��VNmh��1�o?��ˬ�vYC/*���?;�'��
�P�\�[���\�^S�*���-�w���o�"H5�9�)�a�;��h��6ӝ�^��(���V+���J�t��+�e�~����]J�ky�#�y^��Q�0��e�v�	ڬ#���ژ�D��]�p�S-���7��� n�Q	d�N��x�5e=6�:�޹[G\C�P`�;��qc}�'�*Մ�Vd�w�@����u|�2f� [Z�qN��uy���M�m�Y�[y60k�=���m��>$�[b�����r��z��qM!�*_��O�2���̊4*Bv�n�~����ɇF`�I�Ys�Q�T�l����P�e�y�1��r��A���5j8�5��%����f�EH	��r�-֡[�������i��#"]��{���/�"�1�o�=��N��6��_�2Y'�O���>�����.��eΚ����A��5`*�t���������G�8ػU(q��P]c�=�7or&��ݗә��lN�x��� 0%��Nސ��?0f��7��cS���󮙒ޛ�J��TRT���Y�ŌN�ʭ5�dz�z�&{32�ܞ��]�qg�O�Cϛa0�����'US�L�z���9MW;�wv^2�M��1���}3�?G�<�4=+��/�#J����KV/ǔQY4E�nZ�q5<0CC���o����~�^,��3JUI��4:��,��G�0��Lчu�mw���n�!N�k��
k�I��Nd[Nt�Ϧ ��p,�`��i�>�]�����9yJ�.�v�gU��p���FQ�i;�O!��M=7h�k&�gV��l]+bI.`V��� �b`�A�*t�M� q�ܭ�:��ګ�iP{�8��o�Y|C�J��w2��0g;6a��;3\ķ��cO2��[\m�c�}�����Ο?m�ߤ6HƓcF����{���-�j6�5�}~�"[e�xO��(5r#۴n̶5n�4���E�Iv�ql���ѓ���p1O��u�)�ֈ�����ĥ��g�k�u>��;�e���M���8Έ�m�A�4��r�L7�hҷy։���*;�b�'�� ��3]r�o:�u:Ƙ0n˵v��e���Z��ź�q,s�S{��^�u��Iv"j�������w_q��CHF�r1k�T�������XgDWa*�<��ڵu�))���~|�S5�>��~�+e�-I�n���w�Ta�X�4���G��DIt����l�E^0��P�6�_shT�WF�)�]CcZ�;�!��Z����h��=�&�q`�E>yDQp5�ڣ�wm��9S
;s|�چMD��S�6}�d\�+gd��9�_���E�?�&(E��S�ڪG�������x1ku���{i�G�?U���Mz~��
q/~Ns �&[�ݛE������k�d�EuwN���|�a����)�ҵ�]��`�m�ʎWԻŅ���8_�����\��Ca�v�ӑ�Ɓ�sP̃>|�_�_��@���Wm�,"�{qo��%l�9�b�a���3Wn))\m��{Ƹ<�4��rM�R���4��Ρ欫/���o�Z�SVHL��{�su w*Gt.�M���y���<�ǿW_:��m�#Y�#c�a&ٶsϾy�:�~~�~?N~���u��M�]+,tr��t��뇠T�5x��vT��s���n0h��V68�k7^)����<X�!x;����\)V���r�V�c5�׫*���o���-�Z�l�N;j抵��S�7��݆�Lԛ ���s�(I�/^�lt�Ǩt�����aɜ.�X� ���2
�ymP�]���Pc���;5�0�}'$�	*(p�y��}��q�m�x��K�bk%D�N��w]�*�Wݎ������>_�N �8���w�3�ט�pW�#�_�u�H�oOun�iC��m�0�5����~�G�W��a�j�=�P��{o���w32���=�b{��U���+�_t2x����sM��*bz����e���ǿO��(s�N�Ȇu�mJ`a{����
��:d��,�l��εV)�xk`ܢ"��c��*d4ˁU�V8���V�@�"'����k����;���|]���	kԦ��=�8�*秶g4����K�{��/҇εE;�P��m��#Y�ͪ8��&�����G7�Ӭ�NNTJ)�S�f�Z���xNvP;���-�7?]��E��r:�Ka�g��u�dج/Y��y�ز�5z��B�VU*Th�*+h�/��W2�	���h�b�t����WKkx˛���~S�ޝ-�ΞZX����3ݵ\�l*�]�u�ߞ���������\}������o�f8�f��m#6�����?;�~�>�+j��k����n5o�c�Tь I����U�؏]��.�j��ކ�h���Z��Lt��NB6Y˅숬u�M�KW�_�]i=�;ヂ^=K���o��*���4Uw�"�ާd�jZ��%�O�[�5��9`ߦ;�3�i�A�~獼�4�h�λ�F
�Z��Ý�]fB��~nSA{�M�%���o�'%j�H֖��L�6�W�=~���j�/FFkԸ΋�=s���B���q����[���;iIM;�Q��t�j�r�c�HM/�Dc��a3�L�v�zO=<hu�H��FE4�{!HC��KG>���r`��6~����Zx
0��yݨ>-�9����	bkds��OuP'�v�&��n�S��t��zY5+ґ��TEz*ZUQ�QM�1Y�.d�t��A�і���,��^�=����IN�#@�ގ3��_��P��OH�*K墾�|�g+��>D]��`�܊e-v�؄�e�?�c�8�Ts68x^������:<���R�
{7ʿOO�6��D��V���<�!:��e��oJ5�.��e�,������m�k�t!�G�]0���V\|y��H"���f��t}w��6��j�s;�GK&v�l��y��sp�� 撲�%-�L���O�[�����itw}G��|��_���[�f����`m�ḽ�m�￟��u���?��qmB��x����~ �A���-���p��*���-	�����XKKT'�(D{�
Ǩ]�#��op��?�A�zZ�E�mxV����{A��$�;�<��~ވ��͈_������Y����G��c_t+�x�����V�c��z_�M#�KVн�ku��յ&��Sű�	��vH8�r���з՗���u��Zc0�k��2s2��x��&�ؼzqi�,n˨�����FFH��@bk��
anfջ�!�F��0����s���a�����J��կ���A8�*؅«g��Z����ͅץ�k/CS���;&�jS���RdtTO6�*Vw�X��;�D]��CJ�������]�ke�Ip�3�����z��'l�0��)��	,�lO0�E�-ٿ;r����K�,�+.����::�9��u�'�U(q��P���\D���k�/l��-͕��-	�|#�ۖF�$�d�ñXA.���=��P{#KO ����:i�u
up��4�mS<��R��{�;N�cڷ��9�Ǹx��[�x�w������T)[m�o�Z�I˷nfb���.A+��X�~:�QW��K�{J�kf���:�M>��%;_]��Ff�ˈM����Ǽ��?)�z�_|���~.��9��?u��2M����pͷ�^{�_������lr�����E��z�UM����c|]��iG���W��{�s�b++p��&%C[JN+M~s��(������2���R��@?��@ç�:/8gw�
��IO���K�.�B�����;fq�B^(.s�OS=.�����Q���&�Ns΁]����}�3o��н(5䈑9<\T�JO��Ml͹{<]��;��$����7�V�8��p=��f�5ި�ό�����Pۡ��4s�*L߭X����v@����������9s%H��E���\=�P&�<�z����v�O�>�	n���u�M'u\��?I{y\o��K�B\��Ml�
Z�#W�X�c�<�D���-.Z��R��G�_����"�&HN!�h���\�ƿX�LA�Ntr�m7�����WB�bڈ{lw\���魱�����楤��qk��P�5�h�0���}�2�n��n��Fm��j�QQ�~f�yOn\�<Mu=���p�4��dU˶C�˟F9vC϶U{%��f���m��u���roҽ�S��]K Cߎ^��kӔ��v-+��"&v) �aq�U�(�����Ck��T�2 R�q���0��S��g��a� �7!�c�����_M�yH��n����pE���B�ֶ�qE��6Z8J��>�hm�-<>���瞯|�뗝;��`��m��3%��lrͶ�翟���}��ׯ�W몥����8˶�	"u��,��Ɣ�2����E�g����m�r9����zyW�g��)q��p�B�rS���[G;k�dK�%��Kȅ��)���@荫�{��-��z���L�N�8�~bƉ]�	+Ue ~�^���_�ڙE�Ĺ��i����EnT�md4����B�`n[�^v֘v��l�x�C�e_=2q!�*v�鰳pܣ���^Y4���x��g���r(י�uUkW�k�cZe�;�_�۳�ܦ��Ԛ����^�������
�r��;�/�c�oG`=�&k����ܽ��i�zV!�s�&ocj�И;,03�a�F�k��A��a�a�Yw�=C(�1y��ǯ�a�����M����JP@H93�e�����X[��qeEvl3�lCH�iۡ�J�٢��M۴��	k��U���O
�ɳ��mU o[�{�})JjQ�n�}<�0ꓻ�Q��iOx�P����<`���2�1�ږ)
wЋq�	WPYR�A	.�Y�UV<�jm5�V��xSL��XGo8mM�f�k۹��:�7�o�x���}]��o$+`��rs���0o��Td��FL�E�����mP�[_�*̂�DI��8r���EN����Z,h=�O2���5e��,K�˳I�׵.B�l'I�S�\��t�I�O>Nu�s��?e�	m��0Haɶ�G����럟�??]{��眖�?X��6�$v��h��2�⊒ͯE\�e����:�$��x:#0I���o=0��*f��-��7xD����Mu03^}sRQ -|�A��,�l��m�VV��ߞ��}:�����wk�2����s��ӻ\� ���_��wE'\�E'7妅�����B���s��v�OsZwXz��aU�vld/^RM�!���O��Z�a!�I��ec���1��n�6Eg'�uj�����/�Z�4��)�v��OD;�0�Q�u��\{#
1�	OE���ޒ�X^2��2sL�~��u�+YC`Ԉl]澶����.z�73L'+w
���L�׭k��5��i�g���.�y�����E�a�s�3�i�A�7�5Dɹ���a�R)�*z��~��E�"�om������_V�=z��u��[�Gw5�7�P*�l0a��\;��7I� ��k`��K�:/~ۋ�dU�T�iܞ�l��5�o��IWo��'���zߐ�7L����ks1��<�t��z\v��I种�'��I\6G� Į�7�c���b�t{
�s�^T�]aFު<����;&�&K��]�c�]��+L*8�&X/&��T]w`����E�7�5^A���#w��is�o�������A[�3M�ZfH�Ɂ��C�4�p��7��'"�u䖘t�o{�'w�{���}�}w_U}_ųd�i���f?^~~y�8OT�;1:ۯa���`����!�y�vlP[$:�5��23�`,�����4dS��*���ߐ+^�АS篘=���C�y��%{!86�s�U�b��V��١;C.e' ���m�ʽ>G3qg�w��]�4�%r��1О���M�+^�L�tlL����J58�{��˽��si{�=�� ;o���<O�'�ly�s1U.�|����6�O��ܛȼ�#��;U����u/X⚮�#�1��ːT�Aغ*�#�	!���X��Zp��gu��UC�]��*l����@B����FWU��J ��j�D��J�f�#\	�� �	V���f��<�C��h���9�����ᵘ���{�W��}<��>�]*c��Yt�͗9�"��U���jۆ�˴4[z4��W��g-�6VA[ǚ6�+?-��-q_|ɾ
KPfOΊ�.�ؼz�yCo����>��SHp#
�ǻ+��Srɡ��s5�X�*C��P!�+�i�+���s��Sv�§�H��'�v��?3��x{�{R����}}k��e���p2��TpýNd��.�Y�e7G2\"�sX֥f��`R�v���+e�kӏW-�s��)��ۂK��L;VW7X��A1�\d#2�9W�uH2�����(���
�N}��رG�$�P6�,C�h�����*Rͽ{%̇pviM��B�����o
������,�G�������^"�
V
s��؛V��[����.�ξʅg9�ur���!tM��p�n�����4�RN� [ϡ�h�|T��M�X
�w{�%`xvCV�F��S�w�z�D��ݝZ�
�����UM �4�V�&Xbn��W�PS'C;A��9G6��q��-l9xwqۦ��Jn�έ�5�
/{�Z��V�/��s�tw%�WJ��C�'��q8(Ĥ!IV�p�-Իd7�G;�������x�aV����%�s��̓��=t�r�CdT=B�ԵlF�txI���1�׉Y��(�L���[���!�[hvL1
<n���w��pU;�L�v$R�d�w�(��s����4�D�u���N@o�Ӻ�[�;c7�^YL�4�ζ��Ll�F2�(���������87]y�ֶ�|��ؼkh�!�*�؛1�!t��w��t��#�k�9`曭���UF�-ɍ:�&f�\�-��n�}02C������QkH�4j��ɚ/�3K2��K�*-T���d�h���÷������~�vb��E�^��2��lA��j�M❨�b%JJd��ustKV���MΡO:�X�N��z�<H$F�/��/��Ô�&��YZ��0Q�.��閚WG�A��A�Kaɹk��V������]i	�J����ǎA.jh$cV�[��+��)lmZ�Ǎߖ.��� ��L��r�;�:��%8ĕ�T�6��U|��V�:�q�^��j�/��~@9��ӗMӛO�ۗE�je/�:T&��#�[z䕆�mH�]A�r��"xghʭ"1�u@+t�(���c�۽��$�j8�j���8����S:�G�/�:ܣ�k�D*Ir��i)���U���2+�)H&wt�Y�:��i�`�p{���n��oeGdARV)��j�WV쁹ϊ��tk�Ff�)��3�����[�9o��%]9;��Y��
6sunM���N���(Ud	ŵۯ�U�*��6\�R���\��p��yw�k�eJV�ʾ\f �.�k�;&��u��\3���LpO����@Y}I���s�NTE�k�Fi�r�gM$ ��PR1Ib�L���J���ȇt$�uqw���UR:��OK9��^��+�������c��v������&�9�h�����J��7_#�V�r���^H�Wӣ�I�$���WY
����]Ԣ땫W�p�����o�➜g�N+QMZM��:v�������z㞭�*��3����VV��q��R���˾�4�Z��ox��������%R�S~&��Sz�ikEj�R^~w�;��K^��۷������X�s��+jf�[Vի	Sz��.��]�M��I㷏o�>l�2�i�n^�rVVu91J��[rr�)%j\�"�\������j��[o��J�9ME+wmʶ�l���ŵU�FI-���S�u�Q,+)�Er:⯼m��L�,wR[5jڱ�rՔ(%X>\�;�"�(��Ǒ���Q[*�Mw͛�(w9:�3+���u�;���]��:��v}�} ��l��}��zC�=�qf�*�d����\2�����mFr�s�=���΃�v���ߝ�~�m��a��d�w0�xxz�4hy����ҟ����zǔ�,�=xm0��b��T�=���)X�����p��K��G6;t4�hwb�#X�&n/��ɠO �ƌ:�b��aIt�q=��6�N���4�+]J�#��	�R�<$aJQ�	Z晘IՊ�m�*���5�v9���l�����;��i��2�RX-ih��A���Õ�����ZZYZ�zu�B����̶^w ՘�����p��Q��῏>m�]�x�C���J��t���ݡ�OFз&N�h�M�i��5���k��5����!^Nn|.�YM�yP�t�ӷ8�o>X{i�'nk)��B�gu�>��m�7������e���!*���3t��_a���0��M�+fS�����s�w��ЬK=�7>���4�{���d�Hm�Ii*�d!�Zc
�"3��d4�2�?y���$ƿ�R9�G���~��T��7 ��x�(ᑏ��U5�L���R�	���<�>�]�k�1�>�؋#��pn�p{�L�����y@H.��\Q�K,�ۭ&��gd�r.��v]�)���m�&Lת^���p�wY0]	B�^}�<�?\��Ί�^���a��s� @�Ȩ�VNI@u8���E��罏q
e�r��.vЄ�㊰�ې��>��2�9u'��^���߼ؑ�M��f${����f��� �	�OK-��7�iO�u���`t+�0�/=���]ܹw�.���b	�L+�=��?*��vN��4�vW�����ܥ��(�[�k�Ty�O*����p��{�z>�g?R���u��ٳ� ?�3���-�CE��T#�K
�L�
�d\����7_�ei���'�<�C0�R���v�B,bz�^w�b�v�p�s��hvC��+0�9�a^*��v��b��ӕ��"0��ަ�h�Co��C�*[�%��B��.����Md�}�+�y�+�)���a�S�Z��:W3���/��-=)��+~j��!���Rvԗ+>�sk&��oWN�ɬ
�;&y�L҃�^�?n��L�:Q�<�e,�3�N�݅+��O�C���F2ak6�F�6#o��kG&���6W��n�	ܷykT�ipͼ�e:�	�К��h�S{T�+|�?$=�
�X˾�w�����������y��r�֡Ů]�x��4��Gc�����,k%׃�{�!�8�K�| =}��a�f����?46���Z|w��n����L�g^�Y��u��2fo*�&�qԭ�׼�7��R��Z7���J1t��\�ve^�\%ȸ.�,��yx���j7rHm�*�(P����լǕ"�x9�^X�3.��c��xr��ډv�o' �ϣ���Y�
���zS�����/��z+��n�KOB����z�}u�]����=��#g'ؖ	6�;z'�ם�������뮞�k���P��	�r�H�yT�_,��3����05���iw��؅I��-0�߻o����*�o�֒��ҭ$^~/��©R���m�e3])Y��my}7�^fRl�؎`ؾ��wg��,s ���cSi�׌�Bz�����|��%AK�4��:s�L�l�sY
�"�z��T͵]�٦� �!v�SE	Uތ�>���C;-�w�}<�����"��Bj=�WՌz���B�2p6��ͯ@���]q/\�p���N���p������4Tm�I˭�kѳL.$�sR:�l���A�q,�,rڦ�	ek\����Gd���f�ޝ�1,�/;�X끙iݮ���Nl���&ߚ�u�%����׺�il�
�fI/wh�ثze�ձZ���_�ް�^1Ѝ�S�>�dy_F��o�J*��&��_;j�OKe�en�1e��<�g_�m���7&���F0�)�� �#��p�O��p:Me�>����E�����̜"�;�|�2;\ٹ����bZ��5�7̹�ypZFm<\v^L��sz�����3�]�]�8�:�;=�b�{�ōU���5��=`����f�l���Ee�*9� ����6���ݒ�&V�.ueJu��@�'�ݓ`���oJ���LQg	��W�E�����L�f�ؖ3��_<�%��u'M�/�kw�P���X��_��;X�����o{}:ĺ�¬��^�s�`��ƭ~\:���x���]��|�Sv2�f�4���[�'���'Am8�V�e>�z����ݵ��G0�C�yh�Eꞵ�M��Ra���	��Ϟ���B/ot���^��2� ��-_�t�����󭟛�p��O�:?=�r]�R.�j7��rȨ�Uc�(��XC��v^~�s��>�k��%�9��bC��C-�%�(nL*�w���m3�9�=[��b����1�����j��e86� ���/^��8z� P�|ws����Z�� @��|r���9"��󢒼S�[f�>;���@�<;�*��K�^��w��.�!	�L�'����ْ�z�Y�{�s6:,�ͅ];<�Sp�1؆k�0��U]�馳�#�ʗ����N.�9:��-P���t��7t�4��@*:�dKe2��Gx<xrg�؝Ex�3K ߅up��O�~�����g�k#=�����������uVKL���wӋD�̸ʰ ��§S�ɹ���X���/���y��dݴ��O���PS u�m�:��������:O�ኁ�;|���Ć�ɛY%]�1�z��G	��RU�
�Fɻ0��Hk��� ��J�ra⮇fE�j�y+�����7�>y�a�#K4�,�wl���������p��J<����i�a��\�<�C��ʿ�W�Wo�C����F�G�Ct&�<~�1���j�kj���t�'���킫u��յ/�v���Ѧ��S8qR/�K)�7���kA�h�O%�N��s[��O��	8�N+�x�j���cZ-�0)Z��]x���~�ۚ��t�N\�~��B�h��F�L�3�.}*=�z�bg2c�����4�uV��b�Q�E,<��r�\b���L��i0�jS��.#�y�ڧO�[�.��{��!}!����|�N����@L�\��\���]�R��V�=�,-�/�MNӚ�K�����x� �R�ΫE;$(�ʎz�a�����G���
P�
��4Y�S�0S_Z��jч����7���XIa!i�V��k,;��a��=���[6��;T�t�������+�J�oa)u�*	��-@���֮1����7y�CJ=�EO%�y�ų3><����B�52(\�&T'9\5�+�c[׸�3�ГRX���9�!�ː��
�DϤ�&�:����d,��udz��j��~ˏ���z�}��㕾7`ܶ��hw`�Im��q�u���5���3�XP
�Y�"�mpvڛ@�{�����˦+:�smr����NB�GWj�}���>߶��K��d��g#;.L�N��/��rDLܢ��~1�4`|o���m���/���01�R�-07��#'?��{�{V�$�#�0p���j����
�:��bج��m����OfJ��ɷQ��l�F������_k�W*��Р�l�x11-�3�^��3�!��Ӥ���._oٺݫ���Ww�=K�>R�9N�E�]cCm KH����<��\B��h��Bc >�����\}��0.P�q��M�6m������	�ߕz������+݁S�DH|F������-�����y�ϗ�p�V7!����>v�I�k�Y?X�4��l�{hyb�ض�m��S����ƭ�x����t�l싵X�4Z��tIaC�e2�U2.p�^�xݞ���g��z'�RO��rO� ��Qd׷3�}�S'm2���ן[��}�aI���]0�UIm�zJ�g�����ZԎ��W&m�j�a+{�F���æ*�+���/�Ƒq8�77��5\%L�4���[�-���^��ގ���ua��ܱN�-����9�_�\K�lӅ
�t��/�R����mfv�l���V2�[�Ik��jV����U���Di5>v�N�g]�w1I�Yt,ӡN�]U�U�V}�6pj��G��c�waA�@� ��mV��Km]C;sX�6��8�y{�I8\[�e)��uׄj9"�&��O��iȀ���-$��������Ͼ��������:n�$[ߗi�X�r{
 �G�װ�sN�I;q�A+���!3%^����S�Ϻ��\�↻^��eXe5o���*��yaEܶ1J���֩v�6���u�����W����5(8��u�/��U2�V�[����ǳ~~%�?�U�\Z�؝�7��klJ���Q�Ԙ4����ڠ8.��n|/�)߳�kp~��|c�O��H�l�#�E�5u(�s��t$jZ�{����͠�a@C��_�=�F���׍��ک�[�h�m�mM�QN����4^�E�OR#:~(C�����S5��J�Dm���;�����3�3��e��yn�<�\6遢t{�R6&_�J� ���+ء�J����C������E���+n�2}��*��7�;Kz��ivӪ�h*�F|p`o����(L����F�`Y��mnE����-�%�_�Wsl:B�+מ���$%��y�{���⋈�"�p�V�F�u�
�\ԥߋ�C޼��Q�H�������ڢV���A�}��o����'/��|���۫K���z5�#`!o�>٧!8�n��g�>5�qTSL v��L`=0�=N�_d�uvI��cc`�ɱ�z������vm+����ʐ<��4�Wa�F�LTX.�j��>m_0��ھ��n�����c���R�X��ga��1�;�\�W#(Du;��PFby�<��������Y���;^G�g�dR�礔�l�T�=�Y/�6�TG��;�BP͛���Z�`i�nf���#sx���V!�Hӂ��q�Qi��P������5/�;˯�a^)�z�d�����C�Q�u��HB�d9Jgm:�Cp.P��>愨u�$wJ���W`��xt�_�&`V?(����u�)�����ɧ��ŧ�<i�yD6�nW:�s>�c=���,uɐ��ut=�,��f¢5;:�u7�	�=�1�c��ڑ<�sʅ�0�jF���c��'׋]��G��k~�4��F���1|? �@��]@q�Q|��S/��7��'z�2��i�X
5�>�B����[���m΅0�Q̣�Ƒ6a��IME�WH�k
����	q�c[ɳ�����r��a�s@H�l���%Ơ��Ư,��4�*�׮1������ /(�C�G>~����}�m2��vU[M��A����as��	���?
ȼ�A�^2����Q鮙*��H^t~�5�w-���z��X���/�2�! ۡu�x�� ���3���j�� �k�+"<�[%e�j�T��OJ4J3�x�5��'/�g*t݌'7��iov�f��h�ܙ�=�n��#����V�Y�\fb��1���
z��ft䬮#�ò�~����]��m��:ۘ�\�	m�!�c�נ^lZY�O�K5��=��tk9y+����r��BZ�K�n��Ȏ�"]=䈙��"b��ގ�fS4���)(�ltY�9,�g�C��dAj�Q�\	�/��K>�;��uj��&�5��
�a�f�UK��C)zJm�aG�'�|~y�H�5R�-+�o=1zr%�=��D7�H*�n_�:�}s�V�Z�:.�<f�V���v��U`�rCe:��e
��5�)�W1>P�>6`P]���AAO
�vq�T[�E`��kdL\��)?^%�3�H�*�,�a"��m�M�1��6�yp��k�����U��:f�3��[2k���*�vU�{hU������ke�c�0��{���**hɳ�xFg��8�Hz��^�5�۪����g�D�.s�Q^a�H���B	�Ui�o3(���	���N�x�:�ئ���G([�k��Jn�^1R��*K.72|ܣ"cg�v����`�Uoϰ�\�S)`�L�����x�/��}�u'��O#B�����V����Lw���EaW=Aݧ�y� �t-+�w��uđ>KCxsC�c�<��ν}�8@سhs)QPh��Thn@���ލ�eN��'ׂ�>F�h��Y�吶���b�3R̃+O1R��قd�5h�̛�aI���$��˪ }W�]\ŸکI�o���qRY1<�B�z{25Z)�Ԉ�G)����Myl[�NSQ
��'322a�w=���4a�-3��֣��_���kL>��y�o��3XuϤ)l	z@Y�D3n�l���-�
�b`�oq8�g�B�s=Ҫ�֮1�o����l1�j�*�[�w�o�>hA�9��zkUsLX�r���/\W������p����J���{W�g	x����3H3n��lv�*T��Ŋv��tly�t�*��5<��`
�N%��ry]vgn_{�́����ؖ}sB#��DB�'�6�f��;�2��g����q�ٮ�X�=o�m�(�hC�H"|L��q�hO@t�몈���d!�(��.n,|j�Q�26g�j@���4U�ydZ5�^7�/@�!���~��b4_}q
|��SC�.�/YՓvK���ɴ�6�	�Қk�=T��`�!4O�Rz	�W"qѷ�$bʈy�=�,�:/�X�?|���b�/~��8T�[zs&���E7r�Nw�@l�{$f�߲V�ïzǼ=�􁽘��*?n�e=���^�"�Go_ˋ�;��z�x��o�� 죶�^Sc%1���]%>�wB3rۂS3皺�r�5.^:i�4����hR�"��
F�N����Z	�����(�i��7�8a%<�Ĳ�h�Y��կ
q��]��+�4���׍�����w;��H�2
�/�����=�μq|�+m���RHu6_4��y-|��(J`w9�I̔+M����Q�0Q;�˔���������t�-��\�;5s��D�F�$��.̿Vm��q����N���YZ���^t쩍�P����]wG���m��Z��Mo���!$�qN�hgr�u)���`[Yy��\s���Ceg�a��C������Ye!�;�բ�d��P�Y�i�+�WLQ_����}���t�U��;Ҙ�Aj��W3�����U��b3�,j��N�&h�.���Ar���a��C�ר�[w�*��9>��.E�+�Dz�WR"�S~N۽���}�0�M��˱�s�Q�sp!6���Q�f�\:- ʛ1pڋB��V�g�<�/�H�j���˗���t���ù ΨDx���
�o]�u���6F�"p�ݖ
0�ں���/]ЮC�[��Wݽ}G�rZq^ĕ�LK����)VVQ��uj�u�yWL�ĥ�W
V�}�a���
W3v��T��2�V������;p��r�AX: �������S�s��s{:�mdM+:�m�A��Ý��ן~����{ztt�'�<vD�8ݻt�ӎ�t�p����o
�J�S�_60��Vt%_�5��`������3s���|:��ޚ.�td���kE+�1d�Af���YHp)fQʕ�����(������W]��ji�ћeҕv�k[)DxShZ��zf�Y}�}��6���Ш�E�ؽA�@��Y[
΀�\n�Gq�Ū�a��0�M�KS�h����2�!Ϻ���[ܝ+@��;,3wݡp频B��Q ugT���x룱Ql��kwL0%}Pf�{��A��2�@U�T_<�Շy��V���^��5鱚���IF�d�]��ni�ip7��rU��<w5��iD��K�i�۾�{y���]Zk��lt�x��N��.���6�BY�
]�ڙ�AM1�]��4��̺��̻ø:*��x�%�Y�)�dh^��^Qz,�9������_>��a�����l�[�+����m;��n��f�<�b��v	�XGLO�,/eԺ,� pW�o�1����������u�n>�*[|��9=������v������^s,s������nJcSa��*�w���D�<��ѫ62>�6u)ݏ�Y�(�U�z���2x��<�t�WS}ov��[xX]ؙ�1������N=�|��a�B�躕��E�qG��u-����j����u6)[�2��������q�y0k�wr��Cck�)CQ�|��W6x9�v�����jC�0�6iPhѧ�R��q�_y�W^�:��lV�o���[8�h��:�QB�ul��T��-�'�ooo_՛|M�E)���fr%�<N<x������5�ܶߗ���ܭ&�q�_.Z�P�N?���l�V��9l��6u6ެ�V�ݜ����Ǐo_-�7�c��RY���岴�QF��������Ns���ijmU��99g&urQY��soŷ���7&�Y�&$=��-�N�_m�ΣQZ�*�ަ�E�9m��$S;�rۻ�!凓wd�]�6�ǫ9g\��r۩��wlR��9eV��C�0� 0�"=Q��#_/v�t��@;�l��HΛ�Y�g܆m��[��,AՌ��@�Q']{�#R���x��bP�F\w�
DU��(�K%�UT*�S�@�ëU� ��F�����.���!����k��A�!ట�ȕ2˜!t�n�r�<m��w�;{d+�L9�ӘGB��ބ^e#^���lgh=\�<��]0=%tQ�i�'3F���X�h5m��u��cm=Æ���M
�ljxBn�d�,�G
��˽��'�8��c���y�yS��DW>��TsjP���8�r#�V�<�Z�=��Jn��%5C���Mj�е%�"�	�Trt��ȼ�נ�-��������6�:;ڥ�n��[m���,�R����b�X��E��aJ��d�Q��aC�X����E�Z�om�B��������m�΄J���y*ۗ��%���ˉ6/:3�S_F�S�&��V��7{�P��o���f���ە�]�s���C�Z���́fB̋O�8Ϸ�ֆ�N�H��/���ӷ�{�b[r��X��ry���uu�4��^HZ1�ڜ}���T�x�$�Y�W��b��_;�]C�^s4^�E����"z��@r���Z}.,���C��L~>���fks^a���v�;�Ya���?S�Kc�zZ����Ss:��vٻǰMP�d�(yzĀU��=/j:��u�u�Oj��:����%�H�3�x�=1�4-̼�7
�M��|H��ڊ;y� �jN��O5{�P��0`������t���͓ZhC|�L�~������p��"������C(_׺��7�˦�|�mۖ�ľ6Z��h�UϼT�IXi�1L1�Tz��G+�OC���R��ւ�~}y����Aiڣ��gʮ)�:Ezw�yP)Yf�	�i��;P��c��\��l)ܝ��Ϝ̡%�T0��H�{�W:��U����(u����cC&�(Zy�M��žۛ|y?���P�׿��k����xU��B@����y�Y��U��+��MU&t�٩yɻ����#uY{/���� KZ��|lc!��P/iSn��+%�q�3STå[r(0]j/ºy�8`ְm̓.3ҵ�z�(<@�B��YX�Z���z���]4c/4Җ�Mf�qX~�!y���S���Аz�}����B����<Qj"���8���Œ:�ȶ�� �1���hf]Wi�y���R�|�.�&�vM~��j�r��=fQu��܌_Loy��Kl,���A���m����G:s!���i�۴3��%�9S9�	n�a�-�7)��ttͶ�ԑ��0�3f��Oe�F��[qk��y׺�]���;��-5�wW<�xv��v�[Rv�����B,����K�K��O+�ȁ<c���i5A�@-B�ە��Mr��a�x��V��L�S~�r����ѱ��Lٲ�����ɼ��>`��3���I��kg��jh��A�a�ٔ����:<�D���%��mŗx��"�Wi�bA��\Kv��T�=��܃��N����SͧQ����X���`���)����=���֛&�DJ�i7���۷r�u8���"1�ATV�xq��(pD����$3�?�d=��r�_�����FFw���/1�PqށRXez�q@�	���.�k���㱢l^[}��َ���w�7�84qv�����>����!�%YT패vϠo�}�ؾw�b�JW)�M	�d�!�]�#�BH�����b�-C�����4��J�a11m��pG�Fd�Nn�!�b�o�%����mQ�E�3���OnH��Pδ����W?�y4^��*�����PEvU�Ʊ���9PL'����i֌8P&D��~�vI����w��>����\J�e����s���5N�k����7_\�s�]��ֹ�ը��~+(V�F��5b��u��J?Έ^��UL�ߞ
�ӏ��3^n�e��[�ۺ�1�5͍��2祑I��)��Fc�1�nW�N_�՗��nWjSk?C�� J-:�b�m\�����aݎ�ƭWܲ%.a��ù1+Wa��u�h*g/mz�X.,pv;.����P�K8�9�ޔ�]7J���
a��E�[Q���U���B���D{2P.X�7�]�zg_p�C"W3F�ʀ�7�QH�QCv��7��8�r�[ɳ�u=-�fm?`*|�+�X�58r�2�8V�mn�eb�<�m��i���3k�-|z�'� ��f6���S��2��{6�Պ�\6,U�V��{��ܺ��''���#�J<z�he�N̹�!��E���_ �5)�}%ﴖ�9��8�\+k���i)XjR�pD���,Ė�� ����������	���4�6��
��1E��c)mU�5�ÄZ�a~H�dp�a+`âW��UX�t�����z�xAk�١֭�n|k�P���e��%�P^�Gs��-j��,����y��3P��:���썹�5N��Z򃞸�R�M��uXҞ\���UU651��]�qj��Z�[��+����;F0�!����b�_�F@���c��g[�g����jK����)$�72?�M��lY���Wy�zÿ*+�>exe���;�sW��� �]����ؼn���X�k|����7Y���d�&��=90t����g��N���ƥRx�xM��L�l}�g�&@G�XC_�wl�xҏDz�d�`!g���1J��f�t>1��e����M�i��Y74�b��9ѮǎZֵ�A>ں�+���%�w1������Wp}�#\9u��C��׵/��Z�r��yEt�f xo7�*�Uxk�V��v�T3��3y����2���ϵ����󾆾�c�%6��D�'Θ}uB"[F9ap�T
��Y�Ru�`�L��*sLy�xKZ�J���C�JeH����X�G+�a#���bkϕ�r���[	�qJ1�������F��5�b%�z���v�)��jBm⮅c�^Ȫ��}�N�܍�.�.F;T��:�ȉl�e��X|A�.��	2����2�m��ybϽj2�m��)n�K��h���!���Cd�dݐ*8�u���*׀9��Ac�MSss٩�|x�-���ʚ'��jC�0����yj)� �r�&e�C��gd<����>�VN*�g����t�&����v���iv��o���t��xT����24GԾ��c�uqX���f��`dEj�x��Z.-ש�"�E�����J��*��G@��x������Ly͊��ʶ�q5��,��h��a9B(qU��K��g�>�c���J�*����V\ڣ�ln:�q�^9��^����7ga��ׅ*�L5�����`��kT�m�{��7@|��t�+~��'U�jw|A��eɐ�7ѣ*�}�D�p�x���iE:�؊������~Y�Ia0���}ݙ��u.�ĝj��5�Q�h��l�x Ludt�!�q�X��'�0�{m� �+f���g�g�0���/u�f�n�=`Ԡ/ʍ|{��e�� �~Ӊ�K[���;�[���]��V�F�~����é�^>_1��-�Ӑ���hG�豫��z4c�y5�t�n��ww9���9�r��$E�D��d>P����������F���򯩀�,���?k�;-����ά��"8�y���s���*�>%�B���Ft(T>^:c��;���5Y��7��GLc3�Y���Z��⫅VO���S��3����3�%H���'��xӶ��vI��Y���F?c�5�/�>M3*��7�;Mx�A��F]�4�X��n]:�װ��*��Ц�L�3w�@�Z=h�|U9��UUbDdqz��mׅͰ�Z���a��Q�c�sM��b{�cv�ؾ]F��D��j�yZK,�V�,���
��-����P�Z�t ɔ�v7�s4�Jj�[Z�r���9[>{�j����pڢD=��+�rFЈ��֜kg�l��Q�����⫀��q"�a�z���a�N��.�No�dO���S��~*hk>���쮼�>���m`�vތjJL*�h�ӹٱr��i�8�E�Fmo[ӐP?�*M����4���4��1��q�]��utݚ:� ��Ōt|.�ͨ�X\�-��\/2���'b�β�L�CU!NA�M]�f��U�\B]����7�hJf�'�蕓s���8cп����� �|o)a���T�8��T���E�㚨^ׂ����E�H-����&ˉ�)E\k��<�ך˃���[/<�k�>�!}<��;����*-DRp7s�P<��mU��&N�L��2����0�u���#\u4�z���)�O��]���KP&�XG��r����z�;Y!Y2���j��OR5 �뭴;Ux��xhO�rD�P%�W0�,ܦ���lf�m����J�$0�F<Ly�7R�ǜh������@�`-|"�橅�W�Us���B��G�����}I	ִXb�>����ͮ�p~�`?�Qu�� cW3�L��������s\K�j�ќF��2��2��Գ�d����1�/��Pਐ1U�j�W>W�:���k/AgCfr��sn=e�c���{k��Y���碲/9�S�S^3�N�q���ߞ��Gغ�z��4,�{𖀰�M\�~[�vM�͚K(�Է]�Bh�����Vp�)�L��ywΧ�,��~�?tku��U�$�Y��{_|X}y�M
��#�s�g�"r�3�;��Fh�3�.�C�>T���(gEp#J��)VL���Y�3�����L�E��'z��9�}SA�b�;�B��.�7m	�A̾ƚ֌�vm���81��d���w�T�R�j�СW�v�7%^�Ntd����:�H�OBy��P��f��~2��2˿���ۖɞ� �߱����ƞ�[�������)���� ���o���sd\O^d�n�R ��]yth�>�2%�����E�������מb�UDY�b��Ӱ�,��qQ���c�plꓯ~;2��j(��YB���L���E����X1�>��`F��=����O܍��|��{�~oN_}:�Z�}	��b���[B��Un��Y0­ݱj�q!�Ih��/�����,a훋c�8�r����t�h~�I�
�"VЫzUr0��"s��v��U�:�}�r�)�=��P��%�eՒh�h��F�`�V�)�?,�:��q���xu��Q�q��zUb���L[�sst�;�`�,��n�я)��6~�)��\���Bl��n���c��-��n����:���jR��B%�_� N�e|:SA1/@c�;��9����l�B�����jJ��V����5�1 s	[O�<t���P�`�������J�Nol$4�oe&��<n�V,
Y�}t)F댾RX-i�ײ����Q������d��u��3&�c��ཌ��';�`�~#}^��~m
����w�vd�^��v㾎�;ށ��k��B�*����|�U�v�S���wo�u����]պ>��<��J�B���N(�r�m���b=j�X��'����Dk���<���=#5�;����Z�����S0S튊e�қ��걸T�ȡj9��USk^��]���T��ٹ=��5�8ktT������Ɍr�f�ɶq�jz�\��ر�2�t���%��.n�QBa���39y�� �g�^e�>0�a�|;k78:��*�5�{l|�Y��hE3�ql�wT�Q�~���J�j��t���G1��u�i�}�@��W���۵�I��!�3���#�UZF	�*��Q�gO=0��t�?f���P2��ybm0�ʺ��*w��t�+��|m�ٖ��r�\�6בiu���<���ráݤ�x���%K���ތˌ��݃���c�!o@K�j�T�7UN���H��jlҮ�cߗcȪŕ틶�^�n��cƜ޲E(w�^w��l-�u=�`��zUcO�w*d�c�.�����2$f���M�����/����ȉ��7��ǗzkgnN�js�CH�Ar����g:Hй2�л�*;��n�co��6R�,1(̈��D>6��l�0.z�!��4�s�4r���<yb&^�ʾ��es�&ˡ�2J�g:�q?^[�9T�:*��u� {@՝�]Xe�;�sV��;N�5>��U�b�5��*=����x:ή�F!��D�o��ӑ����w����AP�Ȗ��9^��e˨�-�0p�U������uht��V�4�)�	u�n:��f|��W+υ@�%b~^���_R�x������S=7è�h�d>c/�sJ�>�)?w�=�uR���'��N����׫���Z�gf쉤:W[�S���dK)���	��Uo�F �9��u�c�_qP^<I��56��o}w��'^)3�q�%�0wr��s-�����)\5�q��4�*��0Yf]i�l�5��/o~DOZ�@g��h�FVQ}�uL��e����X���|��jK>V��1�m�F�C�����2�oF舏}�(p�5�Q�:.�j��2 ^Ho�~��Լ����lq�)�p�\�qA}K������BL�_��4?77����^<�	��0 '����s~���E^�F(��Mo�PT�ΰ�1eހ�t��K�x�%(!OR#:!��A��V'2ׁ)x�s������K�?Efö��>hi�����\�ZA�N�Ⱦ2��tD={�P��|b���]�?��=��H`�}z-`MƱ��A{��3��4�v����F]�4�U��a����,x;�5��Y����J�Z��t!�ʜ��dn�D��є�����eѭY� s�므]�J6o�c��[�������vZ�u��J�in�ns�t��V����wvv���WE�n���A=1E�dT�qWq���|
��T���R��*�+�G�K�wP���ڋR2���,rFI�;��FS���W��
�k])6K�Z���Aʹ��s���	�V
2���Y�CS�Z��ڻ9}���nsy�������.�.l�̫JԨ�����ݒ�������ࢍ��R��N�ܚ���(l�M�	��mh�K]
�	��2�X0]?Z�=��
p,�4��![}�93cc��[4��*�	0���4*�U�ss� �}���+�r�x�u�c6EH�w�2�5�J/a����7(�챔u��;�9(��䷄
�$Y�2@�AU�b���Ú:�$̎�'�2m�!?%�ׯ���Y\�B�]C��e�oX���Ӄ�0n�1�u:=����c��P��f,�qWe���b���ǧ1)v�nd��S�(Kxg9Nh
�Ӛ��ԩon1
M�2��
�����]_%7��_u���$����G���Lm����w`��pmp��n=5.�T���,��&�s3����m���l:9I��=<��YB���[�a\Ʉ�915��u__y�[��K�'(\��h1;�e��7t�B�*�ڬ��h��?5�մ��k�2-�˙��K�EE�_L���7��nb��*��wf0ɚ:�/ ®Ζ8�+N���y�nƪ���jQ�p��<����qף��S�Qdq��b�kkX��x�G��e.̷
�N��,�5/%��Z\[Q�'�2mJ���H%V�n>D����6��6�rm@qz�vK3�u��W�Ybܹ,1U�# �G����ᙒ�nC��I��f�u1�j��J�u+꘴�=�%J�]Nsx�cx���-hS wW¸����-�r���	2���azВ�ݧxw�ݙ�e-����EbQ.܆��;���%|7_o-��z���PY���MMn*U���г������{MFy[����5��weY�&�6s���Ʊ@�r�w��f�e���m��^�7���ʜہ�K0ː;\��b���]�t��2����{��ҕ+u�Sx��O�O�Ys�6�78�k�L�˲��,����2�-f=귊%zS����8J�u�Lh�/��m`I7��e%Ok��`��2F���⨕M�5}/{aC�"'b��m���k��p�3����F�
{���.�v�Z���K�ȓ�am�;���
��E��,�+l�yӅ@��)�EW*\E�&��!U͛nF�88�wl�sV|�&�{�1���`܊eg��Sg}t��rWIǧ�׷׏ϟq��ely6W��a�rLzM�5i;{~==���,��岱��ڮ��+7 ��r�Së�O<{x�������}��>�����V:�Qʱ�:�v��܎[��8��|{~?os>�p�޸g���wݹl+W-�gٷ,�w:�jܛjs�7�ԭ�vr�ߑ���VV;�[u������gR�wcwf�elu�6�|��{�ƪ7���竘K.�z�s�f��#�F=.u�ئjwrl�nM�峖k���ue91�3�e7WS7,����˻��J:�P�V.ȡ�ٛ���@��i��I�G!K���3���O^�����1�:�C�<t�?0f����u��ל�}_R�l�jS�+���M힛�a�ҫ��OT�b��f5�fSY��}�xD^�o߻�Y�Up`O_1�9R.�d�k�^���煮��2s�l�R�cu�ن%��+�l���\�|ޠ��]?q@K���9o½py榥b�*��;O�SM�W��c��I�tQ	�>���EVk� �[!����h���S��;UF����
w�ػ-�);j4�<®�p�a���e��9=�6����k*�]���6�ɋU�J�w�*�0Fi��!C'�,�/��ۻ���6�B*2���r�K�Ŵ:�l�ґt�ykB���d5@����P���B]�xd�]��#s9]1�E�O������K����3���u�[R����2H�y�\h� b���o�`N��-��L?B����J~����=����W��v�k�;u��$��w�]s��j�Q��zT��yJ��h����0f�A|d����	�Z���r�c����,�`������j_O\G�=���55�<��N�MW'���c��%�]K�GYۥ�j�ƣ�;m�`SǦi���͠%Y�X�shNCmk?u�G%�$V���.�Я��#aLhw;�uHiW"͂L���7g`/w�Qe��N�RXF-3�vA��}u\];7n�g!����T��g��
�>�t�}�;�(/C� Yʻ��2���J���.ֳ����^U��[��g+�Mm�1��^㾮a��3v�����(@�}eo�R=�j���[���� �xX��f�8v}���L�`�_;�kl��tԾ�d*�����{��U}�Xeid�QT���:N��E5�iW?N��$E�����g�h<�t�O$����ͽ3n��>��r�G�TO��^Cّu9)<4�k��MV�����;���1u�!�^�K����k��p�<��ጻ��G�"�"����XwFf
W/6��en���qL�Ǯ�A��j)>�YB��ۊ�!��9�a�_�-�I]��4����ێ�_�9�w���硓���5�x�&\����9����u{ߺAITd]/q��b�NשA�sS�rލnq��3���G�N1mٞ�m�L$�Ty -�x���Ǻ�^8��|_p�S�����Ǭ�A�[f���gv�5	r;Ύ���\3o�T�{��ެ�j�D��,t�d�aP��z�_��YBn���a��6Ar"T�}�v�y�+c��s���]�l%⻻����zfT��\�L�J��J��U
�'v�A�6�^��z�Z�n�7�A�3WbH�Jk��GkwZO���	Evj��f�Z���K81��옏;>G@@|3y��f{�-M}�,����ۥ��
T��X;[c�LV�H��I*>��)��"�r�U����;-�X�U�뻶��ٮ�T�G:^��^�L�>]hA��r����|�y����]j�xx�Q�;����]�ɤU�FW�ڮ`Q�ڐ�-w��,h+d����H�i�!��RżGDQ��Qljb�����gY�Z�����Q��� �+��y�'`��C�97�=�r�m�q[�����2|��^��.lTS)=E�\N���O�B�s=��A�]�+�h�a_K�8A�hk
��S^��kÕ!��L6��\�7��ܬ��q��s[���3v`0�|�؎�y�y�����<T��ҫ����Q�Γ��<P��EcaX��h=?t���D�~V��Y�B��dg3�ql�L��Ta�|�:}��g�&�y�Q�~���^��z�Ã�C��tc�;���\[M�O'b��C\�ZA�`�9M4'������>l����ᜨ�J�W?cZ��MF�Dc�G��sn�k�נ� ډ�ț�r�wz�X��v�Z���$��y���؀�yPx���p!��3oI�#�*��#M�ANk�\o���Gv���P˩�`�%��ZUQj���+96��͸�9}׉��K �&ށ���c�pXC��ﲄ��p\޻s�zv�:�(q6%���7�K�T�'j��[�TeO5	p�f�i������Ht�J6#R&�.ǐ�\5{}ߍ0V�Y���#�06�P��K3�j�k���(4���we+��P���K,4q�+����������3��^Ι�%c݈�����0V�4C�w�Rd1��9X#b@~v�ً��v��H��&��s��cu����x�&���/�2���^4k��깚��3��C*��]��ɉ�Aތ�tb$�aeT��Ī�kۊ�9ɋk��05�D�I��Y���g���7��l�Tںh����.;�iQO�Q��/���_��Z�`y�6��^�W5ZQ�} p`�[o6����9z�!�mm	�?nD��R[��LP�⫓�r]iQ#��,>�i\{����y��[��Q\��'mp|Ɇ��6�T�d�qQkkR�kN5�p*9�S4c�	�{R����}S��rj�c@ڥ�hf���Q��K�?	L���ޖ/{����;!��J��Ƥ���ْq{^3�i��V5ɮ]��P��B=�E�����;~��>G/��~��V�2���F�1��8�+s�9�騅ga	�S|�<�S�յ(����=kg%ָQ�@�p[Ck��ɗ7F*��4N�]����oG,G���n�V���e�N����`ֳ*��,b[��:a�Ht��:��f����*	X�7Ϫi:��O����b}\jZZ�!�\�C6�e��p�9�eUuT�w���_���J%���9�R:@bdck[�Yw�Ǩ`�f���'�b����m��:�nM�v�:+7y�+c�h`��֡.1(�fþ���7�ӷX/ ��,%�9 �T'%�|�q9�5����ygĝQ(c�=��At��c��sFf�ܵ�2�
�R2�1�k�Y�z��s�B��V���Sm��V���u����ϭ�5-Tdqx����t�SB���,�es\�Ȕ�ǳDfm�2�[�f�C���wd�S�����2g�~G0��=���Z଍W�ʺ-��J�QU�������A句�^6QYT��YZ�z�a�pˡ�����N��u�9r'
���y�7���1Y�
}����s������^Joʌ���;��h�O^�qn^����@N������26b�U~Z)ѽTe��}V����u�*�g�����o�W��D�Z�V�0�V�tπ����9�	E��!C'��}���O1 "��OE�m*�x��i��Q0����~^?Add�op������_��ka �:��ԍ�^��*���$ڸJk�}P�.�)K�״]��<�C�Fg]evX��e��]�4�����A͙\�I[ĪN�۵ys�9@@{��/Tz�	���.G[�y�>!��fl<nkX�ix1�>UІ��@����
�}�A�S�ƟU�S�r�m�7(�����v��7!��U/]�/��m�X0����4����%�?����"�R���ZEUn].�V5�w�ӡ�'Z�0Yg<x�<:��I#i]1^eτC?>ҘQ��W��.Nщ\�骳8p�6�F�.�"�0�c�����G)�>!�M��!����G3G��w��A�D>�.�[ë*%]=2���QC����q�W�gS�����K:Dj��|��Z����2�h�+��y�ʸ�6�t�V��;_I`6C�s^Y�f��B̚i���jBn�=�\oldz���Ut��\s��	U�pm>!���~�銬�lc"���\c]��/���|��b�Wh�g���щ�!�s���`^;^�[+]Bj�Ɣ���N�V9=�vfK��Q|(<%Tml������pwXw~���6yB<��{�Z.~4��H<-�u��ނ����7�qR�T�,���(A��-t�n缡�N���?_�f�������}��6I=�W�/E���,��靼:�uIC��5��+��'J�+�S�L�߶�Ὄ���Z0p��(4a�`��5\7vv�Fv���IXQA���I���mp��%��}*�k5���=2ow
�F�يd�8�&�&$?�y��v	��Ju���O�e�똦��׾�A������e
�f�Ko�\�?K��a��᲌9K���8�~����� y]����v�p)��Gs�eϚ������Nc�B��ʽ��������W�R�l����<le�P�����g\FN,��X�����ٻMhA�"*�1M+izC��g�(oj5�c븖��
���ru�k.���`.#]�a9�������ނ~�3nk�>��rƷ�LfLW?6[�x�e�U�����T��'Ĉ=�	�Ε�3���J�����*L(%R�����2��4o����|z�
�a|'/�ԁ���ꇚ�skݵ������A�ˣ�I�a�Wƌ8�"˅\��E�׎`��_��.��1���eO)T��%���lV֦#Z�c����E�c��6��Az���q�
��qAs\�>��2xEݓ�}���h�m��XC'����?0f�3��{����=~��S�;�[�	]C/�O<.��\2��������j�D���%e.�'ax���AΆN�6�o� u���1��<�x��O��q��s�Ř�)�C�k�M���w�NJf�y��T�����Y�Ft{�i��~Uh@h�J_J��[����/#���wsȺ�g#}�ݒ��n����a3v[S��Ӕ_
KX�u����=^�>��Z�b�:,���QZ��Wm��r���붋��`:sO>ԚHM�i�h�ϏBz��&׺6�����"$N��vM�XO�1�FBR;��ܘW}�W���<�v�j�8�V�I	UsP1R�껽4��n#�7`E	S��C5�Ϯ��-�7��v�vN"�&Fl��]�k�ZF		M�i��С;��u~���m3��]F.�����ݰ(ME����f��56�X��JeA�7^�X�G+�aөIm������-�]�k"e�Y�=�FB����5й�k�J���ݤJi�jBm�
�o	���m����~����&O����$t22�����#��U��߭�����~��	^�
i��z#M�5R:���C^��D�W\��T��uT�)>i�%��)4[ �^�n�%��M]vr-z�
��c�L���m����aEFd��xކW�M˶C�˞�&��%	���V͘�;V�*�D�n+�{��x���ؕ[m�8�ޓ9�@���Ϛ"�$΂昽�U�k����Zv,��&� �
�h=�QqA�*��nf��b~l*ǣ[E%!���3�ú�#.��R�J��-�+��^�ճ\���^��δB�{��d����}5��f���%�����Oo^�Ӱ�/F��R�<����[�̮����#�(���7�g���V&��Bh�Y+���( �ٜ�IwB��예/�S������e"�QoW�"@�Sو%�`Q#��	��[l�aV����q�Sc[c��qa����
��s	�z�e�vqYllr�CPN1�c�ֆ�����;Xz�t�_�n���׃����ٞt�u�Q��w*(|���៙cC�{���c��e��r#a�S�N��|����Y���lRh�x[#��P��hU������28�yy��w�3-�vjǼk�a�$*�B
���d��q�m�z�Hȩ1^�ƥ���ggs;�B	����� �VQ΅Ќl�^٭��#Pbdks_�ŗ{VH���+�\�I]p�K���O]�<��!4ɚ�n�hify�K�J(c�e���)۬�͔	iSp��w8�^�vOw�u�~�-P�V7�Z��'�9�,d��3&a�x˴�����>�M�ó��	�H_@��Y���`���,�c�(}�j)uʽ�O�x�O��1�'}�b�ɽ��,��N�W��_Vx�J���s�tF`_z�MY[|NT�*w�?S[���|��Hɳ�qLa����ާ-OҀ�Pt�jVb�e3#�e�{��x�X�{�x`0������6�e�F�e6r���%�����Z~̩Jϫ8��8�����m��qR��F�!ѱ$�7W�nGզ^Hv�.�l�A�O�_K�"�h�wǬ�9�n�ݔ�|���	�M�HHEQ��D�|.C&6�X����T���3爩���h}����z�g?-��>[�e�s3|&w������Y���s·�wE'\������=�%�6��F��ǫ�O �h��罞�p�~��{hF�FG�Q�%�I��ec�Fq9[�+U�0ƨ���W������5�������'��^C㲭p1�5sCrP[�b�^��ƭ5H���"6v�a�z�C)��H1�$K8H��[Tk��������T����d:��R�6xe��O��{���6�|9�T-5�?64�{�R7bIʲ(������^�j���ç��d���=;F=�v7T�yC�4a�*j{(��]�㨼%X�$ný��<�D���^td��əW���D��nu夺J��g)��F�B�Ϟ�r�9���p�i�l}���(�2���Y�������,�3�?5K��+��ϐ5�V����Z]Cg@��j�^��04ʋ�ǫ���-�Y��M��tz��<Hy|0Hu�k#�g���s؃�C��b��~0XL��<�i�B��f+_��7�����h.��ݛ�S4�A�Gtbd����A�P�B�&�Ue���Ghrr�ݱ�)}��j�X��	�HΦW:����S
��N�Tf���7*�������]A�P˝k�f7.��xc%��<VI=w������QC
��Y�z��r����{�x���M�ۥח�Y%��C %[O�Ga|� ��\�<PTEţPcw(ı�-@'ob"���q�=t�TV�$Rj�C�_#�v���Dj��GJ�k��m���t]���i�nM����2�"VZ��U�+,����*R�̎�Y�#�%�G��f�i�/�w�P
�+7�ë���gp�˴��bv�Jy]��l,	�<),��'M�t�s�L�PͬO�*�9l$��ڔ)CP�i���k�B�ƲW>���� �W*c�3H�_d07��[��y.�t�zf�p�6�ZџT�����J�ެ����mvU��I��;�7}Q=�ں�V孲Y�k�o��X45���Ok�yB1uB��kVu�:)������W[�T�W�%��֤���b��M��K�(W&J�HԬe^1ՠ4+���4Nɴ���j۾׬�9i0��v��]L�e��%W
�?��,�`R���M+�,͌H�#Au2��h�g��y�h.�G�\�A��&�h���Vu<h�M��vq�	8��!O;�����V�
�_\9Nۼ�I{]�\iZr�ʯFm�{zx�����ۇOI�ӎ8v�۱�8��:{&�tN���>�e��*�N�f�K��6�Z*�%��ڷ�M�E;ک��%;ƕu�F=T�;`�n��u���h2�fv�+{ٯ�wu��B��ŹqJ�讑��%�gx!U�E݁�72�%$��T��������7eD${���q$��¯E!�Э�.��5����tՅ�����]�̒��vQ�l�Cڗ5�×�GS3���g�F����<�m�ܶA��ʷ���oP�Л|/�/x�د���FHHl� ��@�:�=��$�E�e��x�ehQ;*�,6+�\�$o��8U��M����K.u�<��dn0pht1�bݹF�%Fk�ilt���^Y�ie�ý�0RegBYj.6���6%�ء�>zk��/b����67G\����aY��P¢]���,+ҷ��iC_��S�35<|  ��{�ҫOEo�_F�+f�n��0���δ�͹��/�;j� R��&N�۴�j�pӌm�;�鮆��оҹ���P��4���8��	���8���ʱZ��/�kW ���k�{�P� �T��,a1��w#o�Nܲ,���v	�h)Ҷ������P�\C�)Z���X.pT��l�]N= ;��Y�1n7�M!q`Jޤ�v��R��\"B|�S$*�w� -�6,����mK�W3A�&ţ�=A>rd���r1*rq�P�O#�)�C�H��
m��J��#�.q�rzq5�̭��7���(S+m'nߧ������|���wg�1��L�Sn��N=�x����m�m|���f�XܹmJ̦�Z�N:}}}}}|�m��ɷ,?&rm�n��\ͺ�P9fI�����~?6}�(ߙf܃��G��ܱՎE5
7��X�W9�K?:�7����rlz�=sl��Ef���,ua���,9�)��f���T�Σ�9u�>X�������f���q�c�[c�B��jl��Vw7-�SSV¨�9l�=�s&t�Um��i��N�8�N�=�=+}5��e���_R�իT8�H	�Y�ٷ�
��MLn���X��U��g�8�0�t% ���~��,@�SĽLU�ڹ����<��/��	_Jpm8\�o�Su�޼�q��g���5��^�l*W�v�R�-����'T��tll�F�/��/�[T%�Ec�ec���럇*�[Ò��s�Z��	�Ƚg����	h�i�WP� Sp����:�̋�NIO�.8�_nd&ZX�Ob�q��w&��=�rä�2�dK].��yFm�������I]S�j��wg�v��%�ہ�Q��&)�ꅏ~�tK���/زD�kSX��N�K��/��R�a��_y��wT�z���c�!� ��?�3����U��~��(�Qi͌YB���V�a�m+ЎQ�x����0�^C��h��x8�7X��3�ܳER�>r�;&�[c����݄r�Q+�4�=b���6�y2���B�T�|�Ϩ}�z��*h5��LXi���Zm�3c5t#K��,q�Q�J�Xۓ7�9���z,��}�P�*��J�u�~�ff8���ҫ^I��W��:�J*V��g�'���OK\X�S�ׯP� >7<-�l��N����+�63����S��2�h��,L9ڵ�[4n\�^ioQ��m�'�P�5yu���hN�B�,�����m<������m5�8Q%r��^[�����<��#�p̴�l�\�IО]�XvL��9m��p3�I\�;ӑ�˻��	\��U_ϥ�`��y�oRF)v�c��R1�=c�y��EP�4aŚS�
��<���aI�_G��G�|�́�5�����}����e��� ;�M�0S����~�C�[�ȵ�2�RXb�J�vU�����:�X�6~�(g�t)~� k�w�����E2�����!�w�b{�I|��Nu�%�Q|�&h����2�˺1�=x��!�6�?>m��D־��L]�e�EbW�]�����Z��ɋ���{M�~�Ӂ�??GU�*����aNT��4ϐ�s�����i�k�^��?(���֩3���,�8��i�UI��4:Ήg�.���a�_)obP�f�J��u����~PW�:��++�9s�]���t��`��BSl�KB�F�����[歝:.�VL{8<�j@Z�O�9ܪS���u���60�5�_���������X���1���������>`�T�4H���2��0],^��sK�M7`Je�����Ԅ��v32z֝��`�����O�=�"���T�߷�Ż�3[[XT�P��˂��|Z{�V2�B����_]����˻��eu�p��U�K(�̡��t(	jJ�S��y�5tp�'��d�V��|7�#�z�k� '��,%7dkH��sMf]|��]��F���F���7��_]�rA�ͮ�p���:b�c[��nf���o0f�3x3{�;Z�I)�y59�ڦ����{4���7!����<�D�f �h����z�����;�dݻݧ��jl��NM&ܲ�*��s�]6�^�u�
{��V�5�=���o&��vu�44�lR�΀�!���y��\��]0��Q��Щ^7_�g[��t>x��z�-0�x��j��̣�����/z��n`�gu?��R��r���1�Zʎm�
���D@��YC��� ��C-�1�*e�P(�u�DF��'m|��@�<ޝ�QB({��OaDsb�A	*����Ұ]E=�t瞛��8���aPV�"����i��r)H���F��r���MM���h ��:a7����]��@f͟<�H�!G�/-�d������n�l}���~��؃M�`�,S�ꅪ�5r������{���8.��ʅ��7�7܎\v�[�h���w��ڀ�����[Eʌ��~u�G���CK�@����>�.������G5��ysl�쀽!F���)	����vs����fh�x��/��5��mf�B��fkX�\�ٵ"�p��;���ܮU�4,��om�n���m�X^�3x�m��c�^'B��� �r!Gd��#F�7yխ�(vtN*��t0��M�$2��Z��"�q�_��>��V��=�,`wg��3y����%�Byd��yᛠ6�vsq�	Q�r���E�a�n��9�x��1�Zn���N-�)���9�^1��h����$�i���nW���4���ƽ�.�)�a;��$3k�y���0ua�L;d7�����y"����<`?��H�v�QLDy����>Ŏsu׽�i��g!���w��;_|���\B�|�$��oơ�9R*��y��KryC��0Ӷ��f�ש�[�g�p�s���\�M"�K��cw��T�7�P6��<JbX9�`���b�7�ּ���F��-@Ot�BN��t&\��)?_���aE��x�Ɔ�E��l���[?���R𷾳��x�#T�i���J1��)�q}�k�p*!�N�Vȫn��f:Z��Gqw�{�7Z��޹�z;>y�F0�Y����g�����5*�t@)E��� �|f�A�ge�#�3*�Kխ45�����7^�ܫ���|��)�P����w2<�a���ϫ��:b������0u�2�$b�c[h��*k��>0�d2c\�ɸ�	�ߣe�aO(�9�J��z�a���q�d���T=���B�{Z��/Ff�ǳ�~���(@��<<��=��ڹLֱݘ�R��@�Wo�ҭ�ƶ��*��yY�T���V��^N�Ѱ��-f��r�'�XU���7��c&V����-:���G�١��d�s�2{v���{���9Ϝ��ߺ�Ie8���m�dW:؛ݮ��3ǐ�ۙ"����Y�LZ�FO:������n��a�>0�e�ax��;��rk�ںu/6�^�NZ ��B��L0�l�Bz��O��O4��!��}�/��m P%s��u`�D�2�JukL�����<��/dKf���Rs"؅�gʪ��T3���$���#F�eM�݃cD�c��g)ݧϊC��~�y>F���4����y��e���s`�s׎�k�b��f��.��u\.�ʁ��hxвr�������7�=~i���ƫf�8P͜ٽ��E����.�	���%R�������￷�}����TRk.�e��gc��{(���B΍�upݬKP^B��v��Pq(�3�s�8�Ie���mQ0�!��I�~w�\�6��ym��W�k��c�k�d�͚��r�_�P�my�At�;��/�0��q��G P�l��g<7bz}�}�5\���`T���wSl+��ǡђD�ӽ���*�Q�.�aL��g�AY��qg]�Y|�;�Т%ݱ{o@*�4 ��)�}䡅8���d�1��,�^���+?p�ʺ2�����=؝c ����Jk�	�z3�^�����j�f�<󇷴˗��+}K<,`U��l����e�1�~��mR-)�v�<N|
�/)}�I+�%;�ٿ:�r��5�-;<�]�uj6�\w�f�'�&�v�H���^3��B�
�(0o3{ۆ����N���Nc��ݨa"���_��a�=���������V=�u6���N]6^\�FE��}C�}ȭ�V���T��u=B�V��|�g:��pD+܀CC�k�SD�ܪV+[?DZ�mJ�bd� ��X��O�|���&o&+�zW�.�ˮ=k3��V�MZ��5���t9�G�	��	��5)��)���y��R��Q��c-���N������9
P�M�0.zǒ����$_0�)�
2Y1<�|�)��)k�b��i<��j����Њ�HQ"��X���旃)��=��Ы�C���tTw>5P��NEYQwY�˦u�����oB�#�9���a�׼R"�H��S�[|޿r�C�#0�5����4��9���؋�/q���e���cA}.���g~2|�	���}W4�;v��O��q}g��̽�(��Lc[�5����w�$=��P��DF���9��d�@���RN�m;��d����k����c�N~�_���ޓ�yF{�Z!��G�˂�f��V�2�ǝ&+LÂ����C��l�p��1�
����kQ&�(���LԎ�WB�%����Ȥ��*�@������u{y�S�.��'N[u9��m";&�'���4 W��t��a�ݾ�suo�Q�vh�gf���@�V�.*'{Pϧ%k������m�6�����f �Q-#�6����B~�F�TO�=L�}Wg���xl���ä�P��9�:/0����le�A��iN�ގg��؁~����WݥG�޸�^�V��`��"��䷪EEn����fLsf�$M��2C+��s��oޜ6�-w>}�d��m�4Q��=����v�y�\�7����:���K���V�Ľ<O5����Lqƹ��kzl����՝Җߊ�ԲnA5j�+/F5�\	;�v�F�Ƨ�l�Y�C88��@|'u����@��5�2��C�s<GgF��v��3�y�3A"u_s^�Dr���Y]��ռݕ�>3E^s���8Djv�5��zR!��p��T[���Q^�W#2N�ب���X���63.�sQ�*��ř�n@X��1zlm���c�NCf(������K���kX2�$Z��������C��z'��1�4�O�Qv ����}%���%]qB(f�F4Ơ��s3���\�CP*�y0���E/"Pl�CBl�_E78�����ʛf��cO	$榌vi�ϛ=,*q����,�3i����?P҉[�;*hj�M�>}t:�"#Rͬ9Y��![�4��:�q����]�|I�q��ES�}�������曘C

���?�Pp���Ś��`d��_�g�m�j��˪zq�:��Y�4"���:�-���5��vv��ڜo�R"Ҙ�%�u���s�5��'g�^3FpD�������f����Wwҍi��W��\�1g#8�o1��{\i���X�|���`�wLu���PϙX�� �z�v{3v`��q�u����r��M.��c��Gs,�
�h������\�)9B�;R�zjSV���D��ࣁDd���[N���ǺŻ�b��_v'j�p�:z�bI����
ɩ�Y<.:ef�Pps6�����Y�V�n����3k7P�&�f�u�ϢgQ����v�� �U��)�)z"L���w釽��YB�m�oޱ�ٌ�{��F]����[
���(�r�st{�ղj*�M��^d�n���&K�𫭧U*�]JT\Ѫ�+X��O�=@�On������o��<�=�yG��G���Vh�Rm�ϰ��T�w8�䦪�`�]q#��F8���~� H/��m�՝~�oL���v~��S\�I�W���x�(�������G%���pݲZ_z{%�&�$ߵ�|ׅ5��!f�g\#R�"��r�p��y�X{Y�Ůk��)��O.ϧo�`����j2��C�n���1�7�a��P��x������1KM��ҍ1�aq[�Y��05i�`�W7K4�C��{]��#��<�I*��]<�WX	cCg\y���=7�z֢s���'���(��#���Tm����\�%ck�ڵ��£۵4�Z�<\�yחdv=�`p��"���oeA�ӧ��<�����<7zr��z5��ӼM�㏝p���2����g��WU�nF����Y��!#x{������?N֐�*�e�N���3����c���DЦ�ꀔz�v_N����ɣ'��zYՍ˞��aq��T�@�m3��� +83�K��/�d��f/�4�_�i�����/�Ʃ���eK�4F1�3(�\]�u�٩R���r� Q�re��9i�;)���D�%y���ݢ-l��+��/:���mn�� ����6�ۗ}}k5,�*�
�;0����UL���ц5ei���v���-��d��d/j�Z�V�n̉��S�޾m�H�/��J����S�LO�$d��n��vFY���v�d'��vV��m�t{\�O�T0&'g[C������x�jf�.���j��il�{���>����UC%���B*.8݅u�җ�;=u���Y'��Ǫ��#o#��vc(���&�Ϋ�䋑�C�����m��r�16�E�V�zfqH��M�+�9UEձ�o���"3�uŴ���,���n�vX7%6��g){L�� �����h��0�:�M,�ϰ�Ox���y�����e��7y.2�>O++�#K|!s�G>�J��m�Xz���s��>�K�T3^}K����-]�WqW��Wl�L5�w��X�Ty�f>>��G�pτ>�wK�{cר�qI�+�����7n�Jg4�g�Yz���h�6qَ��������Lvʽ�u.srX�ʔw��;���(݌��S����g.4�/��Be^b�K�vS�{p�s��M�ek�����ڼ���&On��I��ޮ3Y����@q��U�\.�� 竒l�|sx�}yy/��|iI���M�V/Z���f�u:ɥ^Z�3 j�&a�8s]����,x�p)��[�-���y�(<W�*3�&2M̠zŅ}:���gJL�9�Mt"�nT�j�@���yYC�����ΥӯHI�E�e��3a�ͮ�N��3+�\6���x��NWY]�|�T��Bl�D�:۰ҿ������*A�u�_�B��v�v1j���Gz�d!���:ŬD佚�ɖ1M�D�"�K%p8�\!�bM����!����f������[�8z�m
�.�ǎ(2sZk�{\*��:�N�Kw��N��et���
\��7� �N����F���x���v8R�0�����,��4��%eLB�;[�5�e^!���o ��m�EtjWT��`�۩Y���۠D+k����c�[��{��ҿ�Du jl��oc�ow4�g2�����.�wʮ������v�mLb�L�[]&a���teņ�{v��~�Ah�9���5�d�yܮ���M���+S��K;���;Mp�L��Qkܳ�}�������G��r������Zo�־F�cFwc�[�	,H�Æ�e�s��6c�
�<�����*�5gwaٖ������U�%t_l0N�f�`{$���P���� �Ã�:+��[�Q���9�a��W�ḑ��_)J.F��&J\���ŽK*�9͜�Y�V����d���x2�b�����CP�-�2%��;)��f�Ԏ��re�-񎫹��X ��fʜ:��� �Lȑ��PWcw�U)Q�qS�M^�Lӏ;�b[\��ͫ5�3Pt�;�Z�0����뛖>�w�L�V��y��lky��7K�H�1�CI�ӊ�٧$S��5׶���Æ"`(��X�]�u)�m��h��{��a`������syQ�3 u+�V��&��ꖟ_-tC��;y�O�5
��Lq���jx�^��Z�n
��˩cO]��彫�c��LSus4���p��k�L;��5&z*�[U����T����&��0���6fv֧���tq�*k`~��	����b��)NH�3�B]N��Y��ƍ 	JZ�*��%�a�k�[H;Ȼ��f�$�r�Z��n���bZ�P��k);��J���*���_Y�[Z���3*�@ȣ�vU�w1<7/i�h1n�e�7�9�]�=��[\+�b�����{�M9f����R�tKQ.��Օgz6C+6��O)H�kSh�[�l>��T�3kzZu��`	�p&v�)\�o��=ݩ���6n�Wx�����G�M��>��o^y��^u�^��F{�9mw�qjڶjQYF����������5�9��vr����f�m��r
�՜�$�����Ǐ�s�ܙ��X�S��mնVέ�#�EI��~?���qLVPUcVՔj��ղ~m;�YF��;x�����폜�VV|����m�������͜��7��%mw�ܰ�fVV��wu��KE�뛫jح�&��z���[wr>�ɶuF�g,�g&�F(j*��a&��v��m���ɶ�f�KeQ�y9m]͹e5g��ՙuuUV�^<�%�svl}aT��R���;�f;���#����`&q�n�8���C6bZ��u��W&��2y�xA`?0wp:qv�DĵGm~�u���̀=��oO����
3';�)��2r�+"�t��#m�ώW�ވ���2��}ŶCqa�\�d��md�v��Jk��t�C�#{�o��ƽ���1d?im:k�.[��ʺ�n��Sס��=D�x�w�_vm��G��٢��%�<{���1}���|N80��q��oc��3 �7s�iG�'#���O�Y��ź�_nA�L&���3w$�B����Vz�4{և�6�3�T����w�/����I� �s^e9U,��w�w[��s{L�yN���e⽒��R#:�Ԧ�Qx_f�l\��~�5f��#���$.��j"�Mv�.b��sR�"�\�j\�8,�:�^Nr|I
}F;9R��Ҳ����3Xlo6�Zl�MJ[�O=�[����T�/�^��=��#^*V�ɹ�5o�@�˚|�C�Kd
��)o���
�~܆T�NffǏgӳ���.]sǁ~��h�O�v�q����e���"9`vض�źoݵ7SzD�*�+r��U�.ImgT�?iT��r0��-��r�-�%^���v���o-_]i㵪�^#���-�{[��&�`μ�j^��?b:Q�QwG����T�+����j��|���'��%Sxzĸ�s����)��L�g�#Գ����,�����	e�>w�8�}��W�dZ��%��P��4���Q#:����mS���s�>�NŢDeHe��3w���+H~�k�#��vښ� �0Αa�1�~�4�������̤|@�_\s���������(��Wr�P�V��#Sf���rtM�=+�q��#�ƀ����α�)��n{�S@�fǟ��#P�=3�5
�8%�����l�ɏ>�i��e��״!<�pKd�㳐iTx�3��Y(`*�F+3v{�wa����8�B.�gU��~��%szgP�f[�q����EV1}��q������ k6Y��՘j8U��J�@�>//�]�e���<W*���J��'�cV�ma���#��Rw���u�\�t=�Y��6w;�_Ȇ�L��EݡC��P���s��ށUb��I����]h<Z�����`�Z��C��p�{��.fؽ��:Zm�����]�Y[��QE�W{�vt�����n���D�y �1�s�w��U��t�B�V/�H7�Ͳ�0qc�cN��
ٳ}-��;��đ�ҲJ�h�Ԏ�� �R"�j%�{�l�L	�8^�Kk+^���}ͲIHd�+iԎV��k-޳o��va�+әM��ghNI{Uq��R��
"ԝ*���/]�5�(]`��Gn��SN���Ԛ(���5�er����+/ږH�8�"k�
�cvUm��c�xiǫm��M5��\%_6.�����|+xEj3�'�M������R��S\�o�W[�D�i��7V#ta����tOYyY� $�<9ޱ�J6d3�� �r4�SfXi�C�۞�\��ں�3DI-o���c�R*����>vm;��،}�
}x��K����ޥ|d^��TϺ���\�%n��Z���Gc2�
u� k3l���X�;�_h�S�LB�`m��Em���in�.�t�O����<~R�kʰg�*v�E+4{W,��*ES���2֡�@�rD�rXv����:Dw8���{o�b��g!y6u^�&�״�䘤���U��iN2F����o�Iu�5�����Q�:}55������ڗ���y1�B�@Z�q�;BWL���^��'����ڍ¯w�w�q]%�9��D̒���Gӯ�<�n!�1{��C=�c��h�b��WH�ϳ�]�-��!��0Q^:���;�-K'�������A� �� �0�Iℶ7H��v��-����َ�)��N|4��q�4�@���;�_�\�B�3��ɞ�%�Q>�� ���n�������wW���ԫ�W���b*��+�Zc׼Ώ8��yV+��{��;�Z)�v�"iU]��،N/Pc�(����ȑ���@��Z*�t�$�U���*����y��+G[���!q���H���m�2��k��#��Vod<��xL�y��j���qۮ���8h���F��T�ẍ5OuY��a^LٷR/wW�5�D,�s�:�)���S:f��A��r���l�d�ސ�̟���Ԉ���o���O��o�����3A��x�!�!��3��oL�r�E^�Fd�hf�u��X"�x�]ݖ�
K�Wd�4����Q�O��`���s�|���%GAN">XF�K�^�<�1bU������7r��3���Cl'�V]L�L�b��[�>a�]�[��{�~+��4��P�U{����+eY͡-V�>�����a��wtr�ͣ�v{K��^�;�ZQ-w��4��'�	��v�4�ԫ�)������}����*�we`�V�z�W&�D��ޥ��D�i�Q}�%ۗ<����[5@%�����e��:|!��.��/Q�Rx��jWl,�K��A�rn���v�d����-#Z�d�|y�6���QЋI爜W{{��{x5f�B�8s���C��s���}Ŵq�=�$���iO,�w���}��]�x"�a��!��g��{׫<r��_�����Уt���'�{;��1��O}C3=�a_utk�W"{se���x��x������6l�y~0�2�~�C4��y�����&�S���_P�nQ�@�n����w�)���GChk�ݾ�)�f�g8�����e�_O���,2�R�fXO0�{3ަGr��-SnO�3�I�t�ci��)��֭�7x�\����Ê���_W_��<s�1�Tʹ�+3h���W'����
48��W(��:�خ��4��O���UL�j�v}BMW����O���!��zFDwM\Q%[��l�Z�&Zwx�d�d��[�"��lW.�J�ח[Ūw�l��}}�3_�Gw��3}R�9zN��u�wG]w �Ԡ�6����Ŏ��j�_T���b�5t�,�ж�g'<�#K����g�����T�K&ɚY���˗~�z�?ggWAJ�<�P�I���Ka��k�%`�[�M�NS��\n��~���LtlDn�S�7<��#�S@rO�zgsH䌆��72��Sl��^��������)W: ?nQ�d�j=Z�_X�W���±+8�މQ�1�.���:w�l���nOf�38���`p�~r�n��u���4]OR3ӼMw9�V��+��y>�cCgcf���(f��Y��1����#m��ȆZ�L�۝�*�1�\��ܧg�S@��h���!M׻#W�M:]��ȏ{��^#q��5������˲5�-���u���R���l�q�k%�'D�J~
�W2�J]G<���B�R��B�,�}[}�=ĀFȱ}*�-0��/����,3��U��B�ur�M�/��Fks2��y|7����X�3o������ˌ�F���5��zc���d��1��[C��^��g f��*��B�ބ9�p�ȿ[����Sr`,3��O���x1��S52aj��<���vn��7��Aԍ�w8�E�WP�EP�^Έ�<f��E�Ý�ݎq�f[�s.}3��Y��)��6䇌�5�Ǆ%�[���Yc,���x�n-*�~�#�
@�,�U�G�S��e��� �`�����v,U��s/����1ʧ�Jf���
"�!m:���㥬�)����l��o���9�1��ʫ�J��Բ�P*��U�Q���v����y�նuڝ��t�[D�_�5W�%#;Ï��߾�b�rV$��*���{�N���P�L��������e���i��iᒯ��w�M�ѯ�"���D���t����=ݽ@�\�t������[����[��x�6f-�N5tCn���B7��hyH��ULd`�;L��i[�2�@v	�l�s�sI����Q��Va6�n�9���#Y�F�5�|�b˕�V�t��Ү�i�@�-��}ƱDsj�9r�I���ʦ֦��vi�3���ə��u3R\�C�~���\
b��E��8{hs�R��so�D���щ[>���K�T�g�Ԩ�/<gy������>��6����+�1Iq� ��~.�"�d5���u	kԬ����:���ߪN��uqS֌(�.WG��%偋�O�����r��~��&�*��&��LAF�}ݛƴ�,�\)n�١�+zg5�v��u���(|a�D1S>��h���#Ob˾�z�|}��j#e��I�|fw�?`�i�H�l�6�@I���*�$2��#1��	��j�Һ�wa���h�%~�w ��28a�8����益w���z�#���\ђ�Wuy�ڈ��]�~V�jm�&|ǎ{^Z��]޼Z2��'�v' ����-H���`���4�7�I �%�G����}9q/T���'Gc��.�����A�͆�O�U��ሼ�bQ#'ǔ�������S]~�2��x��~*����%X;�kRQ�ڄ�g�q�㑭��,������v #%^/���tǷi*����5�e�ļ�'�����'J�T�_g�Ǖ�OY��X6���N�ٱ��Ŷ�-KY�s�vh�#�i͗?W���Kkw�,���C��j�=�ג� &�=��GL
�����l!M�)ڎ�nfk����(hD��}�v����}{��B~6%M ��qҮ&�n����8z;�7��m����|���u����'$���-wڸůL�YǴ�DTM�$�"���N�޾F�����S�ձ����I/`�P�73�p{��Ǻ��裫Ց�"�a��$��:���{[
���M.�Lq�����:qۋ=�ӏö�Os7��4��{��[�� ý�ٙ:F�1�x�J5����@�gL�(F���1�M"���,G'�t�����s����j׶�W>kd�fp+,��>�?{��3}����uځ7���މS��_�ռ�8�㘲�+Z[l�ρ���f�[��c�m�\��-Î��#"��<�����)KB1�M��i���]^v��{��绘����	S莚0_� ����&#L������']����~�z�F�̨��d�3��N��n���Qu�K3R*gn�FEhry���4��t�7�B��pQ�w�[y����1���Mb��Қ]��k���y��g��s�o��̀5.D� �7���\rr@okm#|v�Gk�cL����\��K�dX�J�U����D=oH�֬Z;۰�״�ZGv�bB&ۅnd)��ʳ�h���Ȋ��!�;^NBx ��Z,__c��m>/�j��T��;[�}pﴨ{�\�f���j�n<��0J�Dٺ�qWs��)�兦ww��]�7+���Z�3@�N�l�y;LW(������F��Uh�=LKE��dP�I)m++{�ז��4����7*��4����]]�jȌS+p���ޅ�܂��sM��R�{mX(bX!����Y�η<�i�����p����|�hwJ[�J�P	�R㎃��]f�L��i��c$3xa���,���pP/F#����*[��H�E�Yy����C�vm�ll�7ӽms��5Ӕ��e��}���з�π��gN�%��S5�a�����5/ ���8A�|�	�w9�B�uY��.��^kZ9oi퓁��B���0���NQ�ys0ˋ�<�H���w�=y3&<���h���V��b��fk���;��py`�M�ⴑ������͑T+�0�g�S-P,�!N�)x0WA��j3�fA5NV*���z��fv
�[Ƶ�ԥ��i���*���U�=�b�m&�d��:��S��<Ȥ�|�\�Z���
��Z�ɽ��_(�X�,Y��H��̓���ӻG��~�\*6/6�v?����>��^�+{Ӵ�]WM��};�v����k)���Zs~�%�{��U�D����%�o
��kzi�����M3��F�LPei�gfs�mj�'��6��r�;L�Җ.M���!݀���n��o���,��;Y7cMVҷR�\�%�<'!�a��&Yi+xأTv᎖B6�G}�`�ee���2j֓�(�,F�c��л{N(2U��%7�;$��q��[����V�k;hқF��Ľ|,mkmI�Ѵ�p���}%<z�g��+��(����7OP�I���M�W��_�7d�L@ɪ��ˣ�!0�&�	ŉ�����n���}ӻ���P]v����]OeJ��M 
���N�&:� p
�;�vxj腸�����m_4�p��uu��}�4t�lň`048�����:8�q��'i��8��È�R�J�R�YJ��2���+(p�*iV�HK���'2�7b�.A]Q.I���j�!��ٳr˾ڊ�.��ud���%w�1ȍ@*��n
�GB%F��f�ͣ�|���z���s�a�rX�c//���˂���X-�+��R��{\0ExU��q}ƹ!*Ңs��L;I&	k�n��'�Y��yB�0*y;j�����j�Е%���026��J�)�P��p��N^b����%M�L�)i�|:���xb����5K�vJ9�@�0:�XvvE{�\wm�Jf]
�Y�
m0-��r8��z^P��������t���>��R�7P6��,�}��z��<l]G����PcOS��P�ڹ;[6��?2z��=��L�q"�rb�K�>Ζ��*�һ�l��).C
 ���V�F��n9���ɕ������4uћ�OawL����L%��#܁#���q�؛��y�'b�)Y.�/0���M�֠��uU��>�8q�Z5�Rf:.���)�gu�ӝ2rY����!U�)�*K;�1��M��q�j��Rt�s9ghxI�]aڊ�&��̕�B���X/9�"rW	$���]��.�TW>U��ь�Z���9�B�9�	C��2�F�On8è)��0�C�0�<淲Ք����mJ*t6�<�7�LN9���l�Ԕ�R�M��A�*ڨ���V��P���P�Y�PQJ���V{q�nߏ����ϖ�.T(���~�޻�icSVV}��q��o�>����|��%���M�9�+圳>M�7�{{{{}}{>MT�)�5lU5j�~��mw��g床���q������{3�[P�;�/2T�R��L�er䭩��Ï8�Y����o.,�T�z�y�v���Um[z�)˗���������mX��J�5��#��خ�ܱ,��j�y����,����7%b�m�MU�j&jg�9\�J�UF��·!��>��R%�׮9���<O'Gi>=:=���������ٔ*R��ބ�oxSUݺ_WNq�*>C�.r����[Vl�V��]O��nF����4�S�����v�X�5(Ѱ}�hW�YN.f;Z^���ģ�|󸯏l����zk�o�z3�?��ʡ�
X�A�S�b�W]o|�;���\�'�5*�O38m��؇޸9{UY�عqc��_��W�
� 3 Wy�)� Wr�
+Н��}��[Dah�х���}�,�Y�F����]�\��3E5q�78�4U[�v��i��.����{+���)�>X�SC�f@�Q��;A��g���JU/[��:����~�ȘI��{\;��a3a�y�qt��[���:f���.U��һ���0����2�~Ep��h'�Re�9�gd̞�k������ܠK`�%J@/.|��-�>x�|��IѬY�\���@�{̼�f$[Dnb���Z
 �<����1��עħ�*3]�v�1��}���A8��1C�Z���Vq>��o���WAi��u'���	��{�v�pn>7ͪ�4�^�k �e�a�.���C��.�D3g����QcU�t*v�L1�	mm�uǑY����U�[v�oМ8�ɓ�8�H��8��k�E�xBWuoWR��-���lLTCv��8�@�;ܺ���7a��}����Rɧ�
�`��U��/�مy����e%9���v'r�ªn���]��@^xrF�&2��>���ދ���=ʲ�&���f[�-�Z�А� [����֎*uk\eD].�ٹ����L�� ��G�)e��+ȐwjC[�Mr�M�t,溛�ۊ�v�3;t�U��د�d	]YQۇη�S��a��J��OmO+�����-{|��q,�'���F�ξ��Ja�ѝNP�S��!�X��R�ؔ����lZ�v(�4Wq�t���xm��^Oj�%���[3���P��y�1�:��iEj�u��Fc�(�ߝ���cA�v�R�]����#���%�?�%���L����E�}[?F�/;NS�ȎYK:��78ۙ�`8��nh����$|6�VV{�["ྒ�k��2�Bts%tE',�N�G\w��:���[��:?��J�a���[t��/��1K�����z�O6ž�R�mr�]�H��.��r��z��-��Y#[�و�gi/�'z���(�
t	y���!�N��b�h�wuς��������J$�}\��9tz���^;~���o�́ w��
35�_��^'�P���]����?Y��jÀ���U
����c&��k�ø0nc��-X�\�D�1�*F`q���v�j$m�J��̦{����NSV�Wc�?S/ 5�=�15�@]^���DĢFF�Y=ƌ]S�0��ۻX��Ú�qM��v��h���p1Sꨵs�3/W�:0i�b�WmZ^�;����{~��X��:[Pf���z_��|��[8�
�J���:�%�M�A��v��G���)�C�/$WT,㩼e���ը�j�4wm�[͝�9�����͛>}�;��_�H�K�j��lU�|:&]�1z�����)�;s�ާ�d{�t��?Yh���Za^�+9�r.�5	��M{�t���g�"�a���ovԐ�@�D�f�U�4��'��ב
0�Ჶݯ��V�TTQ�}&�fc�[����̒l�=l]�޻j���.&Hz�|��ѳ�����] h�2{��w��ݱ�ˆ�ل�bP��z��2L�{{�]q�ko4��Ȏm��T���ϐ�ɼ�� 3^fW��*kz��5�|�(Չ�y��ͤϏ~ܪ6��o�X�z�#v	l�Hf�䟛��gd�3��gL>ù]��F�뺖 X�u��*`戗x�/�<���㺲�5�Z,k�o/�(����ݐ���2ו:wr�y�]L���Ҹ�+���D��z��7ݞ����f2���A��y>�PFd�!��V�����$6�&���MǛ}�f�����x��]�bSf�8�ȏ����k��/�ϯ�;�.�N��aч況������!��n��1j��c��Yr��+r}�7�tן������켘�S}��UQ|���2��g��]�!%"&�U�vS����7
��d��΂�ܡč�"�3i�W��Y�Ly�O�N�ق�ۺ��g5�p�8ʧ�w�f�XAIm�r�[����%�Պѻ�z0��On^����,�b�݈�
@7���R�\3z��m�n��'"L��&}��*Ǝ�c�ـ��P�Qk��]]]*���t(�˵�)�·ݺj�WI�m��JPvsx�]�QC��G�q�L���0֋Oq���r+���N�����%�L���yͲ���@jW��w^k�P�e���E���YC�4��v��.�W3j����[�h�ʌ�w��ݮzd4�2�w��ɲV{ Z��0�>.�����������w��vk$�m�������JW��KP��1#g�%� ["�=.��v��rMUb7bNs^2�������T���ά�s�g��z�y��SFnk�� �Y�r��k1�b���ff�[{}���Qy�Evp)_:/��Y�Ͱ[4�`�R����7s��gV�qj�4J��L<�+�m��s��U��e��:��D:�yQ��1N�b1Ȭ��+M	���:��|S�����[C^��z�����+����{�Ǯ�iY3���{�eY�s^)��eɸpFd�"E�3x�9��E���������u��I�F�u���!���j�5K�3L�w�/;��F����t�����p�ݗt�/
�����~?3`~��yD���iLr�芜ۥY�Wq��78�h�ϔ�h��cS��ĉ��T�Z� �R^���ZH��P.ɺ۾���{����Au�6s��O]>��h�)��`��Tja��z�sj&n_S�V�1we�Y���l�:dN��53U[����Ǭ�v��'���a��U�ȡݎO8�ɺ��t�;�4)�ޓdn�u�\[y*R˭vŏ���c���T�W$#�nU0���U�֔y�����-%!rc�V�㓇V8b��v}��՗�xq��y-J�,􈛙4��}���b���J9l�U}�Y��d��t+��E%����4��t�T�J�P(�ԝٚj�vwJ���{�:Hι�^���c���Ơ7CL�V����m�t���H`�ٙ��I��N+':�د׶
ͪcշn/���AM��Ҝ3ʃm�>��
�nx�K�i�VX(���4��,3"G��Hk�Ļ��9��'Z.��X�#p���[�J=��J�[6�J��(���\Tm8�z|1ݤ��N�aU�T�����S��\K$��w�k�g��b2�駨����mqT��@�ob��#��)�K��-S���Ry�,�:�c�x�x?N�{�c{��&z�z��f�c�㫘�1�VG+����͸���\�x�+����C>s���LV�d�k��e)�P۱�wj� �¥ǁ9Sy�y-�j(t���>U;�󥬭���@����qˍ�Jz�>�D��0�V�:��EGn�̓�����M���5�g4��8k�s��	����wȬ�y�ai�X3j#'6{xdk�4�K�il�F`�5���t��42S�q�m����O��H̽ܒ4ٲu_��S;<l�~���J���o�s�,���ԭ�Q�i�Xg���^��;_��Hզ}�Sω�};l���S��o����Q]�)e��e�6�+zr��v6N��>��P��V# on`���(���8��*�Q�QQ�^HXrۍ�_[6azpٯ֦&�V{�?�J���R?{׵�|���o? �%�m6_
��F���#9���l�Tz*���U�u��/�U��B�mͮ����R0Fb�]��L���.p4ܙ��x���^�#��Dz�.V��,��Y�#�E�8���G�ڱ��u/O[��N�_�)byg�!۰3�� ����7��^��ۣ#S5�穕����)u���X�_u2�G3)/5�0�;�ዄ�Hu)�4��#��?oL����ϻf][(�d5+����+����'�]�u*�(��*k2Ì]��������.�}���f�gK}X�j��t��0���w�����d}�|G�����!߲t���"w^/W����HWb����J��Dߖ�UO�*��%���� ��2��p�&b����ڝ���"��@�G�x�ퟏ��������{�P1�ͦ��1��z\Hʘg���mG�8c+rټ��H�,Ȇv��P�'�Q:���p�UQM�'�P����u��}[ې`
��v�S˸�9�+��Tջ��uP��E����Ře��,��ܮ{��9�ٚ��������p�S\z�It�x�<wm_�1൩����4{��+�lf1@�)�@U*��#�":���7���=��V��l��HE�^��5ph�,�KN�S]�v{���܄�&صj������V#�sQ�����p�FUܯy������@z"�f���lȀ�ȱ}�[-ݛA�g|'�H���K�Ԡr��]�[۾Z��l ؜��]�8Q
�믇Y�>SR���*���Μ'���[�
L���(ӫ�+ki�?_M<b�������sVe��Ӆa,�z�0�H�7(�0sF��޹���ϻ���tl�'f�HU�Kw��c������b
;*�]��Zt+��6�G<��v�݀��P1�	���z�8`�}�`B=pg����sf ק�����i4�\�!�.@h��E<Y��X�Oˣ^��x{�Ŧc�ј��k�A&^�m�=ʝmx�Y�~�����/��{�3�r�o�.���K<z3m9,�Q��{2�AKQ��<E��w�hX�/+�n�pvJu5>ԠT_O�B���C��Z��|��J���]�b��
S�9��9��]��I_K����Yxa�g��%���[�o?U=�f5fB�2f��;�A�j���E��C;���r]^�*���#�.2k%<�F�N���՝G�?go� ����QZ%Uϳ�2(�Ǚ�<�4?�Z���y����*������8�T�>��~�揽������B/��a���۝˳V�ө�m���1��y;���ec�ˠ	Y�	�/[n�d�9�.�SPsU��C�������z�)q�Rjt�������k�X(�`�"[�z��V^HH�As)��ߎ�������<�X]:�F���ؘ1��mP$)V��v���)�j�RU0=������x*��GV�L���y<��}ieqt�n6�ڗ�Dt�u��w�,�\��)���۾��5��.8�hEm�	���3|~j��pې�L�jU3����䯀:�J�5ϊ�����r螮��'�� ����9�b6�ܨ#��/c���)�;p.=��s�����z����Y
~4"�0��2��f�7i6ske�`�љ���sp5e�m�Ij���M=A��gc�����xҷZ��E�a�".Y��	E��Q�}�s��[R��R6�e�ޱs��g4	*�8���a���cع���ZP/2bsx���,�+*��K��/��z^�mu�ٺK��ѱ�^6-�U��.�EV�Xgw8��E��<��^Ev��~{���C�����Z��0��n����Q~��Զ�vqt�l��ڪ�@��$���:Mf{��&X��o�F�P�A�L�r�kx�9ɰ�.��[-�S���c� �*:�fX��^� n_�5Z�6�(�G/}��Q��UGqh{�g�++4R�1���m�F�fZV& ':��`�u�Q�_;��v�k�Z;�;�$r��ᓰtVVh�c��e�=�w�ʇ�c	�eǇ�&`�\���owf���H^�R�-h�M��#��)�v�\�#�;�dgxkN�x���lP�P��6�W]�tگ$�xҢ��ʺͤn��t�}���uk�6B� �PXc���4���;]�E�mS�JJ9զ�{e=<B.�)p�O�f���,D��y�����/*� o6�7R��ۈw�7Χ��ۮ��Tl��5mAb�^�Yק�涍��j��N�	;wõ�?�ޛ�� �ʪ�xl�5������Β;5�mF�!�,�ؼ�v�	�"z�Ө�*���2>Q��v��D�+�S���@��1�"�d�������(7�K���ĉv��:mot�'�J�X�i��qgfιbT��[}�&u��`����ՙ��\:�5|��	�K�b�d�+P�ew
VF��}֮A���)C�q޼��t[/Rx�RO�f�����@�av�P��1f)��X+���VA�p�}�F�.�&6�cn�W9��Y�ܧ�K���-:A\�]��%|V���X�׫q㷉e��H�Fs-)K{�]t�4Qr���P�qL�B-�p.H`�W*��lu�)�G�
���	G�Y#�z6�sK�k��N�Ď�Ẓ��G�1o/f��z���� ��������4�[96�C3`۸�K�3fV��t)��vrr�e�\[�pT�3��/C�a�.�*��M��y��ڧ�%i@�5�	��kMےҶ�\ܘ�Ļ�jE��Pܝp��Q\N�η���n,]�k���Ѧ���uм�r���P;Yy��v�-����m�s��K3&_@|�u��1$��}X	�J��Z�k�q�n\�J�z��"�㫆Jσŉ�y���F��sLfI-��'!��\��/*u�&��ǝ��d :w&�*Ò�om�ɛFv1��@�MJ��2�I����ˣ+h�	:m��ڶe+���f�f�����@u^��'S��]@�ٌ��x<�s�,"o6cG^RX5�$lt���
�B"�`N�Hvk̓�@$j.��4�t�¶�i2���:�;���*:�{&&$��*a�}��-�x�i�ݜ�>��8��%t��M;�[Ip-�yb�:P�Ne���^+3:���kb��a�c������/N�4ó�J�&��]���na�U9;�o8��]L�':)�2�,g�1k�:MjeẾ:iG��ss2��5�_/���}Ys�7�`l�!�f�S�؋j&��ޛsjC%p윌��wF���Ե�����;n�uM�Mn�S�p�3��w1�-T�o�;�Ƶ�}s�b2�&u'�Gc���q�18�n�[u�T������]��W555)�\�J�ܳ�WS+SoN8������=�,>��ʶt��J����9��d��q������~=�s���QO��i��[~\�SiV������<x��o�P��JR���m&����{���s6�ޞ:t����ǯs{�$��U�V�M��MJj�U+R�U��z�ow-�9�\��n-Z�TP����T�T��+)YI(�$�N��[�9ej�圶�W˔�Q%l�ʥ��niU�V^���U���շ5����Ԗ�y�V������MTι�J�ڕZ����G.X�j�VIZ���5e(�eej׷��������GU��#���۝˸;u��}���WT8�����MK�y�/O��>�2�����}_�*�s:���ȱ=_W�2o8>�����~��n=c�f��ʶZi��)��?D�ۑ|�^\=�Q[���<b�xK/�-�RegX� �:��2rR%dOD��,�c�,]pķXߊI�栻%t��(�jV~׆y���GK��÷�%?����9�s9P�\hH�}��@ə���F��9*  ��+X.�S;-z]LvC�3p��}*��~,��ֽݴ��3c�;6sX$�����1�`]��YL|9�_�6*�V曞�p�S>͇~֭�$m��\�~�[7^��4�Of�{Ey���Y
m��jڂ�5}:2�;��ߪ׺H<N�y]��*cg��A>���F4>�>���t�G,�/����=lP�«W@m$��KF���ho��Ng�FO��ͼ!���vD1�����n���$؀�����9t�gxE�Tض���_�)�h�{D@:���+SB��b�h7��e)(5�)�����Ea���������֯~�Ll6\�3X}w�w�ۇ7����\������7��h�=yq�{�Scap�ڑv�E���#��x~a�Y6J%ev�����TW����"&�P��/3sy�C��5�dfkR�]:�,���B/%�u6�x�f<�S�u_�]��_�����`f�oF��`��2Gw`��>]n��j8�1U!���:B�Wr9���V��3�%�=��B�՜�z�ڪ�ߡ���<ܣ���UW7u0U�T��ܹi#/�����]�;�R6�iʼJ��=�u>��t�pl�Q�#3dR��ٛK��Έ��=,-���g���J���Xǰ�ӣqv7Lƭ�1D�3EAl�|��96H
�Eqj��z�ʿW*�:2��+�u�%Ͷ�w[ȈR��p��E�igq/�d�M��-7�j6�oec�]���rus��eߏ�*r��{h�R$J~�Ux�X�@{����n�;�Zx��No�k���<�I����wHkdfpՌ!�igG/oL���H3�沾X�S$�֜wgWf��𱄅��>�ҺY9˚�bl��d�k�=|��zq��e�ur�y �U�+(��J���
�
7 ���0�I��A���vJO�G����k��1cY�m�p=Ɉ�6����3O=|fT�R�Β���U��v���$�ɞnV�g<\V�%(��W$�^?q�V�0�6�f�}���O��"�
�3��	���6^��w9���ἵm�Z�����Ӯ}k�S�J����n��7o:�9�6p����oF�U�mY~m�f���=n�p��;b3�#/�wQ� p�A�u6�A���fDfl_@�[-ݛ"���J��0��jh��؍V#������vXd^=
�?yT����K��1-V��7�C�`;�T[�_�:(Y4��^�n��o�����Q���=N�ǈ�G���cV�yv�W���j-x���ө-�^0����F�n̩��&�l�r2�ж���F3�B���
����x��7u�C�fѣ�8K>�`Wzf�j�a� ���5'�
��[��(U�����lhf8��Y��*�j�D�3 .�M�~�8�S\�L�a��h����л�x���ץ��v�]s�U�f�T��lp00��������6�b�*l��K=��S�h\c��w�R��K��t*4�����1���xxj��x����b��nY�b�Zn�]��d���bE��1VR�V�ُ�,�㹏��=yK����G�o;�w}��;՝4¯�oT��>k�亳�bj�B�1�m�wٹ{�sn\�tx�Gťf�8�+�޻yn��ئ��S���p�ٛ
���u,@JM w"@�7.4^{��d$���~��;7Y]=tl�ދ=;O�}o�=�wyK�\�>q���*���@��u�s�~;�Y����=�Y��%�Ҟ�x��:�՞}�)�ܲ�c��U�QF���H���/��������<f#R����޻�%s�8Ǣb�r[vz㠑�UZ�Έ~v��4�3Ӽ����� 6�@d��:��z���;�����������9��t�Ǡ��ޠ�#����Bbcd����CU;rٰy
"���GtM9�'[{Q�@�s�Fh�z�69�Pd�wh�[C=\FNձ����k�}�R���+�l�s�^��>*�̷�MV=7�2uX} �����z	�4�� 3d׬9�̖�xj�W2�J�6��R�[9sA���u����v��Iw3u�r�0k�c/����-�u�.=ۛsvۢ�ӏ��媥%a��o��Yy��4//}�P�=}�Qe��D���~��ӽ����A���x��x��-O^dF��
�s㬲BV����Zۥ��yޥ�O�ּ�3�5�He?��ꧽ�Kj�8�Q�jT��4��sZ��m:�;��:��H������q�^0�d��e��G��7m[ľW	K:w($���W�]S�bdDz���i���q� YnW(���f��p�:5�9����,�Smx⭠U�Pc���Q a��|Fl����ep��A�Z���*����	e���X,'�t,���,Ȑwk.��E�a�W��qkæ�O���!�v��R���iJ��ͱ� J�ˊg�r�m�j�vF]�-Q�gP�^�HW��I�T(�o4{���J�`�\�Sbu��ң ӯ�7ˀ|/>?��Y��2�иȸحИ���{��M�i��rnz�("�/eyx"�(ٍX����(c,�
[z\�>�M���6n�U�NC|�m��54a� �sk�v�g�<)o*�D�Y%uӷ���"��[h#�-y=�!`�|����!�X*�B��	�����2�0s�K�N���K���W,7SV�^�:�o�f�r�o	e�$��_�U�������.��Ϣf�'�K�}���-ۮ\z46O{6<����s��ss�*�l�wi�|�1+ה[���}ڭyg>�Kt��o��ּp���\y&p�0�hX�\���Ų���4����9���{Nh�D�3qa�ر9z���43!��&��� ��.��a <�{�w?W�h���]\����;����l6�}v�މ������CF�ݴx^qm~��t��*]��RE=#P�`�v�:e��nS�6�=��]6.����GbDhǛ�7�����.H�yA]O�~�6��̐� 1T��/��M��6�1���F�����Ӿ�����!G
G'�M�;<�z ~�{M��}_�庼��$�=���7CJ�
���-6�*/$WU�8�_r̮��ƅ��p軳,����K&��e���"ԙ}��t�{�T"l-�R���}[�����cSE����<�V��C���pe���N����ݖ��3�/��߭��wz���Z3���~�M�@^�߮��p������t$� Ⱥ�mZ{� �)D�����ǽX:�ʇeא�˙u�G*P��+ژr@�Q��ܟA����n�z��W�����g@�S�������3.⭔�[�sd�KdY|[Q�炣F>\p�OQwO�X_TT\�9l�9��5q=ޡ�-~���,����_X�W�*��t����HK��������+4!s���g��G��˞X��i��7����k���{�ng㫁]�&�嵳�4Pf��;�6�W8����:E�W$;�u(���n�OU�H��Y~H�Z�L�d6���8=kgT"׎x�}�2��6""������8��+�战��$���8{l�<�*�W�-���6%0/۝Y)����q�kl}�����BYላƃ�0/(9�z���3�]��z��Ѹ�����Rm���Y]�3ju5ִ�v�2s��<v�����ŕ�.�-sQ�i�n�F�J�x]�u���#��i��t3��=�|��<��/�����aFd�[�a&PQ���!c��8���Y8���3,���q���F5����≗��,&�6�CC��p��f���N�vʹ��m�[������zL���+��G@7n��P�/_\�]�FF���M�a!��V�72�5�G��x�v�d>`����@���k~�̺���>��&h��-p1S6�uce���ߧp����̶[�s��	L��GS��!A(愮r�]o�q�;u���sq��y�2}M����ʯ�E�����0r�}�.��Z����nݛw|�8��{7���C��>���N)a��{kӅ�!�@�~����:�<-�E�zyx��Ԫ��O�;��S�a�Y�G/lﯟ��D
պ�+w���>�zQT��rW�.�7��G.���9M��т�6���B��'����V�����^F�r�Gb�V.�I^����b'8�K�V��ه���_[� !�gЂ�s��#s�<��r�Z�:��Vf3u�wywS}k#{E3/1�����b�Ll{sP��\S�wZڷ���}}��5D��u�u�V�g3������?b`>�"5*����?~�U�S�b\�]�hxM+c鎛cӰ۳B ����қ�m���_�=^h�����n���Y�zVf�W7%�eg�i�X�	K�IX�˸���m(;����Q "�xE*�Fm[��=S]J˜@��|�S�u�|5T�Y���̓�_Ͼ���~Md0yr�1���r��95�w�c�����1�gה���v��gzy^�2r���N �
�X�0g$����-�wH�Ega�C,ly��g7���W���8v[�����Y�菰�f���-)6����u���w��������Ȅ���3�zGn6�� oP��!*R˩ݗ����v3�h>u�vv�Ve�j~K�c�>���"h�a�Ɍ�A\(�̰Pn،��{��o�z�����[Y�1[�Fw�Ti���~:�s��'��>�W��3���@Z�Op.�tf�(l��y�ޘe1~�/�]�!YO��1�~����w��O���O]�
���sj]�je��[U��5��HwV��P�����;�xwU{͝V5,�rM qVP*�xl�}Np��r*��7v���@����^��j�M�:��	 �<ld�zM,���a༃���㱛�&��{!'=[t��&�\o��R�e1�}H�H�`U�*�35%x���w�+c���@��6�Y^����gz�]�C��k��H��4sm�]���ܐ��㫁m�F��1n9���'E@�ӥ��TiΫ΁��o0Gv9#L��|�K�������=>�� YY k�����U��_��M{�`�՞E����?���A�ق4Ϯ�j{�}��=&V���;���W]WF�g��|0?J����­�s�M �Yڲ]g;-�B�>���*y���?��^�b�/MW-P{�c#��u�(�Ɩ���3���dBޟDC8kfz�XR�6g;W�')^�bD�\�G_��]>�������һkA+���ʊ���WʶO?��Ŗ8�ʵ͒�ϸ��{K�M[�ʊ��u�,��p��Vǜml�E*z7޲r۷/6z�[�0��\=V��}��m����pQ/�QB�=\��x�ux�z����᭵]�0#g=�x8ю8��㪃]�_���]�'�(��wm����A�Swr�n�!�^����V�iB=��0�xqO9��κ������������ͷ?��33o��o����ͫ���u���ޞ�m��i3g�lBl���[0B�L�նl��v���pm�-�!3��M�f[`B;��n�m�5-�!��0BfY�!l�5!����F�	�!3#`�0Jkm�,`��\Û`B�j[m�б��B�[0B!3:�:�S[`B%5�#0B��M�Ql!u��"��1d-�,dQ6%�B�L����d-�lMHd#�fJkfBlB�i�R�E$��Ǯ?����{3a��l��eV������?˫�~_���[���K|����O�(��`�>���bo�o���ϝ|~+e�ϯ��b�����@��5�G������~�����߃�� �m����?����9�o����l�o���?�&��<�����������X�o�~_�ٳ�u�����7?m���>o��������M��߾�7+����ffm����X�X��h��L"�i���h��f�d�X�������d�mkf�ƴm[F�[5P՛V5fi3Q�cZl�53Vf�٭a���ؓf��F���ٴ�

6�P0Q�"���`�`��+ccz&Ͷ�`�[+6�f
-��M�V��I�̑�m�����lĶ٩�klS	c%�"Y��
�Y�¶�k1f�dm2am��i�klX�[c���F͞����l����c33j�(m��m�?|�n����g��i�g�ܷ�����oC����W�M�?E�X6�޹����þ���n�??������^�`6m���o���ߧ��f�o��m��b���ï���f`m��}���6��[q���s��z:�5�������s�{���l�_��o��üͷ�o�7����?������o��ߚ?���~�́�m��������(+jڙX�V���Vj��VVژ��P�m���V�0�
0�
�
��2�mFڛ
mL��P5`Vm��¶�V�+0���m[m���b�
`�V�V�[l�VaF�j͊0�چVf�SaL��[a[6��
`�ء�m�m�lScS�(Ƭ
�
�)��+0��±���
�m[fڶ
يي6�͵b�5m�6ڰ+`�°j�+f���`��VaM�c�j�)��1FjmM�S1[6�mY�l�lژ(2���`Sm�cjf��j3(�S2�Sm�l+6�ͨ
��S6�
�+�Y�����j�m[aM��b����VlVm���ح��
6)�(e��fVي�5SP�[��3j3P�+ljm�5m����°)���՛�Y�ͩ���b�b���[cƣ+2�+m�f��Y�F̭��͔��a�1[j)�Jb��j�B�b�[(P��jڊڅb��S)�+j�+�b�[(VՊ�5+ef�M[SV�յ
j+jjjڶ�S+j�
SV+��L���)��V)�P�[V��(+jjյl��m�Y�V++V(V+)��b�YMB�[S(V(V++oݽ6�ٳ�����՟�?����Ѯo��������~�ogߺ>g�ͷ��|�߯�:tv�����{��g�����̛06����z[��������o�?۹��?����e5��4� 3��!�?���}����������H}��+l��M`lʑ%D�M`(h���(��BQT֪�UZ�g1�l6[Q�̶kM��>���ڵ�Mm���͛+ f��V�p�U]v��5M���R��k[3X�Vթ��m��ͭU�T��ʆ�UD��fi�6�c5(�l��m���Y�w���!=��������wW�8ΉF��1*�Ӻ�+�Nh���I�v�V�rZ�ml�j�m��^ ��JR�=�m��7a��v��p����ݕ��R3]��]�u��ݝE�9(ֶ�J�Mk� ��UU��`�]M�i�i;[MS���u��`u�[�%:9:AGnPD��Vη]���m�eor�u�Qwe:ۦ����]�4�v.��I�s�l��Z�YZ�JZ�en��x ̪�z��.N��w��gp�7j�.��gl�R���;2k�����Ye��mi�f���v�����Af�6��EwZ����Ɣ�p� �KF�9���
���.�͖mV���H��+�B��)ЗC�٦M� �6hh�v��hgXt��V���fց�w� 6�� R�\ uL@��t*�s�B@���7v��k  ���nt1L�j��K�w��yڠ
L� �f-��
���\!���� �vs��:��)�M�Kn�x ox4�7
�:�` L�ꁸ�C�p�]aB�dJ;��@ݺAC�� )@ ����J�  & L0 &O�I&�L�L ���` �{%*�       S����J        �"	���A�S!4�&M�Sd��F�&M�l���<�4F�fP�x���9uugfw�;i����ke�b�[�"e�_�`��/Ғ�&�D��P�?q�A�o��y�k~����^�S�s쑙  !:O"�~ED>J�%:4`A�9xe��1�`��ϻ�~rA3���]��7\���_����U�~�s+��Ҋ׳m����_�+��үU�9�hݙgX�r<Z%$��R� ���6��-:2<����d�T�T�i���nT���"d�h�+Ee�e	q�H���r��x7��EeJV�7X6V��f-�H�z����u�6�(]��]JK[���h��z�J��n�M v���Wwbݼ;��^72�5i�ڕ��^�p:�Ҙ1��l)�ek���i�Y���Ѭ��m�JV�њ�l�2���B��+��t�{��Qm��궭�J��+1JVH�@���̇e�Pi�(��fU���zR3b��SU)��Cdd�2D�kI��!ޒp\W{w�Fe�o�kU,������ԅ���/Hoz$�K�a(ó�z&�"����@��p÷� te�P��š�(!�wj����5���6�>V�=�ch���F�/H�Z�2�d��p7V@7c0k�U�R�B=�F���&��v,���k�ӳ�@�m�#�bd�b����A�+o.�q�q��+�K�wt�q��sd���W4-@��Îқ+-Д���Z"���va�Hռ�V�dX�F5���
�KHp�ab)VJ�e�
�5�%��Vf�Gi[F:��0H���$����Z�I!5�fCzz�k�V@�A��2Xt�Oj2Ռ���Xk1���Y�+Xve��un�*i+,P3R"�o���ݜ�� *��a�c.�ݵ���,�7��S����b��+�\ۈ#���֡X5��@�����夑f�V	�$�V�5�� �w��x!h����N�I���u�C24�Ud�Ly��K��r2�Z�p�2�VXB�Q��� Q1��iQ��w�I��n���k4kA��n�h�U�T�"�t٭׎�A�nCg룓C�1eғo+2Z��+���Ժ�7�GBk�F�z6����j������Rx��� �� ;M;ŹN=vL�1�)��uy���)����3b[�Ը^�r��	w&JG+fNl([ʉcڷg @���kY�T-��J�oTmV�U.��3NՌ$�xM�x��JH�!9YEܸ$�Z)�۫�kX����)�ӇZ{�;+{�.e�xO>I�øUһ;f��JZ�
���Nf����M�x���tܱghj�90�b�O��&)��s��m�%�YE��:�DY���9p-?YKF�{��m%KT�V#�2n�6�AV=J"�.�\�uϮ�J��#5�`�K4Vˊ����I�)R�$��oq1oU�k�f�ֳ{ XS8,= W����+,���v6刕t��t0��rJ��Sb�-�^�M�LG�.M��\��x��񽩆�f+z� A[�;U*nF�Vp&�)"t��[�D�:!5�jm���.�hw[*$uu�R+,'8VI�T��ݒ��X	�׍��F�a�Ƀ��S����ŵ���I�SrE�Yw�&*����V%=ej:��&�.�l�?X��:���l�A��jAk/*D������������(��ƌh�tV�x����汱Ę��5�A+D�VP$V.�"�f�s`��1�&L$cs,�5V^�ya9L�V��g�h4v j[+ʒ�M����4�D�a�BVᩥ����� *��<-��E�(��MW�Zvk��ٕ!���K5D!�js0�9J��w"h��{�E�Q�YOX�)���W����F�oj�.���[e^�%�{�#+�xƃL�Vdu�n�.I#�(�+Z�m���of҉J��ܫl�,E(٦�X����X��4A%Ln^�X�Р2Clڳ�F����2m�8^m����ā�q^ʒ���ͭ$U�2K����-6վĘ�PV	�j�um����S�qC���HwF���Z��,Zy�hK6���X���2)4���!��c-(�ݕ�E��(�_���Z+V�Ub�N���n��AXgL�㵖(R���ڣ�`
#t[g	��y�u���v(yx�I��qZj�n��z2����*�Ȓ:ձ�W�12V02]��3a]�ul�wd�4���:ȅ�G�8F<�*�T�;	p�8v!X�"���`�LA
���ױIX[�K͠��[��#
=6�IF��z*;�Y�����x2���e���ཌྷ*t�i�X~�u�U�0�ϰ���Jne�fk��ͦ�dԈM�FV���LJ���۹��mMoi�Қs"N�����:�̨��ؙzʣ�
�+���j Uܕ���U�a:y��H�{W�*BmLv��扗�m�V���ؕ���0Mx�3;��ڥxY*��	S�m�+nڎ�Fm�<̽�.�"u&���*�=F�C&}�>.U�j�6���j�c���`�W����M�ae
\H�V'y2���P�&Ӗ�S�hU�n�U#d�(a�̎�M�����#w`Т0eOa����0K���j���i���!C���ں6�B�e�3-� wf3��C�oq����P�#LH�Ml�,�"��OI�!��Ɩ(���3PT�H1�v�gF�َ�)�{R�:x�,�qX��s˩[V�̌f��1	!���ᬻ���]���R�i&��ј�.�S��SM�4_�h����Z�w&�=Ȍ;����B�A*<sSv����M3� �N�F��A�&Of��_�0�)WK9��PǸ3xv4e��^:��j��S$*]�efdLP�y�V:O6���a�C`Lbj� �E��
������/D�Dt��T��K?�PH�2��n|���' �wKǦE1���'�H4Ԣ�Y�[�P�4�Ub�li7�L('��柞���	��Q,ݷ��B��F:Ӥl-(������b�@��G��$D�I�Գ�YB��^�h��h��yDXqK�K��q������-]�t��fM���#��C�y���,�&S�Rɶ-ƅcG[�OouL˒�6쭊��́���6Btv���70B������TX��݀��V���
�Ϯ�J�VL���ب��`ȁA�zl\f���31�MV��5�@;��&���WX�٤��-�&���hJ�T�yٗ�FA1B
�,e7"��KN�c.��"w,I��vޙ�N���4m9��Ѧ��M�[�����l����؝��kN뭄�S$�L�i���I=�|�u�q���(l7 "���1؎2��#�S�H�V��a]�>�vKu-��FB���D5x`�i�,CvD�OV ���{P�X�ҭ�D�%/��*�Ei�	)�V�Ÿ���^F��V�l82^��/`w""-
��h�د)2	���-�*�����N�\���(��5�D�nB1�V�]�u五,[xi�X�t��*�BZ͆��n����YQ��j�f=C�Mdn��(�u�p=�K�����lac@�,V(wu��W��ԔTF-Rpi��aWSa��;:m��P+:0ٚ���7��e*�G�;��[Q��F�״�ˡ�Bg�!�-�Ym�]��T�"2�͛t��w]T��&�W�nǥ�*�R�G%���Y�J=�����9M��Yaǲ1N���뎕ݻP�!'�y0$�1GWz76�9Rڡ���ѡ�y�l�H�RH�h:���zhEZl��7[R�*,Zڏ8^"�U����B�O�JǸj
W/C�VhE�$p�oT*��j��x�CLT���x૩�A[�Q��tSp��jb�h]e�EA5��6��Tbe�OHմ�+��CE��aB�օښ6BqB#�׌��	>Вٔ��u��S���$ɂ�����[R��=+(��h�Y��v#��X���A����)����#�^�N��p,2���7�\"أ�!A�V��ɳq�ٸ�f�e�v�$��e��jK9;���<�1�V �8�k������m���[	�a�[�0�L�z��,�A�rm�%ع?L��V�6�oJ���j��򵑡-����S5�ٔv�ڔ �Q4խٍ���c��ءG��{d_��43��ئ�4k�#Gfb4MGIQ�����R��\Ecf��ҷ� �� �د��͍V���d�M�Z��-�&N��Z�g5���,��E.o�kkҪ��֛,��b��߬@�%eX��g5�}���^e)I�t��$�)�����)[X�[b ��[�V�J/ԱS���wb3N�u.�����@ad����Q�.��'�f�#�z(z��E���,;��Q雧#��
�y�wa�$`C]ֺS�u����\�Ql8i۝Z����_>� �Fm��N]�j�cm)7z�酉�����]
M��C���&��Q��֜3�n�Ғ�)"
���� �^9�bۼt)*���u������^�I�r$~k�Q�o�!H�mc9]��{��">�W`�]x �d��1&�c���� n���3nM��q���C���ܰn��=��R��$��^�@�iM�R=פ����ww-�����':Y���t��`&�l��n�̀�A�K{�K��/w�G�ȶ���[9Cyc���v�I��r&0�}������]�ExZm ,\Ag�K�P��tk0t���V��a:��8�Pa�4�d�h(�J��Յ\"8����>n�-RcJSj�es�Y�0cZz��כ&��Hr�\_>8)�1������wW@��Y�P�M�Z��j�έ��$]�c7�Ѐ➡������V�ST��}�n�B(sz�J���ޠ��(�7l���e�dP�y�:�dA��Z�H��N�-�d�iU���j�6-�́�c�Yz)��5���򖝥�iul��;�e�y*�D��]��n�%�i�z��OG!���2�h�x)g,�݌)[m�m8lyù:Sٳ��t!��(As��7��S����u<�j�oiN�4�\���R���y�r&�	 ��m۹��6������Z	��J�:T�h�Lj�ŕ��0�35�S�P=��p5}�fb�|��<���h�G``݆�i���o����-�U:�\@�N藫��r'(&c[�a����ޙZ!β>y�>(M�8�S(�=bI�
=@�5� y��ܑc0���%��ܤ	�J�Q�)���
����\CH]b�ѫqu@]�4;w��ɖFYq�X;%�֨�*��
T�W8�6>���/�JV�.��ݡ���j���d�g-�3f�4m�W+Bv.�K��8�U��+yT�n�r*W1��_:0�����
��V�����]���ݭ"IҞ�/H�d���@��ǎuA����!\e������oee�2Ң��XIs�q��G��7�S��U�m;�@���D� (�,�{�����n�d�mr������{T]wt]�2Ѭ����o���S@����*bdr�}:*ʭ���%�:����Fs0�m����q�_϶+Eu$Vݛ��$S]��=;x:���12sY.qX���v�������*X�\b1ruM����3��������^|MVz��'�@��7(Ԥ��3�tŊ[����z�m��I�X�#�7��ڹ�� �).̚1KȶG��u�*N��E������}jJ�Ɏ�=͢̱��C�m>*�,���Vl���EZ�0r�t4�<M��6dO��Z�C�i�@�w\6&�S:�u�L�%1����2�جcb���3�;�x���7j��e����U�r��{N�-�%��%p��ʒv%ѳ��O](���t��*�1p ��N�蔷t��nd�E'�r�:�J�b�i��,�Ư����m��͢p�ݺM�7':<jd"��~�F˗��:�zy�ay��Ի�lk�/��rb�	,�W}��m��d6f��_+yׯt�X`��x ��{vш+4\��,��Rcx.�*��|�=�f;���p���8���6�O-\�a-�lA{N�L��
Kf��u���9���1�Vk&×��q=��܇���Zח{P���ۖ��7���Cd���}n��}>�ح���>HkE�2��ͩu��o]�BSHW�HnN�і�58rȺ������Z�u���$N�Y�'t�a%\m^�VK���I�Y}�(�u�7&;m�tIj A[1A8���DN�yB�]k5�[([���SФ�$�p3�:���������P��hͦv'D܎�A�����u�X�C�g��S�)��:W hgQ�y׸���J��ꕇm���YZ��	�`}gf�)R��~�\��Y���"74�l΍�i�H�� V�M;.���!����+�a�Ů��Y���1����I����v껄��Pwp�,�Q�}rL] r�m^įx���Q_.�t����j�L�*/J�*m��X;X�������U���v�f��2	�p��Xy�s����(������ѥ�9��m��D��,�Pv6خ�B�l��Y�3���7�X�rÙWAn��N�D�	}B/)����6�3�K�x�(�[�Q��[@�٫ec� |#�O��E�cd�9K*uso]M��2�V9(�C��yy7��h�v<�Q�T�L�и�N����h��曈�:f<�^�bM���:/L�	ͧy8�����z��V�)\�彋��T�0�V�`�싫i^(ok��*�ee�ɷ�C�*��/����W\ϴ�,���hd :q״�crVM��ʽ�Dfu�EV�W�81gx����sn�q]����7E�t�36ЋS��˺F��X� �Y��C6��RB�����j�t��1X�4:�,WM������z��zf9�咊�ls��E��ʼ�[�Rhp��)j,&/>���րn8mG�����:��,�����V��z��v��iL�Ȕ���4�N�4�ҙ��1p�fPT�`N-�C����0\+Yy�\a�;�]#:���5�"�eY���PkfC�G������KQ�7��R�Ҧ� �r�c��P3p�&BLF��I��4Q-j��"���7���(��G��V�eƨ�/���sK3v�}�4u�jp�k�ie�N����Bn ��]���.gQ
���� j[;U�顁t6�[=��l{׼v1�|�N�[,�2�l�Rnp�y��\S��h�D/'F�K�G,�c�ξGQͥ�MG��"��b������t��.�xF���͝O�8�gu�+s�k7MH*RV�0q�(��ҟe=�/࡫�2�^Ɨq��2yKeN�%���+�i,�9�>�W�3|ͭ2a���o��bұk��|��=��7b/��/;�:YI��|JU{���'��Ffؙ6��㿐λG0�ʉu�]Ӂ�ʚSF���=�1
<����dC8!��m�j5�lo����:b�X�����if�D���v1�t����4��)�޺�Qb�TVcىS����tb������
�ޮ����W�>Z!B��}b�9�$q���;�a��j�Z��
e�m���I��<�ͽ�43��v��N�q�(]��Hr�s���y`��]	o![�y϶�Dͭ��]H�(M)1cĢ'y�y��`�ƭغU��CAd�CaB�G�G�:Zɕ����u{g{b�B;s�*�l��?;ؽ�K�o��\W8��bXFSސ�R���w���}L�ۦiHK�6�L�1�>�J�u�2����%���7#��"��ѝ�b1ή����[4�U���@--o6f����Q�S�h�&�P'�__��7FY�:�.�E���dL��c�U͡q�]o����� D⧔���X�YA���;	���\���F��G��.`�4墺������Ɔ����Ֆ�v�:U���;�+K焃��9�tt��FL�r�����s����8S�s�赪� D�i�!O])��mn���.�-j��`J�Y=$��`��m���[��0���K{m��x9����b�돕]es�[,w��/�Õ���SSZut!uu�!2+E)/�޷JT��ۂ¹T$��ٹ&����X�UxDKC�䜉�R�c��Z�F	L[��:���;�c�)���|~�T.��T+(�mrY+5I$�I$�I$�I$�I$���!1[�*K˜DY"(����_I$��(�*�(�n���Hc�Y*I-2��j����ٖZU5WF�o+�	!�RR�_,P�l���Tfx��"C�����������q*A�;pY���c{�#�KW��kUSqgj�m���w''�SKz�t�j�mlf�Ĺr�j^"jm�}rU髨���ãjgQ+7�ym�*��r�7A[�s�%�![�u펺}&�wl��bJN*'uqy2'��nC��6:t�W\�/�
W.�]f��+��|����b���G&��c�I�&gS��Y��Y� �D1�6��˙ĩQ�5���L�֫
�#7�� 2��V��#p̃��\z��E�Եi
����K�t�{�zw-Wa3ͥ��1v4V�:���|���&(A]����o�+ɴm��B���[)R�+�
�3��n/�l�4$m	���IZ\���ڳ9r���h�i4�HMj� �em�lڅ$_P�;�#���������毳�f��V���1�F�l���!�00M� ff����-lT!t"�j�h���m�7��ht�!^�G/N�����^�]j�prj��K!=����)W�.��Й������^ʖ�J�5ӱF�#*
���NB���������4�;�����L]͆�N�:�!��4�-re^S�Yxko)��F.��՗�C����	����|�'�;�f\D��-g$g!M�%�)K�N��]k���:��/H�D�Y�:vj��Y��ݤ���F'b�1r�@b7�/��u@���'N�l�ֳ+G [v8����^�Be�s�zf<}M���UѺ�QlP��X�n�5n���X�Q��6p%
줲��3z�:aaż���k����δYC��ǒ�LS�l`�}��5�w�MS5�E+k5���=x�θ�M�����q`�:�(6�nt7���1���@�ҁR��zRޙCx�F8R�U���Ly QdK[����&����A]ժ8L�և(1QH�k��®BL=(4+���f�Xq�g���6<��v��X�029�J�X����J���֌�\y��f�Ɛ�SX�0G��*uoR��^_}�)�9ͩ���������āl���G�4v��ұ��.�vC�d��X�|��n�Qroh��覮�o*�4}��8�� ��A���b0�KN�\gd��Y�м��|��U��f�<����X�@slWX��1�7�AE�n]g����B�]b���pd��*F��V�vݽc�� Ո�dJ;��5���\�9�o�t����s�"
/n��6���=��"�W!Ý�ڟ-��ȥB��-<�[���L�W!���qr8��W8-Ժ��Qs����ۃrZ���!�gj�_	c������� �U�
���k;rGN�/���7O]�l���	s6���X�(Y#(
b��ꇰ�� ��s�ݮK;Z���sN��%�+f�r���L`&ȳf0�{7R��c��o��@�q��g,�/@�n��]6�>]�ډkW�@�h�&�(���I(q�\Àݤ(=����Z���|�#ˍ������>����7�<��gU��l�;V)t�X��Lo,LD���VPF��\d����}�J�:j|i�W�(�	te��y��tEa�������7�֙ �޵p���-�����s����]�f_F8���}4Ń/bS��e�
���f�A�dy��:��dn��o�Q�V���#8�V����Z� '� #YN-Gw��������]j���{�A
���L�m���ٱwʊ��io��w@w}B��ȏI8��Pˑ̾�;�֯%��"��LsuN�[v�"�Tμ{Z�j@s�6�-�LY���6��^Y	�2@�က���3��ܺ��@�,�y��)���W4�x�p�ԃ<��WZ�B�����[\٠"=�i0鸹%�0T���S����[Ö �==r��wQN�p�u�ʹls��!��)���Ƹ�l Nxv(�{i`���׆p\�cz�ݪ��Յk�o�d�R���<�֬��  #���vF��k)�n.��R9���rJ�˦j�3��C���7.�,��֊�0cS�+���歊ڻ���dۨokh���ub���F���3���d��C]����n"[;J��3����k^�����C��pAK|5;HU�b�3)�#^LǓ_ K�7����FkV���;�����iB���Vh���C��R�'8*P&:�+�`������*ѺHb�2�M��Ï׼��-��y�ٸ=6��[ښ��K���A-��L�jn#xB|�.���躍���p,���+�����e��=8k�''B���-��E]"�*>��]�}yj)ӡ����0[�wN}|�r�X��l���P<��L�F�R;J�щ�z����뤹�7K�4���&�H�.x3U��r̠��Pe���G�.=��$U�G"�i]�CifW��ܵL��ږ��Y��h�|%�2r��V�í
tz��lޖ��A˺Q�LN����fZ�ؙhu��BF�뗶�%���8W1\~ռ���D����zvr:�Yv)�0��:�멆���E邎S���ᇋR}���C)�df��Tꑑ)�J�J�`�]�����.��tu����Fݽ��e8QT�{�_�3c�h�YH���+�+°��\��eP3:�n�f��ЈHkL<c&e�=�z�I�x��,Zzq��M|q�9X��㪲ٻ�B[��\�bV.�S
�)���~����MS�3{l&�Amw@;��9��7'��o8m�$������]yÊ?;Vw_c����D�IB\S�o��"�Ā&���0�N^&�e�L����0���vT׻����Qt��t�ī�c����.��b�C8uB�o�eW&��5,�in&r.�C���+�.dU���\.����]Amk������ё�K�wX� *�3r�qe8���C��y:e؜���WjwڪR�v�c��I�ּ�m�p��0�2FF�[x��J	�6�(d�5p�ۧR�$Ȼ��gG����]K[̕ ��f��{mr����s�n��gTJmDi�[���U���7B�C�Ytv��َ򇒻\#)��@`�
��Gg}�,	��]�����Z;�TtK���j�U�|%:����b\�Q�!�ͼ�уe�f��]�D����#.�ut��3C���ep�����G�KYr�i��JZ6�t:ܶX�*�9�(�*aE� ��f嚖��F�]֬ۗ�eh���;)S�_&���YO���`����]��W-y������BGݐtûVX��P3W(*W�ܴ[� ��Om�F�
�OȗB��FXߍ���)N�����j�G:���g������쳼� �h^-�k��ow\j���E�C�i:�I٦1�>��Nj����U��yR0�v<H��8�8�He���p0�Af���px�t�� ܲ6��3f3@f^dK��PTik!ɰ�KK+tu!j^�-[v�0� �e,�:�X:�k,)Zb�|�b�n�$�S�& �	nf+ ��6%�o{-��m�ւ�r���s�&VR��aG�ռ8��^&�`����nCd�Ls�pk�ŷZ��B�f+A�w�=Ntc.���<K�R�M�]�!3�ԧ��b��l�!5%1"���.x��o�+wk��H�d�宮��U,�$5 D�u��f�^8���@�l�`g��u�h��
I���2䐪5���� b�GiR|:���oo�jQ-rsf%�6�ݦ���)�ǩ^
��;t�@�yS���h���EnÒd�����w�#�N�+�T�0��v���G��=�+M���Gf96J:e��)؊�*ʹ1i��P5l���l�dv��v��j.�����휮��V���E�{�v3�X͖'Tqĝ-�q.�y�u*�tm^��@� �쉞�gt�3�wNu#I��%:W:��٧9�������2��I��5�F��n���;������Gv����h%��ql7n��kBt�fr�ns���V���ai��M�"�nZ5a���^���F�:!E*�����~ �\|7��AےsT����h�d_R�3���[H��;2e<�#-�Y1@պ�ը+2S�Mj�鞋�qFa��m#�>�R&h�3��׽�'��\V�ٶ�R�1�3����v�:���sEFm�n=g��~{��X۲3xJ�%Y�[6�E�N6����X$T�ܒ�t8��1�*���	F��4F��b��Ih �J�)-�v�uU��H\ݱ1�؀&*>O�P�ٕ�gt5y��p���%�]��6WVŹ�`C|>�=C5	G��gul�):X�����-2�ަ0�h����n�PJ#Z�>�6 P7�F�]`�G<s �E�B�wi΃m�a5��uc\��r��X���i|��*=YL�i�p��h�n����Ȳ�M�p�GZK|O���$�����A�j��ֶ0�4�<��`�H�-b�{����4��&�ѡ5�Cʃ��m�И�Z)��\ɤg�h6ڤ�F��I���(��K�(bJ�4:(����x��G%�*���i�
)�Ѧ�����
mf�+a<sRp�LGy�.5DH4�Ŧ�j�h(��Z���
H�H���h�E�D�8ڂ���}�ߋ����׻��<�s�`�:�)�����2͠�!ӵu5	Z�'������y �o��@(�ON����j� T� ;H�L4��D���ЧL� ��{���G�g�w�7��mok豪H��?p	AU����`3UY$�<���l�;�t��(!yȋR#�FOd�$�W7��;7���7c���+�Gȕ�L�G���8�췽;�9S�Ơ�~0s� U񧶸	p�7������z�f��u6����,�Am��~lT ?f?�jip��b�H�jo/�l��_��B�"���U�j4�DLq��:-P���oP�,T����qC��E�#����B�����&��c`b����=�G���R��9��A�j���cB��ih��#&=���OxrEE X*��j�tO1���� �B��jJǌc��fJu�.������lP�7(�+/�s���q0�+a$�䞴T�� QܿM�S)v+v��ׯ�+��֤�z���gqM��=�u�p��.4�Q�'!�T5CM���뛬Sխ��'\&d��AVժ����x�L��s�g���zh��~۩d�#�
Ҁ��;��A�j�)�,T��~I{�T-4�F��>4P�
����cld�$]mFO��^8�[�8<��_D-�-�:܄*$v'E, V)�y*�{'��p�|9Hy�F��&2ܓŨ�����2�kԛ��L��E5$��U
�"z�T�d-�L(�&ʼ��˴�94FU�ٱfn>F)�D�q�A*k��vĽaI7�/+�*�,PF�F�(��8�: ��^� ��SG�����~�ϱ�D���)�Rz�ŀ3(��Խᷩf^Y�2����04ј��'h3��| �%^*f՛Y�C��e�]��f˔� `��Ɯ(�5n�n��2}N,�y��{��Kj�b$��)E��=�$*�l�E�t�8h�r)a�s L��r਑�i�*|8AOJ��Gb��1��Cm*�GXٛ�����L��tG���+��!"hU��q���	\�����>��k��gC&�ܫ�x��a����W�UA�G���e;w�τ��P+P
��]���ʦ�Tv���]��D�j����؂�,�����$�5�}�����*H��]j3��X�G�j��qJ(���B)D�fH�J�cY�:�f���tŎ�*��C8���j���;Ǿ��� X�FBǉ�44��T?b�u����v�e��s�(��'Ѓe��p��T�mާ0�>�/���l_e�ó����9�@\�<Ro�*��@�v3� ;��l�ں5*ng`���%�S�D��n�D�}�-O�R�"q��b��+N��2�1!gO���DH��F��[�u�i����U�ˣ7F�\`CF txk5�@��T��x�Z����G�}��y�.*2���调�u�D���o{�甾�KK�@��U�xh~р#I��U�[���αbC���<~u�q����<��FęC��GAr#]�����m�\)8�l _mk�� p����,����9�S����^"jh�}m��t����?n��Ê4O�}���|=B����5Eg�@Ҭ�4o��D����Oz���g�b�a�gDUMT�-�4�����k���Zd���%��ayVi6�5�)̕����02-�����1���	&�,nh쑾DJz��v�OSzZE!��}���Ru�K�uh�}}^�u-f4*8��[t�����t���A���Eb�|��=ƳbCG!dԗ����k4��usQ���?*�P4��p��Y�Fi��xe^�����O���~QptL�����1X ���o�h�-�w�t����� Ѣ�xA8!l��,+K��q�8�i%�t�P0��	�=0Q�2(�/h�u/L��|j;�� =Ċ�����G�H�#j8��Aڶ��o��aD0���i��ĳ�AQ�N�z�NL�-��|�/����p\�+-�d�ƣܙ�yfc�t�����X�
(���+�>0�L�@Oƞ��ESf��{���J�iw�2�
�1��;B��<����v��.e<�ܓ������+�y�9���->Tj�>�#�"���u8V>B�қy-_M��A�X���H-�R��� ~�X�?f��d�A[nM�
�tW}Ƌ�O=8���8�2<h�K5Lq�W��=@�w��J08�<��c#���&B��aXɓ�y�[DofcH]�1�&Kq�f�ڎ2�Ս��68��@֥���a��>:��:򭳢���qzk,�N�d��rd�:)E����{�C��KU����j��tX4�δv�d].��찁�O�ANF���W#�ۨ����Z��j�<��Ǆ!��RO:�$}]�� �l�֪.��xzn�>�r���QF��Ϡ@g�uX�<���c�w2�R�lWK^ O2r_��3�#S)��W���0��<4� �0(Z���]N���o]'E�^ͱeog��c�������^�TǑ��QJ��bO�b���BEn�Δ3�Ft��øF�ʥ�M�$vGj���������}D��?V��Ȗ]���]����Wb/�����!�[�]������mv-"�@[G]��3f���>��46f"J�̃�vm7��"��UFE���E4���q/  �i��8�;��te��A��K!�
4���	��Cj猇S���[��;O��*�{�O�K�7���u�`cN����H^�w�����Hod�9��9,�Eh>���
xU� �Z|��������v���H,>��G]E����#{Nv������\9Ƙѿ4��CL�2��aY�q��]��j4_�<*��4����t���6+�{�G��Й�w�����9B���ok�	g�H7�;wF���s)�|�R#�hz%�;wh"���Ed/n�Lo��h�P���h��)lĞ<n��&)}`��u�ݕy�F��YE��%YY��Fʼ���:r�RD +I�i���m�݇8S�R�-�$XU;L�:~��<�f�E\AE#@���|�����El��2sI��n�B}t@���HnV�9<��bl{��d��!qj��u��B���3>��j(�7:�vf�k���"��xQ|�ep���<��QyEIY�S�B�4yms�]z�}.�^�J��Ƽu|!��U��R+�o�^w�^�Y=Pb�}~����H���i�9qp�7m�ja��=��3�:(N�-���s���_>�C �W��Z��_��2TJA�9�V�m>s��P�f#��osB�.b�*?bw����X8��|�Nc����kh�)̬�'�E�_�d�S�e�]x�A��7����7o<"�=�ZFWk q�>[V��>|1�a��ۼ�H��� �Ҝ�-�9@��dH8Vy�����2�>�~^
��b��U�~��l�V�Sg���}E�#�U7�����_Z3R8�A���<c�k�*G8=B^��%�Wn=Y1�1�5O����pv*C�7f!+7If<��M����k��i�o�([��-�(���PQ�V�'��L�����W:ۣ�' �c��mJY�魪�W�Ə���x\�a/^��q�*�y��R�S6a�j�f`�՗;x�;.�f��P����*����x���$��)�ƭZ�}�n�m��`�|%޺�m*��}Y����y�B	j�̀��ˣ�7[O��aT�퍦���r�FF��d�V��s��;��j�w9��K���4��&�xEy>KA�ڼ�˞
���*��wK����c�b]�TVsÖ��U<���Bj��=aCղ9����������"��Ї`��O�ԇ��nLd�Fz��|M�LM����U�oڭ����j�"����{u�m�/�ł�KQ�l	�['�?�� ~#��yz�?�em~��u�r-{�HI�Ւ�vf�H
�ò)�#�J�sPV��GՇ���
�:y���vծZ�sR;ʮpnJ��;�e)`�]n�5N��P���hƇu*���Ҵ���u�i�wKڨ7N �b��])�/kX�ʮ�����*�M���m�k�n7Eu���U��Y�zi S\�#dn��Q���b���[��'Rj�xy�aRp���w*Ws�.@�Θ ܻ=�1�0��FD��iq]\����>���V�Rw�����b9O.����v\p$���"��w˃�$v"�r�났�I�y�~95d�EVCH}�Df�u���&���(����桺���-��(��H�2JL���K��뷪m��I�5v��vne�f��2-�.�KG[ѕ�E֕�0v$3)���+��״_��� "��du�;gt���h�d۲r#ug��èZO+����6~��*��g5S�w�C�Y���
S�]ɷ}-R��ʷ��([�c��+��p]Va��vm��k7):5�d�r�Y,��sq
¦$R�`�`�x�u�։�Xڱ�X�h;d�ިx�7�n�Պ�ڂ@خU����Vf𝘩f�]�G�@�h\�^p\볮�򅜑�>�`n���$6��W���ۆ��v�p�ܚs�aw ������KԎ���R���葁�ѻ�%�\�.m�c��5w�n�`r|2^���#�)�A��8m���x)v;lT�Y4(���XM��*���7lW�&���Λ���8Z9LՉ���'T��pc����EZ)vgYi���d�65�!��D2�*�J�1Kq!r�:M��;Ok���\Mr��]��ε3,@ԍ��0ێ�t�j��������UL�9+\���Yܒ�EZ�WnW*|�ɻ\}�ׯ��;�����^��h�SXŝ�h�(��[:J(�N�����DS�AKBSE��f�q0U:hqM�Z� ��L��N�	��ڱA\����T\�Ҙ��kX�-�RFƫmT�Ad��l6�J���j�SN*��lJ�ih"4�Z()Л�1��͵TPwh�
���gQZ���Ѥ��cIAZJ�QTUv����
%���UQTA�-�V���]���L�1r��\�(��*�%.S�!����_}�����}��G�t����q�a9#͏3���)�S�|p_2}��C����܇ܧ��ǝ�^g����S����#�{��G�_q�K��!̈́=ǩ�' y�|#�� ����>�p>v�Dm�<�ߏ>|�=����c�D��{����>�_r���C���� �%=ϙm�? <~�>�P���~�^��8t�����O�g�����_Y�d~���0%�>�(~����S����@�H����<~��|}����6��
�̞�0���'b�9��|����Or��{��p��8���D� ����^���? H�_�{�R'�|��C��O2�d�/�����'/���d)~K���H�y�׺'���?�ď����#�}_H|�ԅ"z��y+����!ϼ`>��<aR|������C�av}��Dg�=�o�_��~���~~{��^z�o0~N�*��v�X�$�s��t��H�f�:�<�������
�J����P�m{��s� ��(����;��7D�9TK���w.��.ā{\�hxn)�~�O ƴ��fwّpu�1�p��
�	�GxX��%�ǋHv��O���ێf:Yw9Lju���㤆)%EG������YT/��~�5㙾<^�퍧����hE��ˌ�6'K��Fyc8'x���ͧS���f2������˷S�tWӎ����[��;��%��UV�<�{ۻ��D��O�u� :���Y�-��i`K���Ǻv)um���O�7�7��o-Ǖ9�����@x�xp����:��㳑:�\|kd�ocIa�9�5ڗU@|�+˱��!�]%j��yg�"�T묋Ƽ)!���q�m:C�>�+�z����˦)�r��Q��y�`��uj�7y���V��4����w3_�m��[��~��.U�KF=�KQ'wN��%(w��+𫕍!�Y�+�|��Ƀ�S���ԏ:�>�v��E��/O^{3��ſ@���#��)O
Z��;wo�o�a�}�-��]�ЗO��-K�k%L���!�
�\=V�������ER}KK]���s�͓ݓ��q;*�^:P~y'��T���+��I�또���n�9ш��������xz�[��@1�Eeh�C}�{�� �'���"Hﴷ�ôVh{!K�S#�C�Rd����o(�r��������r̗���͎�F�8h�a%C�qp�P����/Gn�B�B�=�tm�O��'}S�˦w�@H�k�d����}���r��z/�EH����d@��O�3ٖg��j��9����g��d^�c��[�A�;��U�M��<�C���6���`��}#zҜsڗZ������J�5U�����.���C�O��w�(ƭZ;�{ݽ��_�~�����3��~?g���(+>Z��m�pzk�-u�O/����݉�5{j%�ڜW:ݿz�67���+O�߲ҫ�d�3�*�ֱ�������[����TF_v�C*F־�9u�:l�3*z�W�iٷ�0B=}eD����cp�9�8�t�"��T������pwJ���;��M�5�uu˅�\�8﫣��oJ�u�<���
�8��Wy�o��G�j�S\V�{����� +ްǾ���C2��µ3ڟjlY�ٍ��3���"WMf�v��m��ű���:�����L�'V�a�^���J��)B�f7��~�o�;��7"���'�������X�O=ғs�N��N�4���H�T7(�E����:�]op�}�l�q}�(��,i{�Y/�wm��9�/R���?r���o&f�m�V*]$.�zR�8�/k�x�#'fJWj]fĲ�ugh�l?�iM/s�q��C�b��Z?gt�?d�ƀ��V�w@�w�nD���� ���yf��5��I�U�9�pk%���b�]�{�<Z;������/o�_죫{�U3ij��\bƧ������ki�wfj�ĭ∞��43���$+���������⽯�/9�n�Q�[D�t���a������w��S�t1k�s�gz�#�ȍ�����Zru訿��0zo��^���Wx�����hl[�e�`!�@�H4R;��Ov#�cի��o�Pʆx������Ai�ɄQʁ@7<9<h���U�	'�||�{��]��Y-k��jC\�aݐ{��l#�����n��f$�Ժ�m����!��Tof��eѡ�v�?�/)�(Ϡ��jS��x��G�E�R���;'T��[f���X)�$Sȫ��J:W�*��$�������j�?sڴ���0<<���8<a�Х�u�i�:Χ�7�~��3xO�/"1wxZ��U�V@�}׾b;sh��w�k��F�x���ԐV#�.R/��I1�;_���;����B�'��;���/w^�Ԋ�z�{5e�@�m�E�H^��'����IТ-�CJG�q��δ�Wr���W*wÚ�BF��EN̪i��.�26�[��n�\ѽV-m�Nʛә��e���҃���M�]�]��˳���p��*$<],�/��k7;���\�Ib�+�&+��u�n����Y��b�:2e���n��;���7�i��;����W��y���~�w�����i��}]|�H[��E�E'�!��(���s��t�Z�DzȪ�h\�s>D1H�Z��i?X���o�y����L���YbU/v���rqj����l~�V������Er�����\�^ G9��
ޗac�E�Y����X�R˾w���Z���Ϟ�6=%���I�H��z9AW����'�2�.S������:�Hj��T�I�`{Z�{�yI`��s�O�8�l<�S�]����B�՝���V���f���&�X�գQ����5P|K�x[��;a��d�b���4��ʆݓ�s-���1�	���U5�| )�������ٯ�h?-�>���v�o�/T��>���h�� ��i���ʇ���:�h���^;Cy���Ǳ�l
������1|�K�)���<���{���>���ұ"�Izr!H^��5�W�\BR���D�%�w�u����=�L����ؽ~�"ӕ�K9<��_{�U����[�1;j�S��P�� F�`V)k6�'Sr]���s�N<�;گw$Z����O>G/��f�5({W��2��N���:*����gr�DR+��ss���|�#{��uL�J�C!�##���9���$)���dY��%O��XzvΒ8X`n����a-1�##b� ���HS�yNa%k9JV�gE��ř��W��^~Ɍ��[�j6�u����^嶒��v���f���֪����{:jc����&�l���rQ��@�\(Z+n�ͻ|��u�7Q���9W0�ڮ�P��%u��Iz��&V���������=����'1	�
��:3�MI�*���rS�l�UyeGτ��[
^|�{Wv+���y�6߲V�A���+�{�E5�������q:�:���(?9�P��o��o�{����g�E�,��U�Đ�Ъصf����ʕˆ�;o��r�4�AX�]�7��,�[�&4�	�V)�H�sl����i�Xc�KY�����1*YPoKW6_Gh[Gw���1���Yv#׷�d�u�wХ��U�g��鴚�tVl���O
��5�F�
�tN�_#�x�"đ���/U���&������	���
\�;�e�΄c�tޥ���n��u5F�5��S�z����Q��ʎ�̿��jڨ��n���W�]VZO�,�_���Wmy�Khu� L������*��7���	����ţa�[�_lc7zڨҲVe�6����)[M#V�{]�����_D9'h>����8��j@U�,�w�!:�N#d����{���kQ}�ʾ ��"�bvݼ�aR����9w�f����ܚ��a��K�B��VhQNw�5Ӹ�i�r������V���2��C�^�O|4�v߼n���+&�O��[zw�7�������.b�X����=\N������Y�jv7�M-���ɚnqqÒ��	�a��C�졅�ّ[dRw	��F�.��	$�|f��_
�Y�|lr=�"�.T���n7�s8���u�g_Q�K�m�W���o�د�E͟�-!��Jx����m��lE�H��fp��;�&ǖ��m!�kN��չb���p���(�-IE�Ux"Q�_H���Na�]�=�0\��Xy\p�����p��7��u=�5�a%PH�֪���
�̾bhp���L�۷`ʗ�zȋ�,:k�A��A��ɋA�����{Z->��;Ij*�V�W��3񵇪
N��|c��h6Lj��8���L�9��l��Oo�1+���_<�����>����j֌��ٽ�*�⪠Ӣv�a�((b"bLci�b�'.Z&I�[��MPA!V�*ihbh�����J�nm͂b��K��#��֊�&"i"()����.PQ1DV�D��A����#gSD�40�PT�&ئ+lMDLs�9�S1�ME]ژ��;*Jb��sSQIDIQTLAZ�M4�UDMD��DQCMESSQ�T9���C���rV�%���#f�@ܸq9}F�6�w��+5�~õ���_}_U �)?�[W�=�����P7��&3�ä�t _���J�pt�x{a�t�KUei�k��4��X���ι�W�gF��6w��ݼ��������@w��� Qo��M�s�LN�}���/�o���SZV|릒{\����d���K��U�����"��g:������h�*������^�t
(c}8���*�6����Y;�@a�,�O��њ��bӒ��d�I�C,���?q�R�8��z�}9���T�c���-6�n��]�=�,��/#�L7*�����&q�N���o.�s��R#��̞hk�!��U���]!���;�k��u��j�n��_ؑ��h�%��>�}���f�����~����B{��J��Q���t�{Ȝ:%_hc}� �OܶV�+��=�P+���P�ڵ�Hl��y�Ul��g�Z�x���i��g#����p{�����9�ɺ��e���JpsR��|�ۯx �~����}$�OPcJ��w���2W����Lַ��R-�.x��"��q�q'�ܷEe�G�3H��0j���H>�7�y�F�tJ��;dj|�\b�a��!�_7W�-��~<�>����~����whU�dۖ�ו�7�Q��͒�Lh��Z��s-�7��%Z<,��5�޾Iy)+D}�ؕ!�[�r��Z�{���_^��Gm9���7N?}U_W�B��*�Z���t��l?{M^k=�-[��A�9�9F_Ik���Z2s�v n�s�~�f�g^���;����7�߰���B�r�%F>��y
a�B0-�r��bư�� �;Q5������<+ACP�d���a�`t'9
���t|	λ�m����w�����4�Ρ�5��=^3^X��z��|�b�m.��v�V]7q3��D]=��]�ݯ:���T��k���n���dw=]�8d��ň׊��mH�,.�:���W>%�U'��qv)s9T�VgCX|�Ͷ3����@��69�xݨZ����]Ɵm��E'9��k�AJ�bjk|>���亻ö&�C�?S!���S��!�6ov=��e�t�<�Q�t����+cO���m�y{���贼�%�)ne)<���	k�-����9��dz��\��WH��S�����M��|��w�f�-C�)�G�{y�x���mA�W�� ��ʂ���¼w��7 ې�p��f��KT=���|�jٳ�ݷ�T��\���E{���o���BTQ�W.��QC=��K1�\��w"z��+%�t�<�A߂����׫gC�qٷ�y�n)����2���uO
���(�� b&��Zc�ފ�L)��:�f֋bRv���ЃbW���{�����*ڱW���_}��b��x�����zQ�S*PR ��H �?j�O�67�y���t�(T����J�͗��}���xx����tc�����0\����5z����D���G2�y��r��� l�{_v�eV�tg��b��מ�DG)z�z�W�ߍ��^����'C���S�i�u��n�mo�>�&�%F�`��w|Q+��%"����Ūki�Kf1���A<��3i�b�S��i've>�TO�>o*}]���V9:�橵�\�S|����O̝��n�K��^����J'�}᧟��B�E�k�=14
�M��,oL-��9�`�[
�,.ۮ��Q�3ۖA��3F��W�MUqj�q��� Mm�Ԫw÷ӭ�A^����P����y�������Cv�Dq�tTL6��;���K�i�5���������-�ݓ�WMC�޿J*�c�0�'s+d�:��Z�O>���ݵa�t2�
��6����vv����w����Y�9����������ck�B��_���Q�M��+2k>kg������k�^a1����[�ە� �z3
��<����Y1�W2�3�k�o�@�x���
��ځjOPcz�����Iw�<��8�9v�>{g���H�v�3�nR����i�Ȑ->q�����j{ļ��s���k�*��#u��m�����܎���C�p�>�� ��j��O���6���E�_M�K"��~�M���(W�P}��Ht��0j�_�<�%��%�iPWt�����1�,0�q�YzЛ�l�u���A���U����%t,���}�j��v��%�:M��k�H�1�#����)O!�rB(Ghut6����FoA���s6/��l'�k�}F�����Y��M���;S.UsZ�*Ֆ�׵v�/<��S?:V������h��{|�k�S�^�c�v����Wz�h���A��B	�����Ȳ���}oT��4�p��`J�m��U�ư��{D�:VuI���y����U��h�m�-�k9��UU}��n�r���W���.-,��<��b�͊���(晵���GX�m.�Jc~ǽG���������K�~[����ӝ�!�.^�LOzw{[ί�ORH��]7�X���w�4N.쪌��|ռ�Lq�縫4��ۋǊ�8K�;ڒo��q������y_�524�3�t�Q����I�R�̵�c1X�a�^Q�Wx���צS�AV�:��w�xyj+d��j��6դR��ǯ������X��[I�]����@逜v�yc���,]���������T(S:����V`�T����x��L9��(WlG� � p���6�ẾUW���>yO5%�=X#r>+�`����h��P�|�������p �r��G]��ٚ����5��u�ܤjz
�QAT�\ë~��w<�3N�t9iRH�辱bs�k�U��=|_���Hu�}�ҵԔ�4ѫ���1��D=�{��):b���S�J�}���u'��hz-��=��iʕ��u{�� n����l{}����ö��\�99��C��|��X|k�T��z��O��Q��c��Gmf����U�=�������r�c�Ya�Rt��5�w+��2���N��]��Y�|j·:����cn�2�ff��I�����v�ޥ9��5k�vn���}��}��{�gG�$V@QiY����M��2˷��<�b�����'Ț���r�^���5f���z�JAK��:���*�uk�Q�t۴��1�>����=�������f.t�7K��T��Ս�*Ye��e�{�Cg�1q4��ԅ���=YCp9�twn���X����W��NՓyS��c_VL�X�r�Z�.O)����~�:�z2JM��S�V�[�j�5<ˏ���MMΛ��Cx#-��z��k�y\7h52/'�*w�^��
�4�m\�if�T\'�Hu���]cU�"�64���K2b�R[m�dx�P�׏���ʸfJxr�$��3J.
�uUҰ�ɶ&��5^���mR�,/U��@HӒI �������I�xsn�jS6�|XMl������#|�>�F��9	G��J��ԫ-2���L�5��C�ų��橽�q���0"S6me�L�ҵ�0#aݝ
��Z��x��)����x�@�,�8�m�WM�*EȈ���`�V�g�.�):�vd΂�6{%e&>hy:Yŝ:�K���.pq5��]�nJ�Z��b7�M��g�gs@�B{�G���{��B����h��2�2��y������c�d�,�����E1��zFlô��¶o�/�_��V��*�ƶ��P�O��n�6ˬj�E�PG���ν�f�Vj���M"�E�<��uw���@V���'�8�+�;�fC�m6�K�i����}X(r}J��jPY1j����V���:�5F�3iA�:��vɔɶ�[#:�J8��-���,�%	cd�P@��ٵ�`	:t7�k�i�m���J@��YQ|w����e>R�m�C�.���Y}�;�r��&)1)�f����*H+�����ܝ���mO� ��&�|��ķ���7��Ӝ1⫬Z�)u �Es����y��v��r�ҿ���*�KM��Q18��*�4�(�ؙ�%ŖŖR�U��v���-�6ܩmL��-R�˔�PӼ�{ +M���� ۽���§:�,�GĜ��/��,���$�;�����nD"�6�򤗆�~7 @$�	4T������S���b�����*���)�Ƥ*!��*�v11TE1EN�`�����kX���AD�'##A���h��8�vuTSD�sH��$����ʚ�"(�h���� �&�Hւ*��*�`�͡��*"��cV54��A�혨 ��+��ۥS�0EZ�1Q�}o��z��+7G��R����9��f�!�#<zu_F/�aV�O�sTF����W��չ�zI�Ww��?(�0mn������G��|���~�Ej���i�Loڲ������&h/��6���脟>�o+۟89�s�K#9$�ފ}g�w����nw�m1��_���[;J��E�s�������n�u9_PyiQ��<Ū�V�",�OTZU#u���&��:�5V�Ŗ��L&+�S�G_V�����z@}�MA��lJ�������}����>�e�f{�����Gvܐ�.B�R�kU�I�</����U�ejmD �j��e�V4�-v�^�{[�l]��NҢj뢍v�ӑE���O	�K�]�7��\�a�mN�j3�[� � "n�G?0��\V��iJ�<޴�Rb;�O|j�`��l��7Y��R��%4gZR�o�'V��A�?.����<�Bچ�-6��.^5��Z�@�/�퓹z#k-7^�AX�d�{�7; {Yۀì{Y�m��S{�s�����M����vP����^�<zxߗ��Ǟ���|s�׾P����~�'l�3�k��U)�Lx�)���O����t��\��AmZ��l�x+6j�rj���х���!1N�;4�ua�J9H�?5�`BF}��x��3�z���5�+�e[�����7�⟱��+�8V[���=KEJNk�q¯�i;�Q7,��u��k����gM���]�#��@twp�%������}��|>9k����w��N��6�������[�Q��_�^��w�XX�3K�q�P��:0Fn)��]�`o���W�,?���͓��=�ڄoG맋B��է���;�R��L�XM����Y��tE�S�cF�N�w%�x�/���.����i+>�s�Z�N�Dk����e��
���V���k{��}�+;�AGF��&�'4a;�̩���}סC�ƅ})	Ԡ-��[g"�]���eI��'K')Y菶&i�t��wP��۷�:�]���/DC�5�ҡ(�s��}��ᮤ̗*�P1��h��U}_R�(�&�6qo���͆ru㣝g M>E��8�<�o��")�лJ�g�b!V��=\���B�Pv����J�������T�����c�$�r�V#-k�=��D��nfZ��C�%�KJ��>��	�=^�3N��<ʵSs������W����@W���0�
�o {��PgP�5�[
���d�=���c�~?*��ua��|��!G'1,��-�,��_\�Deӥ��.g7v��C�f(�����m�BŐwo".���Z�1�h���Č���=*1�9��9���Ȑ�w�e.79�e��=��U�բ�m�,7���Z[J�T\��^_rt�l��M4'r��G[�t��r����o
�����^.m���{6�B�c_A	�1�� -����zG�^'�n�����Zp���;B��ٽ�,�y���7)��1�(����}}�����=�E�xV�ޓղ�e$<�C&��!��^;�2��A$/�����ȟ-GV&�B�8=�3��={��H^��1�~ͮW]�MV�D:[���e���B㦣��ׂI�Y�/P�PA��i������ui]pUz-����ݳ�x����k�""�P�ZT}��<�}J�
T7Q�x�\iߡ��F�#�����55j��t�0�F�u���Lp��mi��嵵�������u�U�Z��y�r��+r k|�s�p-�Sy��z�p{f�����~U���)�5�O�������mvHkV͕��O�A� Fcذu�Qې��-� .����lvk��}t(��U�[Zj���_��Q�\�/�_my�B-���]}ǥdT��2��q/3��e@Z�r��W�L��]����	��ө�
#R� _ׅ�?'�Ͻ��(�*�xtѶ��h{�XSʵ�s������G]�'K"�Tm�\0_��9�q��H����S�Ni-�R�C�|Y9I�)8�6���GU%�Qa��.���3_}�b����$@Ѥ��"��f-������\v]뮰^�XP��*���;�=��}�Ff3���WW��<.��לi)�kE�/�_��3��)�TǏ/�m����]� r��>]ޜ9f�n!8�7jQ)k�J���:CJ�l�uu}-�\�±(��&��0{�XJ3`	�U�l���,j�q��cڭ��	����r��"i��ɸ����;�O' br���s�G{�t���8��ET�b~��]�e]<�x��������}�W����c�
ƺ[�"	��y*������p�c���Z3bx��[����:�9����T}u���HM���X��TU��d��h}&�͋�"�����k(v��ȚT�}U�TrA�� m)��!�W`B�3e*W9��7�[�1���՗�Q�O��"�jt�'K��-�
����[�(��G*�F����QWyI�t��a-ʔa�:�)g;��`b�;W6q��[�Q�1�x2UԮ�W?'���\���{�+���%Щ���<�<)��t��cj�eA���aO��e���a\�Ǟ36��=\����◜��J�LNl�p����=P�EN^��cw��|�TD�i��S�LU���W��f�+{<Չ�
���ɐ�-���>��N�Jf`a�;��v��si�˰���VxR3S�<{]��Yx��ߢݜ8���WH.�}�}Z�)�{�����m�̹�Yz�8�~��6��秲��tf��G9�sC(ڢ��#7�TS���tr�����$R(��,X�R{5u�#�/����sBFw}ϟt�Z+���4���7�<-&ƾ�������1b�7*�i��O�y����%����p�;[|h����_(n�ޜ)���n��s�s�LVd�KV��̊ʗ3u�S\>��j�^��Rć�7/�[�ڛ�sR��щ�����>�f�A��>�(��=-�j�<�i�Ҭ�:叵�c1�&$b5����]#��*2��wM��o(u���p���.���U$�!�\�'�or١�t��[�~��ꨣ)�{'A���^7�&Q1�zKsq�Ʃe��y�m��g��ϻc~i'���|�;�Ff��9�j���=����c��L�y��hA[�WT�}�R��A�}�q[�ô�߭*fe�*콝,�F뼽�o��=OZi�??a��֫�R��I{"��b�>J�l�R*E��]~����u쁬i�ޘC����2OH�v{o��E���ҡ�>�iz�f,�����~�ILFW�P�GM.���j� ���:�U���:, QD�ٜ/
󁅜���ݬQYI>�g�z��ӈ�[1�3��K.�b��2����,�.9EJ��b��ݘls�����ӑ�f�G��R�� ͲkU�7��<�%���w�G!�.���y%�թ�ͺ����+����H��=r�w-�#�͹gY��UԒ|�=�r�iǑ���u�պ)U΢];��I�L:�Z����l��f������"Ύٜj[��/IR���� )�jݼ���+�M(���a_
�W�u��Ak�Ʃ��{D R���7�����ب�m=ז��y@�d�:jn_$(�b�{�W�|I�~eU��b����h�n�iR��Z3J�On���<�AXhj�Vt�!#3M¶��t&tWvр�%H+��A��;�ӧ��*N����gDR8��o#��(p���UI���)V�E[�$�]w�g
\<-�wR�jZS��̩��7BT(s6+�i񙫻t��BJv9|kr�<�n[�t#'�Q�j�3_+6ֶ��M��MK��ᵷ�^�˛�Mn���c+�K����D�ހ���B��D7��Q\Õ�� �̫9�J������Ѥ剦�5(�(��;m&"�o��*\�ղ��,�����1��`.������C؝]�YtJRF�{��hb2�0�_qC��Z��Dp��;|�]ܱ���6򸅫l���
��t`���ӛ)h�1���j��Xg�ƚY�J�zi%\0&�V.�h���2we��w�Hf���5(p�}�O��e�e,��k��r;/�D��e�7�l�""8�K�s�n^K����n�Y{k��/cu6��oq�ZJ!g1j��FΧ�&i@��ږ�hu5�2��Tœ};s2����\>�;H$~�$h1��ADP�D4\�EDI�SDD�kTR9�TLEW���;f��J��G6��jccQ	AE���(�e�"�8��+���h�

֝kl���ևN�1m��x<���)�(b�;�ld��**(j!��h�J*!�()���N���(Ӧ����I���(J+Zv䎼�ƑZ�-���s5����LV�>r��Ny��]װւ4�/���3U����V�;�x�)j�� ꝨX�T�e�����Oe--�Dj\6��/1v�{ɧ��Cڒ�yQ�Z�S�]�bbJ�d���}�`�U��N�n:ݘ�R�I��
yW����g��!��:���]�$R�o[Pem@����?�)�Ǐ�ibiYtNj�`���U��w�C3T�����x���I�LG=<T3R�4��������gP�3��7�q�{�z�iM��e���;[+y��"o�Tó�1�/���%�YY=��^�K��7��Z����{�&Fj�0h��47*钽8�1�۾���<1na��Tzun)0���	0c���u٪�bU|��C	2p�����	��ʍ����Aܑ]�6Q z	��W؎��:�˪��r��soG@�F#8�ZƊ�C�ìch1p�ᐫ�%����^�c��j^�ذ:Ԍ�Y��!�z%�js��@��-����!�Wb��{s�jGL�uC����֕�7��M���+�O#��yY�ע×m+�&�z�H�Ƕj@:ԝ������U��7��򘇀ϗ�b�4.i�(��mz"珔��꾎�M����Ԩ��ŋ�۩��!��I��Q���ټ�:�Y7������[�,�wҺ�0b\3Y��p������sA�%u�̛�cn$�w=���X�W�TLE�=�?�{�N`�@c�g�:�T90���*�=3����oy��|Ac͘�A������4�����]���Xa��z-+9>�}�<�ت,L�庚fX����W��T�J�oFG��[�y�wF7jK�H���#�8��Nm����kd�5�ѽلr��9��mվ��-�����BJ��9\b�1�s��6�7=:��WtZ�7���B�����n�3?jW�<�ƺ�l�\���m�Q��\�Qa\1X�����=�j�~����Z���i��D���f�"�h��G��m����W@�5�6
�uLU�A<U�����l"F���2�Mv��:�1�*�݈�������U��Rc���}��З[F����G�\����ߔ��-o�ۮ
:����|�@=jOj�*�G+�o���1Kk��2mn�DY�m�����u̐J�Nꗂ�����N<�[ggw�f�?x�v���'j�txׇ1�w����:%D*�i���ύ�����t��sLm^�7>k4�wګ*����6�w>��[��#�JT�I�%33�5j�!t��wz�]O�zGl��֒6D�"���o�\��W���0 |��R��V�����xX��W��j�eh���N��z���="�'4*���2gI�ZE�Ι{ ���}w�X��6)�-��t�7&�׾|����l��ض;'Z�+�|���R����-��Y>�K�O�����Jd�yX}%/f�n�����F?���Vz�ѱxhVl�Y�-�P�9��-�+e���t��Ĵ�{�w�P,t�i�Zw�X�-k����͜�*k�,rP��U[{�/s�L���jh>R�{㮓t�x3<�+��q>g;����|c��bt�-��y�=$�߉��������Ψ���4��i�\������3�{�_<�z�N�~�)�q���ɻ�gKh�g�m cS�pW&�R޾[���+C��Jp���i�j�s'[ݯ�)��a�
d�T�وVAM����Z�t�����a5�\�s�?��Wפ��~d��ɞ�Lr=j�O���m��87�*צt�����9�(yFv�w�&�W+f��J>͏�UV�[�R$Bu��E&XS1���[�W�vf���\�OL@��
�IyeG�h�[0�x���ז�ꌟ��W�Ѫ��!��M0��o����g=(ɒR��A̕3(��4�;+����UBc��d�فֳ����1����H�ä���j(���hd�fN���\ǣ�(f���Y~�Q��6�5�-g f[��
�Z���Ϋ�)�7^<h�n�9��9�b�Z�+̒fG�0�9���j	���{�m�3g9h�%$.Ț��5U�� ��g����>�bf}�7���ЕX��K���<��Ӷ��m����&��v-G&K�L!��3!3�6h]�s��m2��i:�j�1+}2�/���V�}�<��>r�o���}T�xv�Nf�\�|�d�	���R�[6k��������������>��?<�(���
�Zv���v�z�:��;� �sGho���|&[�;�Jml�~����2*���_�̱�i�2#u��=�'��OYϮ��{��m����AQ�Z���Ƽ�����<Ӕ�Y�g�t�N�W]�m;����xPu6l�no)���JN���Ys��BK�f	ם�5�N���V���b/�Y�J|�4���r�+۾9�U��ѷ��fK}T��]%)�+ޜ�l�G���ʔ��Fz���鿸J[�g"^�V�4�R�vG\y;+6�	ޕԹ�ٜy�nq�f̼���W2R�(ý��B�b�L/?/Vxhn�ar:�����Qx��;��V�Oy�c�k4%Ce	����a��t7�aQ�����L��H©5�ע`����nOF�Pi<}9k-wwm�L7k����T��c���:5��&�U������YSn}����$����z��n�]��,�p}�	�2�1�u����f�;`��R�+l���3r�n��q���[��r�|���32Qo�(z�|��F�#�ݵ��V����9���ī~�;^G�s�;6�K:�V�0�H�Ѻ+\��.f�v����D�zg{7����ro��P�ʸ|{�ql�N�;|�\�O4��!�
�#|�m=�9��U���\Z�/c���
�b�z6ōp(���s�E65�[=rl��Zu\�ba���
����-[CVl<����o�!X:L�=�*d̥#�3��~��8�5��|���YD�"�.�k/��,�d|��he�xpm�ImY:L߭S)�t�{ܖ^�:�]H��0<��9QQvM���t�����꯽�����;ݩ��5�W�)�4pv�9�S�渮�|55�!�5��K��f���6!t�i��y���}Y�p��ʡ�5�������՛��W:=^��>₶���=*�kl���l�����I�֩��*��w�g2����H�0���yY�OZ�خ�ȓf���k93���q< Nl��?%��oj[ѕH�:�&�����&Jr���+c:���8}UYi&f<m��Wq��W[�;#����[�*g��ZGV-�Α{G���͟{z��F\\��vi�b��7���c)�6v�M��9�h�d�̳*1���rI��ˬ��j�9��qL�.�urnF�����g4t�8Όh������#�!{��B�'MY���阐}�fq�,�ۣ���a���x���5��GJp
Q�f�����ȫ�������n��1[��4���-���U;i��T�/�9�7M�g�R��-�Ճ�`��r�=���xT��tpn؍Nč7�c��.�H��^��(�
R�֔�K���%P�ف�7�2���_s�mɍ���e`I^������R���2��݆5�,����R���Y��s����aA�����G�,�Gy>\R�;��1��n;n'X��}W91�Kf�[RQ`�өs�#F�Ȩ��+�1�W�I��$��e���D��g�l�A���F��A��,�kŤ������o(�V+b�ѕ�\B��'P�|u5x�`V����0˱�cj���ܟ�2��/��ݼ(RY*�����}���R=M��,�g-셕/&(��ms�Y]V;Eud:��a�@�v�l����t?-�9Uӗ:���͈�Xޙn�
��b�Y5|s�!��:�f��Kж���Q��������;5U��L��@�ڔ��Z��s8��(�����\��m�R��N�5u��9:��2%�{s��k��B�w��Zu$sz��E�N7�ZR�d/��S��ص=g���^(�AJ��Ǚ�41t��!Ⱥ֨�wh��l 8��	AIwF^�h�SP+�U���V�.�v�tKU^f�v̨Cs��t�R�"]�|�4���U�~v!����	�����u�#N�bB�
!4�ш
���"n�)�(��
���("()�C�(ih�QMG#�y��fh�&�
�w���%4�RU1=�3PSMP�b�k�i�RD��CT���&�qd�\�CA:]-ZѠuACCEC���R��`�ɭ!�)�(���5MMrE`�G� ���#β_y�E#{'U,�[�7b����u����؁��]
.v�t8���j]��7ϿR�N��:P�����*re���(�aE�kUB؇�pT�CKa�rƔ0ߪvr�����-����BN:�N�t�.�n+����"jo�٫6�\�.��E�Ǘ/z�8nV9��ݮ&�
��>��;EE}w�]�|Xx���2�1:���`n�s�sg;o�S�UF����7�{����O�{sV^j4`�x��5��X}�>�o��ſi�9�B|��mo�AŔ��:��Ϻ�-��,��^5��%{�c>�kʳ��TY�_V�Xq�)=��w�.�?A��Ѽ�zX�q���И��em�93O�LX�Φ[��u��*�O��6���ߙ��A>G(�	�p�v��z��3-��¥vW��6��l�p9c�'ӷԒwu�|!�zQ3��8�IJy�~�z��LR��h;F�uo@��Մsd�.7�e?g�����r��om��{Ag�A��R���y1�3ޭ"xx��^�3�N�/+�h|�I+z�����ʒ�N�=A>��ST���s�v��e5o�U�w7_�q�!������P�*7;D��	�lI(��T4�NOq]�V�4|�;|k�O��ں��^"\�v��/L�@za��Ï�k�_���B�J��C3�tV�'3s钵��Vb%�����$��?C��\]?,��Jf��-���O���'�kZ2�Č*��ŧ�]<���F�|}ކ��g��j������%���0s�V	�5|g�^�!<�]�D\��Үz�y������=��o��}Κ�>���^���n�-�9}C�"�����#��2�>��s>0mr�]��Rkm*ú:]w(c����g��sP���r{��;ސׇjT��o�Α��xg��^r}u$
%��/�3�a�r�l��u�v�Cg��Ws��M:�f�Gd��U��d\G�������j�1�+^�{l��w�X�.��A��v�=�ļ��.�d�>q-�U������-�X��ź2Q�U	��&�Lw�Z��Yw���0:�_��8�c*Ca��RT-]�9f#����M7�S�-oC�HΥ�	��-����@�v���s��K��cx\��q��k�ݜx�ms�.�^�usnẹ\j}Ȟ�~y5��~�6�A�)�|{�5���"�=Ɂ�AՏ8���o,��Gޖ׽���LQ\�Y��nc��R��Nh7�it�9y�!���к�۸�^�ɗ:�+S!\�o\%H:5���E�V����l��-�cʉ̀��,	��;��-�W�j��zV��dt�������$�W�5:q��zV~��<��~��C]ei�a���M���<t�^{�L�gL�V� /8�ڲ兆ūA��?p�/=� ��G�>zt]��F㖭�`ѵ���+d�-��ױ� �M�����Z;Lv��^�ĺR/�:rzN�Z�spϵl٘�i-E��Ӹ��Y�Wu�:F����=7Z���T�#|�%d!n�'��t���p�1����X/؊&���Ǽ�����x�f��X$�4���ח�%�\���+j�OVґ�ʾ�!ڭt�d���(�0�P+a�	�-��u��n]��^�{2�{u-�d��Z7K��\k�'�U��yoS�D�{lFl���[�9�v4�wAظ���}�Hm���+��)h���L߸���!�=�j>�J�z��1�����=LBeN�!S�c�g����Ts���W�S���Y ��ڭ>���Db���<]��<�ղ2'+���J����}�Z�/l&:�i�Ի���5Ö�p����a��h�cuS�9:ґ�*��Y��J6��>��$��R�s�OS���::u�@�t�1�Q��e�z�&}&h�8��*�RA����A�/�\�T!vZ�(36e[Ѧ���P��T��#�J�[ΤoL��� ��w�rb��{5]��L��2�둑��p^�$zI��ݶ���r�`%�����O����H�:�������x4l�u+̗�'3��"� ��E&5*狭�(�ƫ�_��;��JPP��d�;�{I{��6�g��[JԸngk��4u�z�*[蝩�uOܶV����q^��w'�o�HYԆV���x�J�W�w�^��x1�Nu�����T�m�ln]�7=�w����nT7�cy����H���z����U�3Y��n��膭�-����bAo���<�_X���s�Q�'�̿C;x��o\�����gEeg<�e��CM=ΟLC	�`&���8Q@���y����ϕlٱ�i� E�Q^<�4v�-@��4\�E��mv�v��X%}w4���isnC����Fv���6?A(DC�o�������x�{�����?y�Y���đ-�v�瞹�r����kΒ�+����N�!�%&R���2���Zw�oy�'c1�h_�Aʛ8�Ԭ�׳v�����Ą&�sRA���L������D-9%ך�e6�-A�w٫��gT�Q5�J��a�
n8b*#{�^yTg���R>�/h}��-���ש(���T!��׳x�[5τ��ƘQ�P!�Ӥbؒ�P��v��M�vPPwKL�3 ���b'zOV
%�;X�I`��e¢�)�H�R��JU�_�2��`����{�� S�Y\uv
�UNݬ�����S�1���U��E[��<��-��Mr�k�V�̧�?tÛ�Qf݂G�L��د�Oz�]pC��O�n3	�a^�m��Q��/	�3Uic��B�T�^k���2��B�[V)]�c�{��F�=�gb�W�<��I�缬��h���{�;FY��n>�ct�fU]{(�/~ϧ���;M	a�N9J,��;���wԝ�l��6����hؾ��T!�N�3��DݰtN�=�= �ի��0Õ�o�z>Dg��C��HK�h̫�o����z-�@̜nv Up��J9��=ؒ�����֪�74 A�}dѾƀ\��|��c����l����j���Sժ~�
[a�f�ʷ�7/�ċQ��m
P3n$WGɦ�N8��k��avU��	�C+%��<R�X�Ք�����i��h_l�S?]�"_X���:����7U���+V������t(��=v�>R\轨��*=������=(ͷ�y��|�����
Ӂ��i�[`>��9<ǟ��Lu����B�-p��X�d;��x�v�{��#�r��x���"bO\����(�}�x&�6k׸�ZU7ׂ���m�M����T�r��}ա"��$8�� Ν&��i
*���#|/���v�7��&��&$��o �[�v�[;Q�/5�@*1)Wn%�<j�V����N����ߵ-��tȲ��>�l�3}ؘ�sU�٢�e�l���f9�rei��?9)
�:��+u�Y�5a�\��h�v�{��[|�;�H�;���lҲ�j�����3s�v2�X3���-2�㽅��۩gz��m��\2��dr�ݲ��z��(K/쮜j��pG}+4�����r�;@Qh2Ü3Hvsg/���L�}�(SnT��VS6���e)��Ŋ9;i�̕��hU��Aԩil�(;�.�\��`2�	���q}���n�P�]ܒ�԰\�c!�m��@M��7K�j��A��(t����riW�Tˆ�YS��&��6�{X��UY���y��ui1�0)�5�0�T�ӡu��n���(HQdIy���ŷx]+�,b�A��+��N�r˸T
�zzѱEM/�cU�!j��E�f�_��дR<󶒽�� �B�mK�
�[Ԭ�1^��R'(�=������5�kt��b�a�Ń�s�čK�\
u��x�c�h�K�#y�ې�u(w�Ů��E�m�m^DhRZo��cX�<���(��&���i��^�i9�`׊I�R.iF�� ŶY�mO��ҚػIӺ�����L����*t��{KK���C/B7P�]}xZ�=�%^��ܗ�����Y;b,�xЈ�4Bã���Z�vr��U�I��څ�x)������tm���/�Wu#��c�Y�)$B�r��k�,�&�s�h�juuJ�\�wl���x\�f��*,e���{��)��t�m ;D k�ɓ�2��wf$�l�ֹ����ʽ�����U @|�D�CJ[4��P�QF�64Rk\٥��$)��i*�G�r�R��Onsc��!���!4��@b[���QKJѠMCT���P�f�H�+�:Zi
�qi�r��ZtP���������v{,G*�D�ȤM=�lrH�byd��sr(���y���E'9�C�9���
P�Z|Q<��p]�]�j�"|7����z�Wd�Ob�+jCQ�u wGvL���U�t�5�C�׽V�Ml���0�:��˦<�r{\��f�N
����j���n{��T����w����5�+
��?YFb���I]IpX�.S��4���ŏ�u�~�� ��۶3�el�D�ӕoo�j������|S�)N���9��n!��r����K�2o�nQu&�.�7���(�xwӧ��|+eb�J_�[�tl+��#%�݁���y��x��s��7�5�ޮՉ�勆Aޮ��w�)�9ө(�YoH���3aX�w>��8�;ݫqa��L|
3
����)V�2*��)+<j:��c�1�zV*Q��=p]	��+��'E�[ˇ���(ӋQ�C���`yո�L�P���:��u�p����K����v�^����$��;_a[�ƵVg����2O{���&3��ﳞ�qn��V��S��<2���u�VZ�s��cF��A"!���IW�s��'yl�k�Z��*���}]:1dT����c�+��{ֻ�Rt9�j����}3��N�|�n.�k!����Bt����٬�3-��
�nX�X��P��,�5A���9f0�Gk�7R�CV�]8"�G?<������9	�]��o`]��Gϕ��I�'9�ڙ��G�T�t*���^��I�$�7�\ᠨ�5��x��W5­Υ��b��n��+`�hME�D��ih"������g !��x|	���|�S�p�� ����"��R���E�ڱ�)愷�/l=Uo	A��]:�wC��Y�f��Il�m�jo�4���h�|����Lg��͡F2ʥ�y�پ�?!e��Ǣ��Ns>C���+B뱯9�~�I{Y+4�+l?A=��a��`�k��׊Zv̋Q�D�9Ջ�ܺ4lt��f�wɭ2oͽ��=̦�w�����Y^xW��zL�ѫw����j�fz�HU��-��V�t3�|��:^qfy5��D0ܮ�ǹ��t2���{�"�2�Ce�u��e����0X��}��(Ӕ?j��?r�2�rS�)#@�(ȫ䵡OD�!@J��5�6b�]/LXRJ���K�=�;�'?��&����u�EXt�;^�W��)�G�YZ�BfDX�W���t��3�Av���W�C�.dào���D�J������Ϣ}���M�-�GW�����ڎVKtG�i7<�c��]�m�X��ߩ�r���vj���������2�2�R1MK�����͟j<���+�� K�E�>[�'b���G}[�#�d��\��;� q��'���Kշ�	��9f��1��ӑ�YOoP�k|]���u���y�4�u�gX��{�~���>nn<3L�?q�u[��̖^�^���^����%��z��:t~���Y��;Γ~�ʿz�{Z�H18'�O��:��Y�^�i���vʧ�7ڽ��=Kp�Uu*�-{VKW<s��}^�r;�yM��[����%^VS:L!�KsS'��qN��W��\ևu�4ú�Ou)k.�}�Ӫ��sµӐ�XYzj ����y]�]xJ�f�z����V��_�B�nc�ƻ�7k0���9�n��:�(��7ޥ�*�6�4�Q��Y����=�~@S�L�Y|r�:��m����c�e����<D�*>�A�<�_.��lM�vy�H�1�m�4pB��M��9iʱ��i���W���u�ð�e���l9
zj��%>S;�;���?������KzP�R^�>�Y��p�9�Y��q�{�A���l�J.}v�'w�����z}+DY���^��^��a�/Oxf"��~`j��q=�+p{��MW�ڙ;^�?:��e��д�L���҈Z���K��!b�M�$�Y����Gp�5��[�Y����}5[�ޥ���������-Jf��*���"|"�/�y�z�����)<����mfR�~����0����1ypA�f*.���y���|��QT�15\7�i]�?B#W%��zi�����\��Z�̢y�+wPi�\6��p��������5W�T��>Hn�^e��"�9�f,�l��*�Vg���}'Z�/���'��桨Oz(��_�nW�+�rN׽BEG���	�⟕e%���ĳ����(H����ːϜ���r��s���1o#pn���>0eE���.��Dk.�zO��ImE�aN0�]��F��& y�U��$`ޜ3_\�}>�yLϢ �W1	<����uDR�,#N��٩���ĝܣ3k��^Lx\[�JAQ?z3W��j� �J�K<������M�>d��8|�$O��8dRn�d٢�g�5o�.��n���>��)懎��:�^7�N�<;5������ҽ�W�&�R馘Ý�,�sG���e���[��Nm�\��5ːp����N},aut�)2Zy8�m��P�uol���b��|>��]���<ʈ��#�dθ���lA��=~���;�u������^��/�O�hc�NRPNw�,�F����8�ΔkЍ�u��|�6��ϸ�Q�E�H���hp3]$�F�+끾�8
�4��N9{U�Ж=],�zE�q�uK4W)'IQ�bL�]@ӟcgu�0��J�������~Ȳ��9�!���p�)F��])����]7����t��3P;�P��<�l(N)e�7�|^��ˁ�ޗ������;:|,����D�4�����5��g��}L���5T��|����H���3@��$�?c�j!�6�5��J�/�[�]�W�A��:Ge���R�,���F�5���ͼ���~���'w�$x�9&\qu�#��g��t8���[ҫ��a�:�u}���=��2�rz����e�2��o��G��yA��t�^�|�[��ǎ���j¼s'#��f�7+'=�	����?���p3��]�ﲥ
3���:ʐ�ҲQ�lY�5�}�׋}�_�#��<k#�r�{L2J%� �Ι���S�k��{x�|S���F�*��l2e:�\u��Tz/��Z����ܱ���� WQ`�O���q?H�� *���X��G�԰d;\��zY�^¸qz.a�g���"�9ʉ{�W"Y�?7�y�{�p���N�Q��`"d
�XV2%27�٦��=�0��ꮜ����z?<6�l��FMV��l�	���f����^�(��z_H�;�f�nE8�#rQ�Ǻ�;��9q������`7,������O��F1\���9A:��{BN6U�^r��xD~�$��[� �a>��pW����b�OH�~��W�n#X��C�9����w��:[��<�s-�4��r�t��Cye2t��JOy.WenN{�_S��yI*��|�jK�	���h;1�~����S�lD.�(�E��NT�5�^+7�R>�:`c����BD�㠊�w(W��X!Ts��q�u�H4}�Q'O�c���:O�������G"lدm{����ql@�����L�>}Ш��aG	P2Ρ�'7�<���5�*�\E�x��!O�3E{�|T@a�߃��ͭ؂y�wms7#QFM9��n���>	S�n-ć�F����u<���"�?��E���u������r�F|_����5�_��q��8����}�����쀩̜PM�������IUa-v4�d�p�g�c���b�-�W	w�y�h~�l_��٨�gox=+��8�yH��n,��l��D�	�Z1Ӓgp��
�Z"r��SP� �mv�t�Qj7#�3y1X�/A�I��-��x/���:oZ����3�GL�ϹcǹERW64��r�̧M1��Kn-�\bԝ}]Ν��1��j닣C�eu��� ��f浝�e�d�3lb.�����v�h���8j��ֻ��*�N��s�	�ʭ�fﬄ	��
�h���ei[��Z�E-}r�'7q\��H���A�4T�����s+�K��QN�+x���r^����^/��WtB�v�CI���nޚa��$�����g)��(���Y�ph5
e�����e��G�����/��>��U*�W_T�x��q�R��s��v��o	�>R�#0$:�{Z�}/ �"f̬�\F3ٓ1�A��t-���N���-�3�����z��/頨[Y�x��z�I�2�˧zq5���@������In�/�m7aCKz�L@�{Æn�es޶k����-��8�C`�.PCێ��2u֥t��\Q1>#a.MiM�)�B��u)E�w�x��D�=�^M�m���@�핣	ꋺ�1LP�Yw��7�ٔm�B�:�i����N� �R�8`��]�vl�x�v��	\Rک^m�6V��c��~eq�,��}��MTU��>�+7PѲBɏ�'7�keq)�/( �q�m�(챒�mazJx��f��\��֥{�8�a��Q�*�()�enS{wLHn�Z~�teZ�('W+]ʻ-�u���:������X'Rϡ�AH�����p��c�:��)�²�}�!{�U��Lf��m>��'�J"c}�����P�C�[� �AHr4�4P�Ԇ�{�C�t��]'cJ�w��N�I�]ɤJ
ѪOR��
@촫�\xԁE:���:���(�� ��9���c�R�4��GT��%;���RPhtO0��x��i��NG �Gg��P�"
K«��IT��w�y.�ҍ��Ψj�����[d{O��*�N����I�U�2�:�;a�v��KV9�}Ӹd�g2sM���vp�.�m��2DQ�������w2����^&j[�<Qۙ�x���GQGi'������.Kq��ɑ$�L�/��u¸�����r�Y�%�zk��C~�������'(G�HR�?:�~>��WGl#�dY��+33=�V(��,���Bi�}�1�I���B#�"�o��\U����Z��ӔMF�e�3�l�c&*5�^���i^1��+���ܤk��'$�{�$Ty��b�yă~
�mfx�;�bcLyH�0*G	#%�s��A<���e���>���l�u>0d(�sŨ$k.G��^���\�i�����i�|vA2�B��;�4B���zp�}r���3��̴���-�RW3��̛Ĥfޕ�u�[�.˭��/2!0���7��M�;`𠹞D;�f�.�X9M�d�[� � �@��:�r� �UN*%{�#��#�;l#[��V�ӵ�w�Ru�+}��E�J�c��������?g7L���&�N�P�휉��?t�y;:Y5�g��$�E8��n(s�	H�T�f�,��K�y���6m�;�#z��7�A��e5��7�و��U��n�s[ȁ�v eFl3q��#���d�e����)e�Oίo�1��W�?\隅�3��o�Qފ�רq��V6��ڛ�b���^S*�i6���0l�[48�&N�(���d�}�܄1ٲ={<o�(g�(�����L��E���>���5�~���y�pG�$H�"��_E�:�]����$�z�tֻ�yG��'�����'j�_�/����K�_��OP�YC�ק���F�Sn���(� 6vٚ)�v�o������@`�j����[�P�o8&[��lt�>�v�)	X`E;��<*F�0zkD-���� �^T'��$���a��Ɂ]���k�"ijy���1D�|u�#�d� N�
�J7fz7�Q��z������|&8�s���M��6�k��)Ŕhק����T<�����yu>��K�G<l(���j�U]�fi�����9!L3��c��eD�J�T1�F����Μӗ������>͚4��:��i�IҜK��Pz��[�I�4�]�O@��=P��C�N�J��N�g�������e-�l'���ba�3K������O��2�����N�x����C��M=o��},���H�N?�ᖖ~8*Y"�~�������|/���H�)�j0lq�~W[�"n_�@����W�tӫ�T�}h�c3$�#���G%e�`���u�u��n���R�Ƞ,*W]�u{N^l7&���5��x(`e&-���珎tqҎ�
�p�"�̞&E��=��[�:ǜv�\I�M���,�'���Gܔh���>���㪑�N�����hzB2*4�s\�/�2o�F��u޻���}���ɘ��
O���#���j*�4�`���r����-?n�:�0
?~���xY3K�1��'|9�y6���R=�~���B�{�㠈ۑ��i
)��«�!��S��Dx�R�;�H��4�d���~ܩ/{=���n7��̖��p���P�P��&=�nB���f��9"�LK�0l�󁞏O�xz  �$��'֯{�Ft1��n�Ȝ�Fn�W�3}>�N����{1$�'�
�ߍ��ܸH�a���-�<�~��d���/Ʋ5ޮ�PAi�eš&49�T�\ƹa<��oB�we��;��N�M��`��R�ӵb����6���a�>��L�����C򬽿I��=U������+OB��|��A7�*4wg�e����PN�f��K"R���H��:VzFU��sVW�{u(|��z4kfE��B�<Q��{��8D�t���*7��OWn�z|/�^������8���?�a�P�[j��u��B��]�������M�S�*�O��Z��88_����C"@՚����g��|����2f.I�2.cI3��t�C!oH�[�R57�����"�r�ƵȐ$��2�B��u��s53��P+����cA�>��P���5:�Pw�H}����w�>ٙI����ށ�U��9Ŗ�2��,��q��$��c$�X�u���*�sU*��-�ì�d�4����.&�S�R¹V{��.<����ܷԁ�u���m��`�6	Vi>��rݾ7�}ש%�K=`ƚ$��G-@ɜHu����5�����~e��䘽�Dx��M�aЍa�3�NJ#��,T��{��s�����v�C�T�G���qj	1�C�|���^���>�P'�!\l@s�Du[��S5è�C������Կhd�: ���r��ts����xޚ4�`�b#�f�{����8I�r4���T%��(��qҏP%K7ۓ����x[�����('��ހ�8�F����>Z&#˽�Ωh�DY�9�E�H����*a�p(�����{j�L{�O�d	��鐮<Q���Y���̜(��N�3mP�~ş������슭��L����L�j}q�EL���Pҧ����;��et��T!w�ELE�BJWc.i�!m��	���9�����'@ڏ"���@�\3#����K�x�7z�E��%-n�&��fo�g�ӧ�,��H���q#Au�L�o�����Ь��y�On0���7�'�ƹH�>�.�Q���N��0+��j��f,t���b�b�,��f����I펕BnL�a�^�}v �#�Ҳڹ^�X�e3�F	��P���$�׆�C��["�R|Q��4�G��Mt��|��ĸQ0�[���c2áq(�El=�H�ܡ_{�M�����eK�����eN͖O�?/9�*�O����prV�9!�ʌ���vp�9�7�I=����Q�O�Q�6�uI�O��E{s{yVxq�2=��UO��!��")H�QV a���-����\��sf��3����׬z�%�h������,��'q�Y��`1C���'V��9��KJcv�.���G8�.�k? ��XT&t/}5	����Mf��a0�@=�õ^��[���Eb�i*����ݯ��(����8Gm3uj#i%O_�xo����
$��FDq��#9gT~ݡ�I���p[u緡�&�4�9�'�i��r�0�D_����p�ڧ��dOd��,��Tg�x�*�PVO�muul�>����#�� Z�h8ΊQ��$J�B4�@���i������kP�yБP�,��ϛ�՝B�2{ю8�ۄtntC�����
>�$�L��D��9��g\�|�P�{����7�ػԆ�0q5�
��5�*����a>ܬ�=_�f��^ٌ,��쯿r���A��Ѝ�v�\q[���s�k��C��#���@}�[��}r�P/`�|kD��5B[�*�����VEi��"�A��ޭ
!��V����1�S̠wj:�����H�����mX��v�%X�U��R$���(�r�[�v��X/@����{��R�grQ���,���P�^�M@��Z��0�Nu�C%�A�G�dQ� v9�����$��U��J�_o;��L!�R6���GTx�.���'Ƃ�ӹ��y�[>�!�`��}lTY����S���lt��w�+{'<����7ǣ�t������hq��7�gՒ���О3v����]#� ��_E+c���nGZ�6��4O��������Ng�_@NI��^�ز���J��5C$_D)��qڭi��x,lȺ�CK+:E�W��(Æ�u�H��{K* ?~VD8qE�7�J,�@�Ў\
�^l����؂qǌ�aQM���Ʈd?@ܹ�Ƽ�ɓz�Q��#!diYz��û�K��y����{�����*��vm��U�{ʜCv׽����짩�7�Ҁ�׍\a�������[�&'
�74~�?xTc�I�7pY�`�1���o��4��,���
tux�{w}^}L�@�9q@һ��F��̐yȰ��f��lt��^.e>���8|p�ҏy�m:��� 5�'ٔ��d����D�}�+끦B������C43?)�q`��Y��Ms~Y�Dxf��KV�� @	��9jL�C����U�{x��o���U�'�<�DG��&�����i�uǅg���z�p��o7��_w{�,�${`a��vX�5(�f�-A!U�Gc�jf̱�#àzAr	���[��$w[��f�^W�u�$��/UK�E��+�I�����9��]�+�a�p�"�x�.�
� �D���qҏ�,"�^��4ϩOl	�k�d�jqkO\N5[G2�ա��̢�h]q�0w
����ȲWe��6�H:�+��+nv���"�	gt!�4i١<�*C�5ֺ�q�:\���=�Y�y�`+��X6���hV�/���`"�����!9����c��G\��x�7��uܚ�.0e���9��1s��ӓBh��b�B���6[��ao^RV|�nu`$o;5�L��ɚ�9c
I�(��F�#�8���V������n���V7)��m�F�;]ғ�I�e�����ww*ipu�5N�͓'m{�wM�[,���r1�A՘E��3+n:���Z.�T���9J�Z����q�am鱡FX$[Dֽ=��t'�(�!��d�dW�c/�#�9!���E����syLm�8ڬy.�얃���pXn��[oqp@�\�O�Z�� 6�Sv�����Sxr�W�k���p2iy��)a>s�6�S��x��>\ya�^QK��{��P\��Df.n+�YO��,.ӴŃ�,��5��d8����u})�81%��E*�3���gIƘ�Kd0-D��^�d5�f7�!��p՝!E�Q*vwECo����[.;U>���f��;+���X�Q�[���%ULUcGR ݦggSx)+ R74*y���kMT���SxЙ+�#�5P�q>߷��c�X��'�|"v@�� |�Ιw�tÁTZ�M���<�,��pV����z�D�#��L���1d�2����HWv��:c�r�m\�V�x�x�p�v����Z�`��B��7�!�������kH�H�͛,��(8��~�z��R���w�$��փ�R��
Ji5����^\���䦝#B�QUl[]��ZSO��rN΁y��a��
M.��:�P��&��
rN�i.ؗ��d{'#^9�f��%����5�MkF�-1:
)y.��j��;&��C,C��#A�<lؠ�i��m�����we�@뱥���`
�m���BrMR���U�(J^�Jj�j���a������);�K*ݲWp��2:N�6�RSj���$W�~΃�r��5�̆�ROq}���y�w���4LB��f/t86[�$��r����)>��#;,�AE�D�%�����W��(3�ʰ&G�\��_\�z0��=�������W��ݒ�A?jл�����8`�$�
��
��D�/.����	yX��|�Q���6F��C,�3�&�5�Ow�÷��w!�Q��P;7�H���"�:lgJ#��b4�DV#{L�w����{ޠh<U��#Fzl��9���C�Bp�T�?O�<Ǩ���"Ϩzd��>(�W�@�r�YF���C�(R�mqL���
L@���/�=>(��dTqT�	7��	ş0��5���7��X��NǬ�$�{=?l�"w*��=mՊ^���-�ȋĸQ���خgk�*/�<��p,�F�Ylg$3S#�x�Rd���wJ������P��HYlԾ9�S6�Z�l�.pL�k}�:hD&�'=��B�N1T����D���K}߶F���|,z��<�$��r�*8�9`ƔN�{�Ng�K�����*��MWx�G�$���i�8(�iL=�G<19��^\E������ǈgӾ��a�d(.W/��Օ|���,���8"�V@����>.�8Q<�Bz)�>�^^Ke���Iށk���'�	�<:p��>45I9����}0�U,~c�I^K4h��Q�D��G�(�R���FR���ֹ���|<+��k�#�>-@Z�qN0�Q��i���v���؍��۾_�w��c��s#z/���,d2�7�j����H���y��G��DIފ0|x7#�gP����h�q����YqWf��ث��z���i.�`��\��`�l�{�V��>(�H=��8r��:��5�{�f1�;�N᯾mV�!�n�"��OP]Z6u�6��7l%�\8+d�����3�x�1�NtȇN�Ȩӕ�Y�2+���5�=��m2]/P����ӄ��C'�~�U�������Db��x:8}��.�\�˕��?G��#���������Ѯ�#�Ӕ8��
$=�ANE��& ���ۥ�]����n�7�yG�tx���=�P�;�HU�d��WxEr����b�|(�A>��3��YxئN�n��;�Dł}}Z%{v1����G�8xȎ���:~��qq�z�G{�|ayd�ͯ���}Y��W<��L�V6l#9r��a�����u\*�{�Sd��J<D��H��"dj�tU͟}T�]��}�w�D�M�}s�פ$h	��ע���.��ک&�"���G�*����]���1�����U��3Gd�[���Z�i�%b���E��7i\�Z��Yn�>�
nn���&�'�j�tˍ4S�BJD�'�U�}��J����(lہ�1��{��
�#v]�<h�)��:6=J|��o8-�,�̇7�ǯ&\
�p��l<q�z^�r���tȨ��% T��.�Έ,��~U�tA��)�G~����~(��z}�,���3$箨DƒeF�*�O�����3���${�Ed#X=6g�GP0�t���D�ޡ�Hg��r��kt�F�ʸ}t<uF2p�����OA!�xf�:���}}�(\�S��8Z�Ίrˈ�7���&�1���Q ��"%�f8�'�g�iY�Q3�r}�`gAz�L��?W���¨��+�<MT�Qb�C�3q����_O�ł6.��PiA���8�6{Y�3&��-�nȾ�jnb�8[I��3+�M �;�`��U�=��܄�6:�o�us�q�WV�Xc��by�I�e����A����chtԣ�7���Su0����pd�^t;6��%�%8g
ؘ���#��鸰���~��T:���E8%ʙ#�B4���j���)��v��盟>�5�FlEd�L��X�����I�S�ǌf��x9��������|!H�YCn��;���PM�S���7��׶��(���GM"<Ut���P}E1����elc�O�v����\����,H�r��p�s�JԆ~���7ɠ���Et#�^	��*���"#���@��N�{��ow1lm�*sޖB*cq���x�~驪)/u���x�z7����B�i�܎ޑ�ҍ�3��FC��u~f���ו��]�|N#�k�J���`+e
O���%u�m6���	:,*7��}Ӑ[;�B�%�8L�y\t��'��p��C���K���`�U4ج������\,-��E'��y]g5��=�Z�QX�I>5�GJ��g�G�n��/П#��.��x~Ի���[��F�_��t1z,��-w}k�;���k�G���Q,�����D�H�t�a�fN�j ��ܼ�1�#��0Y8=��W�p�5/u����Qy������������f��'�����$qhk�g�B�O���˳���e^ЗbjGz(:�z"g�2�̛O��E׶5n`rQ\G��͚7P��x���fĲM(.6Nz-շb��wE'`?��Ƣ�V@ܩF�zzt�uz���%^�� �{���,�������L:��Y07
O�ƵI9�vU�~�#��d����n_��P���0�[M�װԷ�n��e6L���v���腯ז�*�̆d�H�k_AYm��ܑLZcSx�f����D|��+�G�3E��5˥�
l����w��r�"�t�2z r��Gw�=鎩��^�orP�q�92E[��g�(~�2�᲎�;u[�l�{�����a�D�W27фW��d.89��b�K��v�U���rƻ9y�|�鍇,����:���x�߳�;�̞�a� ���9*�Q@�^i���:����ؼc���S7�M�c��!�j(�D�:�/�׊�xU�2��/xx_�k���Q�(\}�XXcL���*�'ҋ���v/v{�=^�8����RS���n�5r�籑�ά�4}�6�]�}˷�z�:g��3�ȍ�]�$�"�9d��K}J����f���LO����2o��2ly�<��E��W�����
�y8}48�U����ՂrC��3I�Vں"ٖ9EH��V��3$w%0 Ejknk��;Xח��A�?3�X�4k/UF|4��UzG�=��3�}������B(9>(�[���٣df�3��(��m����8�)P\O�L�rȯ��p�L�W�4ȫ�&l�K۝����9�VM8q�g��"�t�²@��h�`�^o��x_�]Ti�'�����#b�i���"R�3k���K����j �~�/�ǁF�d^9{,�+�}��c4��Ǯ,���*��W���#�:�T(���f�~�Hbt�a]a�}�>7�EW�Ua���(;���	iW�_�i�UGF�.��='��_��_N��FT"7b�'��'I(���h��[w���>"W�Mt�ݎ�s�C�_@�{�j"�Ꙓ/�~��}2h����_m���Hз�/9�\��45�1.��Y�=�Q�)�q+x�E�g]�*&뼃^6��ҜאF��{���r���	�y7�f��������aۀ�n�Q��;Q��:Ӡ�#c�!i1��<��kL�FǇD��2|hD#5�Z��%П9��)ӆU[~�Qә.Wn,�,�E��*4��, �|*ق	ă���s|��d��t�6���ղL}1�{���@�U��%�
=��B�a=�<zI����t�͑�R�l�qS#%�t�JI���F��9 ���d#{�٢9��l[�WmMw���}�@��н��q#���$T�]�Q���5�96��A@������'�2z�l"g����(��<sV�o�5om�[��H���<Q	���T/�/�ZzcMvg�=C��V���쁗�}�Z�k����+`^)q�>WF���5�,��ǜ���`;�@�t���'���,��tD� B��+�u��9;��)�/���{5�'{-�zE�2�9��`����2���@�ۧ���4+�
nYF�g=�����~��W�σg˔��틂�ت��L���NRPw�I���o����#�t�A�2�K��0v*�2`f{a�}h�¬k�<(��T>��3M�ҍ�%z0͹F����=~���7>��**`N�A�>*�r�2����)�z,��\X�ÿwj6X��;�_E}��K9�GJ�gE\��W�_]������`�������=��F @�WP�=>(��h�N�3o��������w`z��gu��2Hy"�d�;�;׽U��/��!���Hg>P��z\�N���h�)��R�盺����`�G�(dx٦ FzY������pMl}��tZ�Q�9'Lq�"'��u/������2��uX��uN�ΎK��ݗF�1��] ����]�(�&���g��g;�����(�T�|#wL��P-.�/�����Ԯ1��oڝ0f�cZ:��:E����W�iLl�[]FtX��~*���?{�y�{�}����j�g�V��z��LEWn�p�p�̲���-��E>�\�B��4bE��-���硼�ZA��*���;;�l�ռRB�.�=��>�dJJofU��(��zxIn���V��!sѸ7;�8�Z��u�v���Fv2�H�7�uV��Wտ[����nk�.�(w��B�z�޷�+ �f�=����2
J!Y�0+8��R�5�v\��v�݄��t*v�AfW�[g9r-Q�N� �}�3��E;�1t�\ hƬgA���wHA�����+v�Z6H4�:�m�^~��e�x�L��M��@(z0e����ӣr�r|9 �ڱ�t������L��V>j����]ۍj�:��P��O�kU��
��6A�u��V�T����V:z��.�^Ɣ���b�V��� �8�)������{b��s����ƍ���2��"Vv�A��f�q�P{���\C���MX�W ��3�ؼ��9VT��&�3��p}�g[U��n��
]x��T�f(y�so���mޜg1��HZ� (lU�[H�/�$��t���Id���A+Q��n
qC�f*Iͻ�W(s����v���q���n���S�D_(G�����1,w.VE;˾x�q.�)4�ޝ]3&�!Q��r�]�(J��e��V�R)�6`�V����eO���r)Vdͻ�
d�Lw�붥����B��ř������Q�m˚3a+m\�rN���������;���CȮs)�t�+s���v�����#��N ���]����0s�����Z�0Qʹ�N�5\�G$5�J�V�K���4��#�s��'5�-�����94�(TJPΨtP�:4]��9#�Ili�rk�������J�Zm�s P���P�NwehK�B�:JCAK�֘�HP��r^`oeo]B۬���VMˬ�mNP}�(h�Gk�fM�P���ᵦ�S�M��'?YUr�	��g�Q���S�C0U����}�2i�>��ĖQ�@LV�F�hd��i�I�I*��fz�����y@��xנ�	��_d���l����D��;ה���r�_������k���Ä���2���8�����1���_B$�g�u�<����d�̎Q/�7���v痎��D%� t��~��IHR<�Y�E(��nu8�M��x�K��O�+Ȕj�F�0��(��G(���h�vgn.�8�a9ꑘ��5�w�n$���:��d��Î�eB�3�<h�L�$�T"zx��*4��n��f�=��^���ʵ�lAtL��5H����g�b��jO�Q&�H~��n{����ؾWW0e�Zt*o�nr��͛ab˴B݇��I��l�(Z۰�еⓗUw%n���J�/�w,3t[{��5����9�b�A\�+1�~�z��S7j�j��>΋�簓y����"~jYj��݆n��'ݞ[��q�F�_�W��Q�ކYۄz!�JY'hz���qRs�w���q�/�"3�:�j,�A�'�6�l�1�U�~�~PO��Ƅb�u��~ta�%��yV}y4��~�y�R=�N���\�x���1]}�f��y���O<|;��՛���}�{��x�	ĝp�C�q�25d�:�,FMz��{{מ��F���&\Ӂ���
T�c�Q�E�`R:�����H�'��W�E�&��}�н�P$���@�XL�	��V4����=1Ǩ)}��,�.�Tk���z/�^�~iU�EQ�x���� �w w�&�A�}RWF�ɸ}cN�X eqZ|m��j�Ļ5��gV�a��=��f�;gG��;g`�l�37�һ�LBB���2_��A��̚���`~�gP5?~^��3�����z������6E_�CM�2l�<L�늸����^���1���g���:t�IM��k�#*�Dd���&4��TL�����=
<#�%��2��s
�>v4�쎈�z�{ݾ٥>ޭ��G��PG�߮Gm]25�p�ҏ�M;D�����g{s�J�D�?�I*'�6�#>��l�`3(���f40�<t��� -�SӇ�F�<��sǣ#�q�7{y�*� �t���D��"4��nc|�V�ޓ�$S�y���p�����G������Q*_u�F9�^�Ӗ��6|ᝧ$��}A��B����B�$;��q*�/�2'�˚q�p����	�x���j�Zð��f.a�Mď\��f��S�rJ;�X0L� �N��IǲV�)�y��Ԓg�u߽M��_����c��-t�� t�^1���Z�wS��)��SF����$��z��O@*,('x��8^��g�-���/#L��7o2���3��6229I3�N��\X�P["${����F�,���ӆ��H�R}�/���O��x3�������*qch=4�+����h\�z9�%Me��Q����҇��������% �S��A�<������i�1�H����^�eF���`�T2�	�l�ʃ��CD����Gz0\�voP��F�H�>�;�m�8�k^o�>��%D����U����F)�C���C^��Q��r���'�zD凌q�	E(��ϡ*�K3CiΖ�"e��(��9��-����M牣��'�NC^wC��^��m�����Rj����\3�ޚ�s"dȩ�L͆���hG{{���bP	t�'���P�.�
g�}��7��'������G�j7=�σ�I"��ǈZ��d�/`��G�j�-{�E�'���O�x��J$�s�L2}��y�&�,��hݺY����
ޟ�����qY٤ F{��c�Oz�C2!�<�]	ǲ��T�;�t�ۑ��h���c��q^��șW����C;"P�.�a���"��i�ҏ}���`��L@��إ���$�D\|��Ɣ�<��EȪ�"�5�y����%y{ٯ�y����\4~\��}�,vL �Y����zu�w�����=��;/i�Q�M��G�J�'��b.&���+�z�M�gE��"x[�!첔�y9©G��(l���vݝ+i`�=�XOkgf������,�vm��7����ǳrD�eB�L	0P�[-��;C��v����]<��,
�G7�2aEu��ޅK3y�p��:�{�D�q}E{�Ƚ��<Q��Z~N�I1>��gfb�<O
�	�B�K>p:�D�d����߷ܣ�Y��p��FP�B8��[t��]yW�ƌ5�J��Ѿ~����B/U�LN����=�H�2f#}�u��Rm^S��xzF�H�p��(�U.\�,1�`@^�v�b{��{�y�4"=�e�z,�P=��j$>�A�.�����f+ٺ�(b �X"����r��3��C.��N�^��O�0��f�ะ�l�$e���&��!}��4�(T��l,BH���[�7�h��`W�9C�F*�QTMp*+YҐ�ڲ�2�R�'�!zd0�_�8��<_tٚ�#&���)�d�<n$/v�����Q�ޔ���'�ur[{&�3,�2H��<2��%f	�On��l��n�3*us�����QQ�rjk��>FOR������c��������ܼ��4��'y�<8�E}�ǲ8���ܢk���M}�(׺lͿA/�v5�D	2:�c�������z�5� ��.������^Bw�q�^����t�p�@��,'��͆
;+��e
��Rj��z��|"��(�8��y:z�C���3�uF�I��euu������>�~�_(gnX���g�`���
��߇�\׮o�/ºdc�����d"*�d��s�"�G��kuo��O�v�}qǩK"w�WC5�"�y��CT���Ν�>ά����}�����
������.��:p�ҍ��H��S����C�B�� %�Lǥ��!���B|��]q	ȃ���]<�W�e�h��k8��W��%����ِ\ͪb�D�4f���s���q4���̼<�8�־������>��5�0d�
kw�9��?��f�e8�ߠ@�@�����yC�+&�S�7N��� ۂvG�Bj3r	���d�8B�F�K���-�Mf��[(�s���*<�Q��;6GMnһ�^����0|�M�;��Dc�zǉ�' � �ᐶ2u�^�G�}�.�F �ᚹ/����C$�S$r���V}&�緾�JGP=���4�	�ـ	�/�Վ ���W�+߭��������ǎ���U�CmH�ߦ�<����W�I�z���C�"ϹH?���5��6����g�[�~<��H�����xnP3�|l�C��ȥ��DQ�og�w�N���ǽ�=��u�&FG�yWB+�d�N~���-��C�ѯ��]����1�I�fY�u��j�1D�Z�հ^&9�<S]Iw��	��5�
�;b��̚5��ۓ���Bn%m��ò�R���]��
:}S#=a�Ӟ�sЌ��,��Z���䢮\v������-�C��ب�p�9[�&�Q�R,�:����s�цOXzp~�w�d�-]��p;c~�1M��U�[��W��/�#}�Ol`�G�L�||QҮQh�%��^���	�����G(��F��(�Io��D�����N?D'm����ӆb/�(GO�}��nó�F����p��$_{gyC$\��Mx��R���ʘd��ޯ�/:k���͂\IW�%L�̄l�#�Y�����.�dZ�~�ɓ�xߌi�[r:���f.�r��F�fQW���>�^įS#C�xF��`$��,^��xՊ쯳5�c�Ƨ�8)���ճW�kW=�ɝ��n�% &��nNg�U� 
yczhݝ
�t��,s'� �eZa�L�b뺍��Hf�Q�좛2�}�Ջ�o�x?������"�0a�Oj<W����Y��A�.Q�yH�Ez��g�r!E��P�=����ӭ5��O~�+�E���Uy� ��P����T傛���¯-Z�eDp�8�E�Y�"�_���e(>�>��3�Nr�=��n�w�>R+}aa�*z,�q�FtK��<����}Ə�jF�
�T����Q�����F�Y��r7(r�I�r��e�.���1pc��q�J�0�/���������7�^�"��B̟8�U5�Gt:�dޯ'ț^�%���P�;쑵�=�t�����P�`!�=��	��xm}r�=��\��Q���z�Ǟy���G�?)� ��*?��UU_�6T9c���@@C���0zT>��H�����g}�ǐ�o�����u����Ua���9����1�����UD�"(��>��@�7��e��~	�-גg�-��֛���AJJ��֪�c����2�q`����ڪ�Lqt��)K�f�Fo�,�X�%�ۢ�2ղ�٦|%���f����i�M�A>���׻�½�*L��HA�FQ?C���-%ݳg��<��I�S�dO(����v�����b�ns"���!��K|���R�F�d���.&=r�N�/ڵ#z�b�G�loAo�%��|�S�]��w��i[��wvJd���'���%�V�k]L5^��r�G~�� ��U ���]�
�@( ��H�����rn?G�c�v��c�H ��!�*��,��ǋ���}�0�pR��wZj1:�[��{������$����z�<��k7v-Ay�5�U��F]�������]��e:p��bȳ4���xuw���u�18F#��tim�������},���"�D�$�u�)Z�}RR���M�p�����~�6ʊ�x.ʨ���RSEa��V��8\�G��fz54c,���z?�C##}�*&aǅ�c�C�W� �!�_1��]&Q��ө}z�e{U�Y(�+21Mqyd��(��jfc������CT����yk0�H �`�vI�T���wB9(�����65�m��q���8E�9����,W��R����=[��ʨ�2<�����9����H �'|��
������s��Ƒ^A-'�.�i.��3�jpl{�F��6�K�-q�)��I)x�Ͽ�^K�]��Q��9�鲌YsF�<�j��SK������7c$C.Σ��òg��v�u��4S�2�t57p�U7�������$�>����HA�)���#JH�I���4�׼��gK��20me:��&Lq����P�;�^;�|Y&┤�r����f�6p���.�p�!��A