BZh91AY&SYZ7r>Րߔ`xg���&�����   b:�|  y�6��)+5"��m�[&)EDZ��54��SmT��	KfB��mi�֬))iU�L(�SZEM6٬�hm���d�M5��֥��ã��-@(P���ie$�ͬ5��[j��1�m�Kh�d��ZV՚k*�5m��ҋU�4֭ZVm�UMiJ�Y
m����m� x7U��Z���jk�)ESi���Ҋ�M�Sf����i�m&ն�Y2�f�-l��ԚMT�SU��
�U�-R�F�k!Zj%A(������5I�   >���uF��մ��n��w9���5��nεN�AZ��u&�ݴ:�b��k�[�M\�{�z��mh�Q[s��wV�t�v��lє����UMm|   -��B���*�����w�<��J��=�S�R%+�U�xJ��R=��EM���N���T�U-�\�+l)=6��ﾯ�%}���_;���	t�O�/0�%!*ХM���-k�   �{���P�;�=ޔ*IH�����}%T��>�����2���<�*T��w�}��B��8=�z�i�eko�W�P�mB���Em�v��x��i")y���mP�m���2��f�� ���]����w��
�(�+�U��x��<��*#oo�B[�*���ݕ+����^����J��׻�Pmf�Է{zU�T����S��I��fh�֪h%�j�V�@π��=U**�����Ɨ�*���w�Zz��w;�˞Q*S�y�MG�;��UP؞��{j����U4��g�R��T�Ӻ�EU{7�oeZ�kR��3,̉Pm���z;>�Yj�{z�yM[=,ҽ׎z��R����<��G��<��UQ�{n�J��Zݮ곔��=��*^ڶ��g���k{4��W7���j[oI��%�TZe��[+L�j�ֶ� ��_u���]=���J�ٝ�mw�R�m�#wo]]r��z{v�G��ǫ�)P��x�Q*�{i���u�����J� 6���B���R��ж���F�V50 �� �O� �Q�Z�kkw}�p ���=Ph/^�Ȫ9�g@WAr0�
a��@u�� 8���u=6����m�di��V��ƥ����� ��Ѡ�W��� ���� 竞�V��9���٫:��)A�{��x�h�T[8s�U)����C�x�ͦ�3*l͌��-�e�O� �{�k��F�N��w���zP
缸�Z�����Ӧ�(�&��YOw��
�w�[���E=�{�@(|  �    S eIT�       "��b��� �  4  OɈJU"0  &�&�` )�M	J�4B`	�0��   �?!0�UH        ��H���4�f���̣�(�i��&���������k��A�$Q��;�L�yI�}��v|26�f3u��~ {���NU<{����=�|6���ٳl�鿳�~��ٶ���8���[��߿����߯���������7�m�<�mg�:����m��m�<�Ϳ)�lͷ���g�&�������K������lo�M��6<,ُ?����X�}m��Ca�[m����6�}}}m��0>���A��ُ�fc�0�,6>���0>��>�f��F�m�D��m�!�E���m�}�DfD�6�#`�#6�b>��,l>�m��E�m��c{,1�F��-������&�-��l�豘�!��-�7�3c�D3�D�LϢ�o�6�-��o�È}��C}7�6}�D��[7�� }m�X�D7��Dc���XϢ�����y����.�����>fX��k~��2�G\_���&0ӄn�Y� �"I86�ݬ��w�z]Y*��纞G�t� a,VJI��8V�������J�21����wq�n'���{yx�����T��w��,�n���\K6e��S�*\���M
_L`�����	��'P��h����/ql٪�YD>#N����:J�ߛ�ʉU��mՅ[Ɍ��mjU�h��F�V�K��0��&�:���Z ������$��:�.Θ�b%��TB�bx�&؛��y[d�O�D�v�JVX;��%�S_C��c;֟�����	T�CɚwL0�Q�kP��ϢгE=š�q�\\�+v�4ĭ�N��D@oVҊ�;�a�SBuk*�An�z�j�%�)�؈o�FA��@��Q&��Y��yW�[���P`��a�W�7���u��T�U��PʻCܚ���e�cʘ�C�726A�n�h��9�]��}�ջ�D��O�xxӾ�vM�1^r�^Vn⎅�$m�Y�VMOR�zWՈðV)�o#���#B��.�ئsU�oG`x6c^�hn�ڈT F�+&��M�'�3x��]��a���L�DXl%�8��̩YF1j�2V��o��\Z�f֏��M���b�i���?�.�.�[{���G1��m"/tZ��Y��8r4�.����NGB���C �#Oc����x]�W��
Hm�V��׳v,]tm�ӬU���V�4�����Q�0�l��2��CjY.
z�(U��R�l�.����iU��������r�	W�a�s&K��+Xh8�=z.mJ��ҏ+FRW3�s��Ѩ��A����_k54�;o���^f�55��j1f2�
f�2�Q�b�rõV��ʓ�w���`h[Im�L���lK��M��B��O�]X���:O �QKr�D޳Z�eE!�S
T@*��X뫺��J���0�,�O��:۷	�zSRftь^q�U�dc�=D��Z�b�o$h[%`D���c�
*o_�U�ՊO$t��r�w{�%L�+�c�K�}EN���t�g[흕Ө3WLeWt�V���e�S��s�n׼$�o[ִ�4٭!P�)b��݃�7�{���"��D-���C$A���=���֘m!O��y |��Y�԰d��O^�jd�"��S�I�����oi� �i�.k���݄���˝dJy���a�B\�2^b(�]�&n,�~ئ������/V�u�cK��h�{N��׼�M�U;T�TF�"&3lɰ7�\:��j�X/k#,���*����q��WA��M�nd4-R��la��ɬ���4��:}���6ܣ��;tfϗJ��%��@��TL�[*Q�A�y��xt�t�ۊ�����I�f"�������*>���x�+�YyW��m,�x�N��i�#�1�u�l����U;q�ڳs]���攱�G19��tN�3*O�e�&�J2u�0�X�H��
�Am�0��*ֆ��X���P��H4R̦ݼ1i�Ve%�A��`1��w��FfĒ�l\�7�J��-J�2<f������SDr�PT�GQ���C5Q�n��2!�h�SdU��*�La�P�i1��Ѱ:H)�Ӻ���u����y��B�@���s%(Zt@��q
��CV昅b�T;+6��V��"��kL�EM@;YCKB<��[hkٛ�!y@젨�F�F�Z���S\zoc��<eʕ�lZ��� ��GVQFիvpF��f:��wr�[�>h��ae��6�*���������A^�,X/kS�.��m(�:�N���1|�3)h���i{VF��3����.ٺ�5FT`*+��e��O%�J��YoQ�q7���e�5���Su�T0U�3A��RǠ���(f\/�o1�^[P�N���N- ⻤-`v)�a�=̫c�mn��A�_0�v�.v��5�+;#|0M
�J|��|(�q�N�{�]*2����.�̨��M�ɛ
���+كfb@�PU�m7*�:Ì�ieK�0�凷�#ŉAM��c"?a�Z3e����:�ّ-�M�
���8n�_�GX�q�[���CdZKIDU�����+*\/-���[��ӯ@J�i�ՙA`�^�j){�jAF��`�R2�M�J�t�[M�ȥ%l�U��MF
�
rKٛ���ܴ��j��S���U�VP�������j�͕\՝y|���.��7KLX�F+�e��ZTƝ��^ެB��/�/�ʸ�lSH�C���g@˕��Uf�����4i%I�U��)�J�[L�Wie�+l	�6�Y�#r�M�c5��/v�<��h�zV���<�ScGpc5#���t�Z-^>(�Iw�Aok[K3Y��v�MЏ
̡F�!�nD�01YݎWK��xgc��t	�P�,;��Y��r83�r[��+~����@�u��`�IQDPـhU�!����݆խ�%Hb�� j���90��n���f۷k\ee"[yYIkm���WtH{6"+h�����E���s�*���$�>R�F^lΠ�xswV]kmRX�6�h{����(��5���r��[�f���Ta��j'����e�����J�m�h���F��fV��QǢNJh�a���&�42�[�	9�L��a:D)��5wYR�S�t7ƐV�
�}��+Rk�xv��H�vhܦ��H��R6� 3G.�6�{���F�������z��ɬ��9KRt,�n�.��r��i�#�⫭����ٌ�%�k*�n��L[���Ҷ�2��4�k)�7%����cy�'l�t('�f1�I5�lE[�M_u�V[�M��"���20�4V�Z5�5�^7��FLqX���J�Ff�	8>�!�e�V=#�h�J��iP���ըtH�5#4�]�[��$���rQěy�YEM��egu[J��V�qg���YY{.�)m�|t�t��՚�)!��V���hf�̗��GZb��(Ǩ'0��༲��XB��"�&����������uT�R/FM��JE�S�d�5��+kT���R����8PO@�/~x��R��In�ڡ�Y֕���2��G�X���:�l��a⸤�cM�#UW��rA�ykŎ�h/rk�hn�B����J֋�B�E�j�SSpɐ��V
�z�f�^�`z�L��Ӳ!�`��dÕm'G �N���D^��^��G3[�&�԰�4)��4�bV���V77ovˤ��5
�ݭ��i�4ّ��T��t��v�m]K����
�"�ɑ	��
�7p�E�d�pj{�7���Ks%X*+��v�l
��¡��ʲ�����Cj:h����c Y�X�-�c^<����흂1Mm2U�ՇZv��kE椵���-Y�K&e�ŦT��Go-8DܑGXLU�Q"EM�ʓ�4�@I�
4�5��7۫��-
�k#��;)�S1݂�j�j�A�[��/j�[F3��J����J!�WY��1�&�RlM�l�1:��nl�L��y6]րko���d�c�������܀l�6�Hn�A�V�X�3h��;Jٍ�f=�k�b:��8TU/%�q���]+�[����Ip��"�Z���f�˼+v����ɺT�˧����J�J�VP��Ȭ%㙂�X@�cM=>)8��׏.��v�lX�q�a$dq!��ue]�&7��:)e)zb�]j�1a��v�O�U�:K76��n��p�j�[�ZIf�6e��܉�20�'.Sݺ:!��J�[YL�rV�ڕ{[�-���R����)V�9l��W���ܘUu��oJ�VH���:�'yz�̈́Ʃ�w���U
�8���۶s�&��DTxbTj�EB�nu�A�t��;�#y�	��i��u^���5=���
�sZ�X7���G��K�ئEw]`�Ǣز���rf܉셩��d�Oe��(h�+T����>�T~y�XJg��cZ.�w��j�<F���	z0逍̋����}����	�w�c�������cG[���+\ƋQ%�����"�Ő�7�m��:5�mӓ�����D�{��@����"4Yk����òIZ������vڔ�ҁؘ��8&��˗�
y���%!1ځ�"�+V�4����5�Zf��c����R4s`�J�h(^����X�O���Y�n'kFj2d�h�6.��%@�ke1q�í�Z
ݭ����@�=�d��,P�n	f޶�'�a�R��cN�V��PL�:7�4�6���1I��%]
�ȝ�[he���q�/#���=eK�Ow�QO�K�=�D֝ɪ�z["N�`�ާO޽@���L���\� �l:�[K���X���fnnQ�R�E1�͡�U�0�3i=$Vշ��E@��N�Ѷ3oNj�z��y����m�%�IŎn�&ckݛu�e�stmk�&���a������[g�[e2�m;w����V�q7q*�M�z�������K%[��V�\5)ح�Z�x����
�{l�N�n�,��ӽ����G�ˇ9�MB��[��e�����v�r�j�vJZmc��fmZ"k;�+fUɭ���c-�Yר�ӰU��L�q�U[��:�[j;yeͥ�1�&�{��%5���E�����`R���lV=b0.Q3KVQt&����"*N�0�[F�_Q7����D�� 2��Efc���Dh�3bJ��r��8���Zl��&����]�pA�(n=K�C);��z�׃sYH#&����L;.���u\�5��a5�qjV+%YS-͕u[65J��T!P�6e2^��(X��Э981�n2-޶���[��j�-�e�ٮ���A�/ۦ�l*��Xt+faʰ�+ZpAw)�V����mok.j3(X̑36�&kf�6��1V��Y�p+[�N�%H	�iĻ/h^jT�0��0����.�����b!0A���n4W�C<Ȼ�Ay�o�EU�y����An�m�yR[�v��ۖ���	�R��WBAP!k2���.��9��z-m8�76#NV6�uަT��D"������*�iQ707]+f�����f�,Ŗqj�[[��#Hnb�n^؆f��+5e�@��P-H/�-b�H�J:�cl�֨嚟 �]`���є 64�OSM�G0�1Xwp�l*����;�q�N������n��{��剎�VV7B�E�q����6����i@j�MS�����d��t��_��ܫ#"��+Ow3�&>7�5c)�i
|D��Ч�+o7rlE����n]��r�ؤ��
1�a��,�i:Υ�Vs���bGW�>%�6v�!���#�n&�JP����$Y�mm�[N��Յ%5����;��OR�C�.r}��r�ևjjZ�Ax����w��=�w���+��)Q
��c+5<;���� �jb�f��yJ�F-qnj�{�(2���r�֚�jh�J��jl��`ǿ5o7N��k-��b��-'�)WJ��� �j�"шG�v^��wJ6�c�yWFo��x�,�+v�%��;5��k��i��66�˫��X���^R屔V��:P-��͗��(����4,d�;0P�t8�B��k�,e�{���TR؋n�]�A4~Ԇ*��+6�ֺ�7��Хz�$�Õ�e��
�q��Ӱ�,�ͬ`{Ql�F�#J�3�f�6h��V���%.�� �pI4����6�GB5��.�*-'�n!LH�U���TB��ճ���0�cL�BnY���8@�����K��"�Ǌf�:��5a��3#�Rm��6��	'����ԝ3�f��g�����CQB�wۍ�ԓ�<ϊt��u��b7FU��D^��
j1�P�"��ǒ�b%Qu�`�&h��d��{v*)����B3��y�AX�����-��ս�N��[f�s^��Շ�ʴ;��T��l[V祦8�A`�m�Đmk=���'s4�Ew�`�����w�f┲�D�W1b�gj&�<���,A����W��F)ɰ��Z�%��]n,F�;k]7n�(���U�l�{�$�6����WZld=�:ZΛ��`-�5�Α�-Gh�l��m�KG�z���M�R���ѱ (n�T��,H]�q��r���� A�G��*��Q�M)�=#��S��&� �l��j&�ȩ
�����6��qkt4D6��\�d�Bɛ��Z���e!��혤�cn�x�
9|�ͧ�Z�͒�<�Q�F6�$�(6���T,Sֱn7��tF��i��Lͫ���5�R�)Lڬ�J�Pܫ@�v�QӵaQ��H�����aE^^n�;Wm�m+����3.��t���6UH�_NR��AB^AX�֙AV ��̸m�����*YV��:��o3l�)W8���kȨ��-\�Y(T�� �3E��9>�AI��j�_�ӭCi���VNV���j
�H��.��x�v�/�.&���4�Y���3���ڧ�kc�-�c��s�C��ݜ2R�5���:OQ�Cm:5p�X�f֋Qͱv���Ct�!����MiS�7yƆJdؐ�ަyZN���ʋ�@
Xj⨪f�r������IZ�sa=�;E�=�d��һ�7��l[�g��a��ׂ�a�Wy�0VT��T���u�U�wQ^^�O`�k#�`2��3*m��g�ZEl��i;�M)�Wz�¸����#�̟+JvmCVM2i�YB�48�������d4��᭳�Q��
�8iYB�4���=tg�#l�Y�Ȍ��B�4� � �(Vq��5�f���Z4� F�9Ɲ���F���heP6oՇr���F��E�%�#t��!Ы�pQzj��#X���~[����R������_�t���*ڪ6���JDL��c����%�cv+P��*2E�7���>�{|>��SO]U�������$�I$�I$�G�Np4.��I)�I$�ʒI$I$���N���;V�VX�iT�@"�J����v_>�(����!B��e�щצe��K�'f˶�y��XS�f�����I�����Ƈn9����w��Hp�Եd"�P��ո������ޥ�tH����RZ�|^w:�} [��gp_1ie�ۗ��|�7����}�V�6�Z�6�^��r��t�i\+R��F�ʌ���\�Mw'��f�� 9>3M�2evk9��iM���$�htz�gBV�r\ed�v�W]o�����'y-bmf�;!!N�wn�qv�ǃ�F���\��U����0C|��%�<4s�DA#B�$@�Ҥ�6f�#���ա\DA]�*ƻ-U����c�Sfص�<v
�E#�h��)�(C`�;���:���V��S�\�K�{V-3:Z���gkI49aE�3p�ϣČG�%��S�Y�k��Q#�u�ۈget���G;�H �pcS�/��5��UEq�zl�{|&❏-�,�a�#��s��i��Z�&7�ƕ3ܰ�W6�b��u]X	�wX8)�jΥ��\U-Iq��8Y�˰0Y%��
�������G���l=ۗWf^���vr�&��>V������4�9�d{�������lwF�#m�BI�/3H�L��r��g9���*�D��z�:rd4��k��]w�7n�IF��3��߶1N�#]�l3���	�yd�)՛��d�͉33�6��V���1\���bw˳���PV�[wDDm��^KK絻��ʻ	�Iu�0f��\�2��o��8������y��L�Қ�h)��nir�[eU�j�)�{�7B�M���*<A
oS��J�;+�����-k���H���vSĞ��JV��u8�WqǊÜ6�j�5*r�*˻�e�2��A|]m\m�]�뵽��q̣�{SF
"�][)�-4�b��,���I����܈k��y.�1V[	U*bY����Ҁ\VU`�5���[��r�����
��,�q=�\������_5�r����]�O6.?�l1@��ѥs����.Y���VC7�S��]�-�	ٳ��LW<U�1�W��p��	R��w;���M�Hn���	e%�1���鶚u����bxВnM.�aƫ�v���|�C��ml��i4����&��yx��� �����chp�W�����D�v�zW��3ybd_��Q�D�]d����m&�МY�e�ܻ|"�wM'nWorw>{/�/��Ŗ����zl��X+3�7X�UcT25�ڢ!��U8Ty�Ʀ��e'\�:���CЇ��(�J�_hT��D�u4��vN��^A[jmĬQ*}��[3���q��u5Fas��4��`"g�˶+E�G��&�\#ٮl�����a��c^�K�a9�[�[q:�l��E�&�24���
|zh�B�+���#�K�8�+l���r�MQ[�p��6-V��$�ĝu��2,�:�W���(V��ko0��g��t��CO:Z���ү����}��.�Cl��<�]aǣ��F��x,B\}�����L��v�=�fRzù7tb��]iQ]�kt-�P/��ev�Պ���^_k��eα��R�3kf�Z�f�q�p�<3r��*Mޑ=\�vs��m��TwV�k�{��Qkɥ�PP���j�������V��H�U��[�b�CR�oP�����b�f�;��6$��C�x�P5τ�a*���bw��ޙ��Qq�9��
�6I��-�݊'�s��=�}���4����̈́%vQp��i�ȝSiȑC0 3OLU�t��
4[!��.ǜޮI�!xY��\v�2Ͷ�㋜L��*�+,<��L\����5��<4q��N�4�ɔe.��+�׹XiqsC�h�=�^���Qw.��`��i��_Z��( e�Ҿ��W�:8Oi�ܢ��:�Rk 7|3hʹ0�y�S���jqa��z�lr�''-�R!�`�r��R�Joy�8(Wb������)<�w*��+v��jvnj�5(]�@���.fq��+a�o��޼犃r���.���)"+S�i*_=��!Q�U�����t�XN������]d�\��mJ^M��q�+]�f�(���"��j$|�]��q�����D�Ċ<�F�����$={ū���!~4֧X����bI^ev��G1͌H+1C5�7,e^�ev��svQ��o+	���%4�lY8ka�,]/��jn�~��f5cM4�y�t߆ʑ�;⻭>��[C�A����\�Z���k�Q�K!��sQ��vۏk{M�z�ֲ.�
Fع}��{�3tk�Z�N�+�N��A�55�q��=֮n%�ܳ(�b�$8��8R��)�����^�e�D5m޼�\afm���"N�U�
FRZ�Oً9H�>cZ�K��E]a͗�����&<�QVI|�8�v*�.�c�L�;x����EBuY{N��|���*M{A�]�边5�sa^���\�U6�뢬=�".%,�VD�tD�ˢ4-�c%m�K��/x%��V"���k4gC8#�H�a��e��W)n��N����Զ���B���u]vD����,ѧ�L �����­d���b��c���:��K���|9,c_-=��r��&��6bgoQܪ��h�plŸ�͵l��+����SI��(��R5}����R�\�@����wclP��Z)L1�ǹ�5��v�Δ��CX^ee��B-�؊���ciBb��Z������;�o(�oWR�nS5���*r�R讧-7�cBxn���^}�c�b\�K!�&�j���p�k$|��lS��)wD��s��01�FL����S��opuM���YQQo8SYՋ^	���JS���vGs�p�܂���9Q�7yO� 5}�v��!y�;���R�9z�Y9ge�)j�� � �{�f���-M& 	�u˚�e�=4�cǖz�����࿒�՝z����V��������u)�빓�6�6,+͝q��ϵ��=.$��C��GF�¯��%ٔ��� ķ�R3�&���»q�l���uM��Z�
a�(\�}�ݬT#�������ڹ*�il+VO�L�n7$z1��ͪ��S**���btS[.Utۻ�����_V'�; �b�2��[4
�3��Y�c#So���g�5�WMc_D�5�5t�n�,S����;��vҲ#�o��wJ�f��+���t�(�d���s��h}z��ݣ�k�s��F�e^�	���;��8�gs{X�b�u޼�t�����7J���Z��(�Y"��n��6T�����Q��er6�R�}���D�����B&hkU̫���Zo�#�U�z���ְv�%9���zw[7�a�����ӊ���b%�k��0S�Ú��kd��Ɋ�=�(�r�ˊ�l�3����5n)�i��eT�[`[��S�E/��xܻs��	�n荊�;�a�|����-2�{�㗬��B�k~4I�;�⧛�ˏ��gb�1uHm⧅&����=�MV�A��V��%�!�1��`��x��n�j���wu���K���/��)eZ9.���[[R��݋w�j*�u��C�R
Zؚ;�&#����Tnٕk��Y�Lc�y5Gn�4��Wk�i��P�:�m��v��K�@ٮ�BRʛ��"�%"�q�p��ҩF��n�#x{js�)-�\$�L3�@�cd�KJ!ݷ�.�z�-�n���/�up�Ϥ����IW���C���jt�Y�u��˪Y�r18��O��+@
<��~��E�m���<Z\If�����_�\	I�g:D�qgX�u�zj�;���s�*�q��83��A\�N�#Ո��4`X�-֝�~}@�u���I<��1 ���F�=�E�U�L���1u.�R��]����pu:�X�NU�nb�Ǐ�5����ԋ:��6IW��t���j�Yp�o/33�x���7��4�R����k�i��Y'p*+F��
�n��)��F� ���졯�uc�oo�iJ�
g���%��U�{:�by��M��c��k5'���վN��N��<��hNq;[��**�ư����e�s����6
5�-�.�Q�M�_J�����x������:ZJ`��}�{�@�o��qt5��.�I�g0؎m�w�!��rmr�L5�|�Zn�w���	�����!]�Kq9Zf�֝�x� a���=���tPY��<��+�%h�IZKa"�]�"ɽ�@ڏk���0W`��s���,e�J8�F�s�[�V`o�d��f!�*�[�N���;�ؑN�s�7�x��nh8��D��]w^�S�#���m�mp9s���x̭/��KyW6�r�M��Z��㇯g^�>�&:|L��\�-�-�/pXy>�y���4����un^�ek�"(�����
��'�Z�0�+\�ʂ��Ǯ�K&�cS�]���'�`���쩹�Ps,�ti����Z�ީ���c#��K��b���uh�$HV���B��$��:�9�"�Ӭ���ZNh�ץ����el;;i��J�}��A�H��wxb}�u|�m���k4az��<��G��G)�X9�+��'%Φ�Ĩc+8-�~��8�9MhƳ)�n]*D�n|��֞)-���I��R�O
�@!�,��k��n\\=5�
�8K���d�/��J��״�H;O�;�L��M�[n�[�s;^��k�����ۭku^λN�V�W�>�Q���$��M.*����1��O���V��uAZ�9%�2�W¸�u9jT�(oVH�`�Λ{ys��g+��������K�"-��[�Y�k5����`7gqg ��S)4�g��R5��l3�c��r�v&�1�kkh'�.�v�XoI���&<�q�Ef�{i�r��pe#�zZT����n����A�z�f_Rܢ�����ԁ��]"ĄE��n���g��Vŷ��u �T����]r����Nb})��g-ݱe�)���XJU�ٙE���0�_S8lj��9ti�d֡�v�$��Vc�W�h�]L��k�2���.���͋_j�Xy7Knc.�4�.�k��Wiլ�X.����vE�9�."���y��-�h�K�'dC�����'ا)k6��'�яs�`���o.hh�f��}���Ԇ��W���˽`VŌp��E`4����s³��5���*��R��J������H����E�}qPn#8��*�}:��"j������G[W�`�����a�jkNfu�E�]�`�E]�TN��u�m�b�Ѻ��W�v���i�W����^}�&X
e��us�iV���b��3��w�HT�9ͦ�Vm�LX�ў�5f��fs��q8�3�l��sKc5J��j��̘6�3�Nq�,4�xz����vr�;8G[�;����|��6�`����T߭��iB�\��x5���E�ݞ{w�͔�_G���`ue;�yyM�wZ���׉t���,�}OT�MZ���R�>��m���%�O���dm��ih���Zò�=ۮ˝�݊�a��ls����A3���؟pcv�D�q��}J�wF��b��W+�%s�%[�����Wىskq�JWT�6�](�q�Ž{{��Dɵb�e�.T������wx�n�x��ݕ3	˫��&lN�!�
1�/�d���C*37��[���Օ�є�7ǎY���wa* ���bЮG��^�!�����epJ���v��ۤl�����0f�}�,l�	;]�ޚ24TM�s���t�0 b������N����4�^����޷$���V�+m�锨ޘL@�u��V����¦mk�9֦�7{C4�v�{Kj�E�m���,ŉ��[�
j�����ח��P���;����*ʵ��t��[����K�ugf�]��k��aa}0$]X�U���zڲ��봅��D��{V��l�k��:֋��A�Š���w�:�ޑK5/�*�Cc;�i���ga�I���Q�T��������gw���C���Ѻ7�lب���52Q�2)��/m�y}b��ݍ�IMVZ�3��ң����.܊�[�;#��sU� � �#�>˂s´8���c�z���G1kQ����˂����d��,��H:�	uԓS��;0�Ъ�&)f�I��9�u�����^e���c#�UfCm�;��\֫zq���\���kD	m`|:�˼9*H&�RJź�஠�FCMDH�x/7d5��ɭv;�a�Z�p3�����K��7M�,��|�*��L�.���av�V�y��z�pV��X��ҫ!�#͎�W^�O	��eQ#�;�&��Lݳ{s�Ե���ṛO5]ޭ���<� 
c�Ki�B�:��J�
�z��N�O�%W�]�ՏyꫭT\��M�� ̡�7kNu�4[�v��NV���X�] t��wc6r�8����������v���ܮN�LZ����\��o  l2�V�{��J�=Z��_!`�p`�uɪZIB���� O{��.��o�_�,�D�O[��p؁�:p�N��z����$�}�T�A[����y(��n!��7S8Cs$d���\3*md��1J�Y'���jh+�'_"���!Q|B���A�!wdR��S%��=}�dJ�-�S�Pه��qk�nH�ΒM7��q�$��T�IG$�I$��D!]WF��P��\+�/�;����﷮���y1�57���<zs��9����3�m��|��o&������o��ن��~�1���������|�����w��fcfߪlc�s���~��ߟ���|{��{���}��}�wo+?�"���E�w�G�4I��1�U�`�j���F��	�)��Xrd=:�s�+�K��2^#3�r_���NY%c�Y����wPs��Ð��-D���ɇ ��#!�Y̓�G�8�Wsv�/�_)P�Ņ�X�.f8���C�Yo�P/M��n���خE�*n��E}�\/��g;�*<�Z2�n&^����h�1S���F0��jJ6�*ۏ>�o.\Υmt���nK��1�3]�w[�p��6�֮�8��2Eɦ�m}��d1s�Q�4k50�m�)F�I����8��`�jAL�����Luf��4�������V�s:��衠I`8��-l�k�;g(���/����(��LI&U�K7'dxJ�2�5u���
Z��n�ͩt��At�U�$aʲ��`K��ӆ�U��J]*����u%k��p�4����L�V��	[*��8�yϬ��0�#vR�*��������Y+n�]����>�OFPT���� ��3#f���h������V�K'I�3j�g�J�kR�ɚ�N��.�TG찐���˕����K�Yuj�yGT$Սtɡ@g*�I`���z�S|
��~pT��Rr�|y$�4q�}ɫ��`7}}//:�����%���ݖ�$ǅ�P��´��TZ�oP������]7��ݫJ�f
�ֆ:H�s��O77���I�(5x���V,2����\�fu�ov�Gf�Ҡt'G�Wy:�*y��$�,vչ�Հ���V��1���B�NL�@�%�мOA7��u��S�+��4�m��O�]$���6{%Z�)ڱ����i�;�f-B�HV���*�֯����m�\�p�S�ə{��ȷb�\�w\�'^�"�=q��F�Z�`uNׯT�.�if��ȪҾ�skI\cǹ�ap4�Vb]WY�rG���S�e�s�|��m�j�붮�R��2yʍ��TC�f��}�Y�y�x�Jm��L�l�2�S'4`���ɬ�z;o��;\�jw|\�څvE�e
����0�#�c�>d���h���%�p��8\�?4m�Mj<�u��L����.i�����W<�kN�Ӵ�u9��t-��v0v�͝1��m+֫�!
�(� �Rȫ�Jr��h�0�k{Pp�w�22 @�ƅ
�xQ@T�T���MO�rΧj�N�u�t��CzQ��!"f��E3
�	sR4�X���?�VcZU�+\����6�@^r�h�]���q|�rŁ�+UݻG�+E�]�����<��d��b�v�"VH��U��+����Yb|in�2MlL�y���1p�X��Gn��Pf��L��@�=غ�Tj�PVI �ݲ�o�ܗ�^�2���mdr���N��^��t0���#��b�X�3wW�3�2Y���˔�6YF��X��kZ�9㮗c�F)*�{9�����V/ �][��(-��.2�I}O�w��1A�Zi٥q�t�.�pWa��nEZ�۾��J���Υf��Y�E��q7Y���pc�L���'LU�YPp��z��&+��&�7gmit�&��f�:��d}�q��[�l�Z6�F�s涊����(n��q���-��t���h(�o��������9�i�#���q	cWB��{|
��|��n��2sw/+Y7pn-(e�L�\Vʃ�x�PPn�*yt���mZ��a\�tr�]�'�v��qF�
k�ޭkh,�뷓���o4es6���ӵZK�ev����eBrr̮�139��Ԧi9ݫ0�-z�IT7Ξ�}w����lf��o�T9�n�bMꝴ֠���mHv�������J+�5P�9�W���]��3�q�ۃ��*�nv�V�f��\�v��c��%Kod��� )�c,NEV�h���h��2�᏶*	w1���u��\�L&zP�\ƈ��h�>YF&�mVe�M���j\�svɑ���V�㷋i��)gҘV�>�wIQn���=�b0�i�S- Sx�M�ɥ�0�ԉ�/R�֨dK���n�>�T�{R��v�[��Ͱm勾�vŖ�B����T�[�`�[��Q�$���EM��G�p:��J�%p�:���T��'+LǑRݫʀ��A���p\��pPK����6�B`R�Z�X(�cK�8�go�dnj۰���f���!cw�� ���Թ<ݲ��XF�P�2�)nS05B[q�ʊRd:Ǯ�����Xԭi��`�*vp�!e2�a�r�f�����B�k�ݽk$� �U�8%v���MQ���1�c��<��� 9�k�������e���9(#�4=��_��p�����ie��ڽ��;�+W:�eêm�rS�9`��GS+����޶�H*f7Ơ8Q���6#[i���4.�K�_W�]Ǆgܸ�14k��l��E]���N��-�Ui9��MM��૽���]� ыM�-f-αt(J�	ϛ���v�[���.\*J�e�h����Cj$�M�� H��!�L)j�u�Fw�Fm_N�(T���2Խ�7e���/�ۥ��Ӝm�B��q��6+���A�A�+n�b�j�e�
K�.f�}Σ|&	Ղ�3��Ќ�*EwAR��P��U�(��ѨJ��Vƛ�q,��(�+�K�ںҹ�Ż��`O���V������J���g�5��;Η���F�`50����f6U�t�]�<u�']�`]�]ef��<����+v3�FhO�ƞ�/̕vS�2��Ȋȹ^��0zvA:�P�M�2sLjT����kV�Ç�:��
}�H�⺭5�h࣡�S�ᑓ��j��o�����ݣ�m�D��	׻�ź�\�t�]lVH�'���.���֜��T��nWp��H��3+����\�	�cA��Ry�z/���2q����s���GH�\K�W���c2���,�|�Ǚ����Pծ��=�u��ÿ2i������1+�:�:��3i�j�|��@��j�r.�Ki�n�+R�b��X�X�I�ӹq�Gp��韥mwY�Ȣ��� n��F`:�KhM�EZ���3�
F|��TQ���J4%gT.�Q��4P�;;j�q�Y-TxM*�V���!�4%�m��wN[z�)��B�t�J�&on���5(��A�Ī7������z����䥯Qv� �Q6��e�7�v�A��Z)��ܮ��a$@	��Q��wV=�ͺʁ�,��M`ݸ�z�+o��hӃ�3s�V�" �L4�]a��&��>A�#��Mۋ�a���k���(Cu;owl6���	�J��
�V
2
˼xyT�9���o5	Ӧ���^��#Pm#�^F��v�Ř3@�`��|B���sX�C͏(Nl#��ҕ�evb7����C�6.��5�8�P)�۪R�$���Wp��1���Z Ud3{r�\����<֯-�U�R�7H[ƶ*��j�����;��I�Sy/Gc(Խ�UrZ�]���g �9D���ՙ��i���lg�L�ɬ�{u�`��j-=jwD�w,�2,@�W������D�$5��n[k"���2�n�;i�,];�DQYW�4U�|�()R
��p��wcy;�'Q��ΏN���i�%������0>��ע��y�N��q99��8��3�ޞv��xcְ��tq���cvz����-?�1��1�]6�SƁ��g5u�0�tB5�n)$Њ4�s���*+ڷ���m)[|��>v���ͳ�֢9ۉ����a�z����f����Q�4�i��Z�\�0!WG^Τ�jʄ�R��_D�J�[N#��
r��Yr��&��-�E�<��
Im*�����.'���L�-�M���/l7H��1m�4��1u����!7��=KT^-0P�\o;v�����	o��S�`R*��������77k��U#$\��I-N=Y�b�)4v����`�E���n�8LKABf>��힛}S�u���rʁD�`֎4��v��r��1�B�[;z�X�S�"�����Q��^PV�P��ZeMw[ <(���1�/����W3M5��g�ʜ���%�B�c�&t��ru�T|X��։ ���2���?ok,t��X���j1ʇ���GX�,��(�I-���E;� Їg-�5�gJ�Q�����[�����9Z4$A{r�����g�;R���l�����&���"�[�q ��gY���@R�(�&m�v�k<BT.��6t=t��[T�̤�~�q��^���+�,�Dͭ������У�����s=\q'B��ŕ�Wi�����k:�^�����ۃ#w6��B�wz\��a�w��}O���,H�˕j�A�w0�	Cz�B�-�z�Z�t�)="|�Sz��Y�ʏ:c�(֬���%��T�����l-����C
2�wt{7����6l�8����:e�tu����n�Th2��sA4Tˤy�I`:z�D��κ���ʘl��+��V��9$�5^˰��+M�A>�����P|��7��%����ʶ'o,����6F�.'Ô#}�*�tx��!d)�O5N�v4�˭Vţ��gma0f�i�bZ�k����F���k�R��
׵���>�_hC`o7M������P	:��Iܼ�IU�<ث ���34��)`����is1Z�F@l�|��I4����.�!اL"���lY�xbN�l
ԃs�Ҥw���2��]3t����%�0T��wS�G��e�	�1�C�8�=ϟK��DJ�0��CO2��R�<pe�k���:����2q4CeE���W1ܻ�̣jE�ĺm;O%�c�{|Q�\np�� ���І;AE#گX��|�����p͂�V-���Ҹ��g�!��1�f�֝�z���n<,����2���2ͬ��F�6f�x4��h�n��`�{��O�wۺ�.#%�l���oIK9#��CJ9n�9��:ȝo���M���v��w�W����4�l��=���ug,8�bKh
���z�,,���[k�F�j%�d�j�s�Ȗΰ���h�q�V�j]�_j��E�	֌�ξ{�����.؆7�+x���Nϕ�ﲲ�DD�cf�j��L�\��b�vV�n�k[b�Sn��(�rY���ݕCF�S��e*��d2��Ws�@v��l�FP�K���6��N{q���\]OzᥩՄE|�W_sھ��L�2ҋr��a�W���-���I^�JU�×�!ߵ��e��zc=NcJ|6fBn��؋�9����_q���8��MK����J]�yeg[$#�sw �uyawb�Z���E�%+x(�X{$әܽ����jғuE�}lv-T^fv��Pr��G�F��-Z"��Ύ���W}R�����z��eۨ$�K�0���hV�B�e��OE�ȶ��4��p�i�7k���lZ@��(���Z�kS�%Wl��TըB'�[������r+x����u]>7S]��Z�@�&�X����W�moT	��|h}���E�%�4�Δ�T�YB�1�*?b�U�V����z�ꕓ�,��[����(,�W��c�f�71����
�:�f�� �e#����M�2ʧS�Y�O+r�&�v�	/����`tvr�v�:M�x�0��t��L�W:�E�Nj֗-畘Q���!���Ed�9�Y�t2��'URj9�O��n�0��Eyw�������V��7�v�P�}��K&���e�j�]�.�#]\ ���(֦o:�����w7RTy��C%h}�e��gQ�{�!}$`ԩ;N����,��K��Tܫy1g:�oQv�"�µ�FP�u�l\��*�/y �T]O�^�6�'<���^�5��M��Wxqbe�meeq�C !k;�f�M�n�X��ڕy�:��8�
�]-�2�X�F�EJ�aL���#�Y�]��ܡ�7c;�M��{�C���%�ӣ����(.[P�R &J�\��f�u���A!�;k'=�h����bWVoQ�%.�$ޫ��5K�F�!��'�e��0Q����X�+&�L����|���'M��׻��,������5ۥ��M\�rs.6���������\Ň�6�����-6��{� -s�ñ�k��#��Ƈ&�3�A��}k4�t�WA9��̏)��N�}f�*��t+��He�P�d�yT}��1�S`NפL��S/�a}�_m5�,�y�(�:N�e�H�.��ʲ�\�*����YI��I ���U�pu��Z:��â�wX$��F�,t/sgdX�S�旎�˥�.��#�Vvv�m�n�EW<C���M
h��u��̏4w*���JG�7�ͪ�f���<ّ=�Y[�/y�[GC���]��ۡ�SK4q/x�c����3��h��cK��%�lm-Yeu1�*�El��{E."�/�X}0ۮ�Ռ^֋�v����ې&h۩���%뜟'ن���m����Wo?�q>b�[����C�*sT�xe�q}:˽@�l^@�m��f��ţ�H�����-ڥ�T�w�.�_�Y�l�<�ka᜹�@CT~�7���c�L_c�W���s��Fp���Kцس�9�IS;-7�:�K�ʼ�ZT0�7�P:���׷�]�S�Wq�zB�͏����-9�|Q�{SH��r#7n�YY�3'>�M���M�1�
�ed���M�gJS!K��51}����s�N).x���w��}���9�s)�H.��J>/4���\�*���(�S�t3�]6Ĺ]|�o�}`*�o�,Qg0ՙye�ѝ��2�`�"�Sp�ɮ��g۸
�VشWpk*Y	����X�2�1P�������2;D����	�  �x{������W�?�9� @^�G�~G�~��?a�?��~M�3w^߂q�G4O>�磞s�='�'��Oh�zI���Ӟ9�U�e]
�>c+�蝧�����2�9Z[ٰ�uZ6v��l8��Q����k�BV�a"�P;��X���
�Ϻ��%Y���s�P���X��ʗu8q5��
�ʻ�;];� ��j[�U��wPn�;�o\,�:��/�4ښ��E�M�9�{.������Ո�D��]h���Jݧ܅m�[̔�ڼW�
8a�&��,�0�9�ڧFA�e��K*���=��jz�v���Xm��G��lu!G�7�WW7$�q��"�'Ib2�h�����<$���\SnK�w��s�2���s��q{kS��^$o���'���V��XčV�z�ZtҮٺa�]�n��3E@�� +Ӈ��Ʈ�p�N��R�e�ީ��L�*>�z��� ^�վW��h�Wv��4%}kX�Q.�
na��s/j��g���on�cg���;۹{r��ݨj���Bs�����Ѐܩ�vo=4�;�D�V�ۉ�$gX8��ܰvLe�w�B����Z�v8r�(��5����3�tCgFz�JǽKc��oq��F����X�O��ˈn���f�k��K!p��M�A�A��!��r�Y��Z"=�J�ڻ/FԵ�;�SE^=Uc�?� q�ڎ��<�H�����j��vwA�Z�4�'Ye�ɰ��|�ձ:�4�z���LUt(�ѫ��Uu��Q���>���Һ2["���<x���z����{9���s��Niܧ�{'��x��ǝ��z�篱MRV_�U�R%$���J�EUy9R�j,�J����T��Z�*�EZZ�iZ%TJ��ʒ�R�u�V�T�$IRT�]D��R���ʊ���JZJV�Z��)ZJ���V�ҲU�I%�9%j�Q+KV�UM))*�U&�R���*����Q%R�U5JJ�V��Q)jE
���%%��KZ�-��UR*^j�U-U�ԕe}��J�*��V��*)*^\����ie+ESV��+���yvUT�y:)UT�ZR֕U�����kT�U%V�����ME��%Z�*��%V�T��V[�s�qW��Y*Z�&�"����9�"�䪥zo��A0}j���cqh�ѩ�%��s����Jĵ�N$��r��2L?�y7��Ic-�-
�T*%|� ��BDrD�^݃&��(f��'����7RJ���}I�ݎ�F���SȽ8�/Z�����\[�{������e��w¦��<�9l��s��r����Ć�ɘ�񾭞��썟j���,��yo/��ois`��ǧ��ǹ�,$����R�/�"�^��`�L��)��5��������Ʊ�����9=���ކ/��̺<�W�j�Gz:�a~��=��1�u.�y]�m��/PO�K|��k�Nn�j��oӲ����Yr�Ľ*ޭ�c07���;���s�x�������ўf�6�Hg��[ǹQ�L�����3��`��߳kZ3�6^��y�:A�9ޘ;�6�c3�ﱫ����y��=�V�"�&t����=v0��Q�$��9Α�[k?�Hi{V�ɷ��j�=�]=O�C���-�]��y��f�ݳ=����a�}��S�a��5��n���eu��7]s�U��R��f���PQ�n�h{/���3����[�����I^E��d�US��<1f�;����]�>�b�e����aٺ�溈��v`:�u8o��qo��pũ�f�sO��*����o��K�e[��j��/��7�fb�vޞȆ�� �ܘ�ޠ�#}�1������$Lt����g����:6�9ݏ�1�n&�k��G��"k�P�����:�<��f�������}��{�z�n�Ǡ��B���<��_�͖��Vi!��m�%fߦ��Ի8��g�f(�s�g����[xT��=Lx��%���f��$�ڦ�!㡌ǃ�3�>�5�~���򿻪.���䖞�	�6�ԧo�i��0o�<FK�{����u�{)8�sw���nQv�����_zG�Ի�&�s����1�͚���k�$Yp"��w�������U��ʾ�`��fN���5uC�dO�Б�0nU\�Yݞ9\)��Rq�i�鵾����NӶ����K��}�#���Zo�M���_-X�ez����!�ZM��jK�z�,<P�&Ls��)�CP@s��1֠\2��Cy��'r�c�d��:��r�o�%;�Ra��a�ʾĸ��e-�0�x�OL��]�B+�h=zw���1fV�yW����[�x1���M�Ǐ]F�����j�X��h��{���M��}����f���KU'������;K��,�e>�>���/���r����<��Z^���|zM�]��<��{ �0�V�۷G�Κ͞S�r�~>������R6x;�z�������Wя8��ߥ��nl�}O�r_y/X�qdL�}�Cr��Ұw����D1r�=�%���zx��l��~���nN�=u��O�5��ҏ����!�-]U�ħ�c���Ok[��~�Wt��ʆr�_��o��j����UԵ��\��1��R���Q�u�L���s��O>�˃���������g�T6��5��*Fc�$OS�|mW3�_��o_����u����+������$;�:_f@�E��:k �R���yU�O?�;qw�o�T�w[@��OB��(�����W3m�K]�Ӹ�Dm��/�;��]�G3f=�n�7a4M|o��s3�_[���­+���/^��En��v[s[O�C�{�[[!�V��͚�:�]�k����]�?�j����w��yf�3Y�h�Ň�㐁��|���T�eq��)gվ���0=�Z��Y��K���#=5+ʮ����rN��|#�we������E���)�M��{U	+�l���m,u{�9�k�s]=�gbl�jsޝ��:�k����W���銿|��c�7;<��م]�W�����2@}�^��߼�g��yÖ�e�z��ek��eOC����4�k���5Ȃ���OPn�M����f�������_��Cj�f���r�[3�=��0�<̦�Y�����G���=tR�}�}Y����{�K�.O�N���w��,���u~s>�v[$�Ƃk�q���'f{-�O��w�}�=:[��S@Dy<���L5E�	w�rh���VW.s;�������"��S���8�⩧��n������s�B/e�ss=t��r/(=V{E����C��ա���_�\ ��*�NW�z��9)n�]u;�*�6�׬�mG.��(8��K:Y2]�3�6�T�7G�s���7WX3����GK3k��ڮF��x�r΋]�ޠ��é���Ђ�݋���tY�c���j�g����i�d���u]N���E�lre�(����X~����ikۑ<�ƝEbD^4�N�@��I5�����6�e޿}Q씼)g��ݮ�u�m�x����	W�U�����/�>C��lg*�wB�����@�?��_�+S����U��^<&y�������� ���C��gZ�24�26�����G��30��y;����N�ǽjz��u��n�{���X��pQ׶��6"z�CL	��^^ں����ɩ�;��go�/��u��rr�⍙���)��ڒ]V�Uj��V3�I�썟j�=^{�w���{5�nC��j%�ϖ�r.s2z��J��9\�E�xEWԯ��uL�r����I�����z��λ'�~��zs����Ii���`�$���N���`? $�6�y��g�����w��_���z�ӳ]󖫚 5��[^�e#Q�<B�`����ǘ��_"\f�7��
��49o`�6kk���8U��#�ƌI�FusD���S�	������b�����!�+s���\v��rD�[�Xv.��45�mY��5�1��s�R�c��EeВĹO�N�����x=�j宫���HG�uy<o�d�aݑ���28@m��~�<"G��J�s}�l�`����k�qyl�[:Y�s��='�7��`ļ9��۷�q�ͽ�;�Cp�����&&�1�}�HWz��Y�9�u�\�37��&+Fz�GeQb�p�㶗�<��������o+���o��Υ���$�~��,�p��O�
�σ���U�������~�����NS�w|u���aN~��ތ���sḩ�iW�|WC^��D��;��{�1X=������<�zĹ�>.����5+�b��c�#*
G2'X4�͈B2����nby��Z�A��F��=�`�S��*ozw��2g9N\��|7s�*��rր�J�z�����U�_=�O�/h=Q�Q�TH��,v^2<�0���Zr�ɍ�2������	�i^�Z����7���i�Z\�uox>�Fax�Yh��{��e>)� �&Eܡ��ڛ���2�9����^�}�Lr��)�e�: �Uȥ��\l��Eɪ�ц��N3Lw��5��y6MAg>��:��M��	��Ko�U��7Z����]�Q�җ{"|�[�u�����������m�� ���Cz�(7����P;a����b)�E)W�}���o�� ��#L��0��99$��q̉�j[:Z�j]�ati\�r��u��^	ꞣ]�/��o�]�o���׾ĪN��oo���B����u�=���g��e%��\�l��sƀc&���Mz={��oq�e��^��f�D;��@��y�<�_�m�_�Z���2���Ƙ�Yf�{,�~�$gw�/?wY�L�e?��p���Tw={�T��7\�b��M���ꮾ�{s�!���S(U�({UQ���,�[z��֯��)wc��z|g=�w���za��b�?c��Z.����4=e�7���6\�7մ{fH&=�=ѷ�Ò8����
�f<���S�~��P�c�C.̾6��N2�z{�4ѧ�b�@m�Xt蝾F#�U�c��+�W�46X��-���%F��e[�l��/�+�B�yL6+�Ra����Įi�9G����X\��(�گ��P%oDr��Mh�ukt��g�e���ր����fs�R>�����K\u�W{%|�4�����my�7���O���<���O@�1Z�z�OFb��+�/}F��4f���Oeutis}+_ç�u:����dr���K�=�A/�Y���9O w,:���e��K;���{�Z껏 [U�̘�$�F���P;,�=�LgFx�|,��Q�Dܺ����E�N�n�Sy"ٽ�P�����{t_j�}D����P@w�[^[)�j�7��|�Igwf�zm�趢�u������X��E<ɕ�{P�ҞUz�xo����֪�c3�zgZ�fl��y�d�x��Wʡ��棯(���H��9#�Jn����(��EܛP߼���Q������0�A$���<o"E�M�;��;.W�R�J4߼�;����_�Z^��u'NsYs3y����{��L_��O]y�M��Ѝ��uu׈y`QrݕD����,OY��FJ}������8�5j�&���8վ�ƥ�o���T ��s�dٽ0�d(Q8��&�>w�TT��j��]f�ؚ��W�ƥ�!Hޛ�ޓ���>αz���5_*���Wi�Ü�AT(VW3��|����}~���U���xC`��h�U~qc�3�0��5�&ץ����~�V�����~�ߐ��*�QO�]���{ދ�(z�U�k����%G��i�C���:��es�a�>�o	y���q�SE+��k��E��oֳȹt��z.{^P�_���J�og���}s���t_�IDz�/]Z���L��T3�ӋG^�O�Ϟ�u'��vw��~"6nK�s:0Ì�}}0Uk�K��ܠ'���K]i���=Ϝ��$ǫ�j����!AʇC_�e�O%��V�ɻ�M��>����k2O5&��26���5X��Z{fw��=������^���t�n���+�TU^��{a�aj�����{sI}�< �L�ܒ���W�&��q��ޯ���w���
��>���+_#�;voc�PK0�-�݅��W���\s(�,�1!S<U{Um�c�묾͆��C�$�fr�Q���QGԳp/gg*��H!FU�J#X�@�RķU֎W�1�+,����:�U��K�w�r���O9S��Mr
��`��x�J5ˢ�i��rZ����U@bj@s-S�Z&��ɻGe'���S}�<�o��V�ۦ=[�7Sp����RO���xG:�w�WO��y�|��fS�O.��^N����VZ��\}"rz��UG�GK��:���O*�m���Zk��w���ؿi��==�d֛�����[@��^T�e�w|�x����gA�M�CH�����׀aݐI�c _W1��e�7��Y�U������=I*�T���}�a����y�1k�S ���=.���P}�x5W���,�'e-��}�~���ػ��qau��4��/I�վ���2��z�|0h�@��1�ͪ4��Í<r�ێsK޾��w��'�_��ph�|�YA�aze����1Yt�l�Q��"����~�}�����'3�3-ͣ1��42�QWF����`8����T�q���Z���3@}aъ�̛7�įo�jtZ�ڷ�o*J�+Y�Ume&n��G��&�k��1�	vB��f�ա;��lζ�)O���k�w

�ymd$��y���K5�2Pg�Wv����2�|�U{�n�٭��~����� !���/��e�u���P�rn\6����7A����';��m�4��(Y�R#d�i[h,�m�Iۦ�H��֭��:2�;
���fT�_.a�\��J�fd}7o(��<wl�а$p�94� ��m�`��:���k�� }�&���QO7����z;CXt�xT�&'�j֌1s�gs|7]k���7��^��*�K�$nw�f��{��y�����-��U���2�.�4F��v�:݌h�ں��2ھh��g4�B��Y��˝SF���)[Y�!\Xξ�֏�X��[�y�v��<G(�@t��T���;�ݺ����<Q�M�C妚�(��s�S�S	M�deH�C�=����I+�/*c]ֺoUų5��*Y���)���'3o��´��
����X�d�}���<�d�1����iKN���	���k$�պY/D��&��c�1̂d��ڜx�wPn̤��l��;���Ŵ[al�km�;g'w�l[J�G}�!
����a�q�@���2�Ir�î�5Ϸ��09��{]��n4�B�6����n�<Ѕ֒�@�����ĸ�U�5��ؙ8I���)r3�f#���ȇq��嬲�V������Y�iaW�zyd��d
��MG�}vX44��+�r����3��>�s���ڗ�.�n��o;˜P���``g�V�mrkE�B���k{q����.:�; Χ-|0���;��jR��D�W]ew"������*:޽��қfv�TD�o<��`�D�h��5���&�7�N�愵[*7[��v��d��zQB�h6 F}�G�ꕨx��.�&���n��f'�X]��,��&B'١���l,�q�V��ɭKlJ=&j�4ݔ���ʚ+B{�wfݽ��q(��n��(g��R�n<2�:<&��S4鏺K�o
�`�.���6YY�"��ۏtE�X[*��8�^*��d�^6m�a�3�M�G���5��ʏF���K��E�|_[���:�z�������T�E2�K�I�i��W���������fi �=Nq�Z���q�h��R����
����Kt&$w��Ǝ�z���j�J�t�Qȣ,b�To9�)^������޺���d�U����C�W�͑��AK3o7�G:n�d_BQwc��;��>�W��%E	�|�8ܛ�m�]}cl���K�Rc�[�s�k�"ݳ<exq]��ѥS��k�쇥;�+C�j����Y<Q�h �.+�1�.��S!ns�H�٩�엷
i+L�aj��e�r�'�׸;�\v�wu��7�ER�V��TK)$�RH��ZR�E�RҵUD�K%R�%��MJ���h�VU��ʓ�g*��ҫJ�V�++Z�T��jM)R�%�e*��;RJ�Z�IV�Jy��ߜ�T�J�I-ZԒڊ���i*�ʊ�eTIE*MJ�Z���J%T�+$�^s�ie�"�*�]�UR�*EH�yu�����R���R�R�55�Y-J)��ΩiZJ(�%����5%RV���U=s�^�ʵd��I)%jU��U5tw]Z�Z�7-KT��|]���U���=N�VR�2�R�Z��s�κ�V�N��֫Z֊�ʼ�Z�[)IR��P�%-i$Y]�*H��J��,��imT��Z���(���Wp��ՒD�'yΊ�Բ�}�֑Z���Z��R�|����$_%�����iK��`{�ՀX��׃�l�gTvq��$��ͺ���;P��W��;�ff:u��Ӈwg���,t̜�27�s#[���Q�Ǟ�����J7������`(&��{_�)��z���W���ho��4ZĸߔV;6l��o�%t�(	���	$����ӧ�}�������ʗ�׷��,$��r����Ş���M���̾�G���`�>�G����R�4�<߶��jq0�oԱq��Jk�d}�j�ק�}q>#hnk݊8��Eʉl�/Q��N,;����̝S�?��a!l_�3I��Ї�yu�.�4�eԂ�@���^�*Ʌ~船�Z�ْ�VwU�<�_�W�i�ns'+��{�(> �ل�} ����ԇ���VF�Vq�]X�6�8�Z��WR�覻U�k^@�x��׽�r��]�sVM�n�竴��߇��7���uz7��� v*������J���(��qu�YV�Z���|��?L"#s
=��������}�}>a��fO3O����}ݩ\5�\"���|&��!�����wɽek�Ee��=L׈bU��hV���`����<��9�R���ʥ���.�p7���>�a{�|���?)R]WVu��oj��pS�+��Z�<���y�r�08w.�e����&�'_�v>�;�����${}k�غ�9���"��0�;�m��l7ڸ�S2_]i57��H`K7e'K^ ��Ntd���l�cu���{#�J����ɷ���Ψ뻬w�� sM؞�Au�={���WPƞ���>0������/5�qˑ<���S=	��w��]�vu�-� ot�8�OO1�x�h�{U�Jʠ<X���Xq�	S��o�vH���}��=�����m��hOB�Ϯ*�z�^�ƈ�>�C3>�@]Pw{C)ͪM嗯r����W��c�}.�Efŧ��uy�?8�ȶ�"*�碣:j�A��+�l�7ΐjs��nM��;�.��[���%@��i�yc�1��zg�e3e�v)�������"{�Wƭ0���
�'kV��=������w�n�]�Ec����d�ۛ0�	�o���%�zvA���>;�8K�YT���t����&���VX_s���mV<D�xZY���a�ه��U�&qd�f���f����@Fm�W�<ڢa�]����SԽc����s�=d�U�]R�M����w�<7�>���v��C�t$dK����xkP���@�d',D*���W9FwV�< ?i��Q��e�0��g�{��1�1E����9V0����!�^�2͈�|ō��F��#�R������T٫p%X����+h���MV{��=�K�7@����n�3�U]�~"R�Q�g��]�q���s��]8jca���YR��Sn�7⺰��:���:E�kЉ��9�*��C�`�����]IO
5�|����K�^.Y����ʝn���E��L��QE��ܡz��8��8��	2k�,;s�����۾�Na�#�F<~��0y�(�-ퟅa�_F�-������)�>ͩ�¼S�nwd�!��i��mJ˝vm��� @�Z�������_H&F��e������aǇR��=���E1��U�_�磨��N�uǆB�7x�?q�}C���-yyy�~���󈇷o'f�0����(k�g���Y{lN���]�A�iIO�E�]�ëݳ��̎e����-6�K�g<������6��XH�dJ�!�RU�Ո�HY-�{�8�F����nz:p_ME��F�;	j��������83
�.0�]N����%��ZS�ơp���jߥG1��qWu��1�7���db��P�&]�k�������J��I{���SYb[����*��^�ܾ��P�p��c�b�ȃ�!@8��_�B��K=�i֚�o����OtW����ju��ز�?��x�v�@'9"qR}"'�ɾPKXE���:z�%K�=�>5����3n��m�Nǁ~k;b��C���&�#9ܚ)LKRrd�t�ߝo<'��!	��)p���5u�$f��	^�j���/8��͘�e_.MI_v	N����mp}}Om�L��dΠk��R�]MFl7���c}�|�l�|bs?XzF�%�
'��>�|PV.Ϣ=��dDʜ..�U�M4���FE�ӷ��?���&�:��斯.�>0(7A��E5Cf'B"NG�g�aĿUVb.К��y
�g��W��u�P����Ü0r�|dM�G�p��ޤAo�fN���Co�+wsri��aD|%u�Y�ʦ�i�L��CuFΰ��)�l�t+sn�s�Ɓ3�V�g ���c�ޕ	��+2��-�BEz�r&��ŬwJ�k%K'�TגJͨ���fKM˪��0���X5t*�����[㾧�B�D�v�Sh�r8v�񑑂�4�.&����W��b��|Cڙӹ`>���t���<�VEs����I�`J�gzQʘ	�?
��[���(�:oN+��A�Q/~s�0��SwbUm�I��1P�lr3&#�gv���PJ��<U��f��ۚ49l[�O�܇�wi�/Ɣ���)?5�n*�7yT��>�j����8���܆3*>r"#V��qm�.{C{���T�v/��W�H�r&��A�C���NM������F��o��{,jf-;w}ԙܳX�>K/CMmF�㔱wYRN�ą���%�R��X��xʭu��C���d��3@���ݕȸs��;��Y�q;b1k"���m&j��@�zh'/w��K�}������99)�Ͼ���S.q������pb(3�pa��_�!6���l�����JKZq���f0k�^�7������CsfةG5sp(	݀��jfĩ8g'6�|&_ub$���W'�+n�i֯>]<U�9 1��5�.Q������聆ސ�'��%۟������꼎[q�@�K��1�(ޥ��{��A���@�W��Ʌ�A8�"	����)���K�>�����ӵP k���P���r`[-t� �P�B�J�*�6Ӭ�Q\�:��{4n2xZ���f��-�Y'$���f������D��T�p���U���o�ݝ�v�f0�gI�OT���ġ�&�%?�ߍ�X=���3$BV�n��ׇQ�tJ>x��ۋ�W(��{D]4F��P��~�[��CݑIYj������u�٬jnjS^�[y��ou�G�/�k~+8�s�⡼�r��l�yQ5R^�P����"��
��5��76��*��8�k�ś^�P(j�Z�vd�=j%�e��M�
�ֻ�a�^�u4����1���|J�h�S�$<�U�Sɘc���'a���֚ev.ES
z��}xN���ާr쨟ѝ.Y���il�7��Ya�_+w[��e9��;oq;�i3�u��h���и��۔���+P:�y9:[	�Z��%.�C��ӧ�_W�P=�UOH�B��wj��4ޙ�:$����s樤�kdSm ��=�S���3a����Q3��R\���T���.��'�����q�Z�/��]�ǚ޷�=���)����'��Š_�Z	�dϼ~��L<���
dO�����k'�&6���#u����S�׎��s½��V�:r�����{ܹ�k)��n�{F"��U}+��>PY���(���Rbj�e[}�1B\+}�Υs����l+>��~`�J��0�y#�J��k{H�q��,:a��۾��2ҧ�.܉d���C���5����}��JV�1$w~����:~.v{��*�Zhh���C��or�{�F���L��U&~;<О��y��̓iz��������b�uv�������:Z�Wbf��j���4:�bgS�(ȶ��B6���z*0j"-��ߧ��E;�����K	�Z�3�}:h		����~��c�_љ#h0iށ2X`s=�:����ݛne�ޠ�(LZ��JX�(|�`FG�W�<�	�ٹ��ޜKH�qs���$�*8O_[��)�]��"��4$�l�r�I��}I��®�эwR84�&�2�؉�[>�u�%7�N`���uV�.�cS���]!��:TD�K�e���J|Kqd��:ۇ��ւ�����Q��TUk�9��Gfo��A����0�����zVY�,#_ �B	�Y�O��ޝ'�ՍR�uqHW�"e��x�W�X��Z�G��H��v(�;��6�kZ/����<52mO��i3�Ԋ���l|q��!N���Q����3z�KZ����2���5m�fa����P�m#"[+S���~���G���/k��rB�Qx�99��e㐕脮]<z�h�/���c�L
���;�Y�udQ�w1U\��zWr�m19��V���F7I[����%*���Hu8w�6%�;ɗ�qE'�r��p�I�%�=e����3ku��Ɇ^C��ލ6Ӎ^�)�M�'.�A㫣O�t�mZ\�l{��F̘^��V/^�켥�݅mt����$z��Z���ˑ���} ��NsI��Cv�R�̋��5��O�<]g�E2���ԍ��59��~l�����t�U|%p;��C�p��o:�r��g����x��Yafa1On�Ru��9���hS�:���V��gw�Fe�~e�mŞ�nŭ�㘗��범P���q Q�Z���������0�,��|j�v�k]P6�'.��-b��H��!f#��u����x+W��U��7Q�?�vMa[嘼d�ڷ^���F�Tb;��0���E���i&.�tk{e$o�@yp[��u�9i�+Cj�
�m����]MG��]ܵC��7U��˚�e�J&V�F���y���|n����=-�{�f^[2p)KR���YT�s�P���2���b�A�G%r�,�=��o�cA�^�OU�N�;���<�&5{e@ϋ ��5D,k��.}}]e�`�T2�Sϐ�ycI4��Tm���0c�ɓe��}�Ӓ%(�z�C"D��C��^,���u��Z�v2�N?ki���k�-Q�o^F�����<�D��9�D#��3�|�������X��䕾��Q.���qU�J a����K�f ���\�:��f��Ց��"4^�7��z�����˛k؎!w=
��sK�i�o�
�d|�h���X�N�a��42�v�"��ln��B��`�Q9]���7���7�ZGd2�Tr��"n�դ�<{!mT0�-��i4FBG��M���]�2���)����*�ֱ�	-�Rk��u�J��2{.��,���Q��4��}�O<����Er�]��<O�ܿ<7'��R��+KP�2������#V��k�@��~��m�|"=�|�����<ʹ���1''\�=,�Ҭǀ�hhҬ�����Y��Ք����3*j�X�h�o�ĥ�`�J��-�G%�;zoIC��t3:;f��S�C�U�r��뾷�i�N����ř�5�c5ܫ[BRFe1̃-o�?�2����i��ɫ�,:��}����f51�ٺ�~������Y�E�!�^5�Ì�e��e�R3m�.�ȑ�=�֓����dgT�t�62E��es���]WӨac��SQt8�~�!-�z�-�i����������v��G­���2�V��w�;��EAz-�N�,G9GM	�v��f ��!N�S�=�E:�*s��kN�9�XUhC&m UsT2��}�g���g^z�H3�_� ��zT6�P�{u\���	�C��O~u��4wB"��ܨ��Ob��-��nEB����܋+�|��c�0I]�t�{�g7¦NN[�>=�̿�M�}������U��B��ytKc�3lT����'6B����vBo+�S6�Xњ���D���wY���FR�@ʒs���� ���R�V�2]�D=�-�
~9��+�>��Ϗ�ϲ�3�i=T��`ٟ5~z~�*�_H�3��r��3k�������XM�#�yf˓w|"<ָ!�����1����`��Y!�c}
m*RT��s�"Y�
��s7w�ؚ;L����,_��/����@�Q��2E�'}��r��<("ֵ	L��By��ٰ�=X�R��[@�[�\���.����D�w��؎3�zU����sr�c�Zy��Z�Nݭ���%XPU.�:��^v������ʔ�q$䜻S�
�h��:3�ƒ�@�#N&xtk=QE��磌F1�&�r�m��ڎ[r�u�mF����_	 �I?@'�C��ιL����T����5���t?�C<Po�ߊg�++���ɘi��q�iM'A:k^ ��P뻬~V�a�Di���!O�ޤ֙K<	ח��"����U^�cL�1�1�|���8v��m.՚�޸:������Lf��������ɞ$f>��:�TóC�N�{�gD�f���v���<~����Q��]-"�K&6
ʦ�+��|ٞ��<4ۆ��5۴��ݍ�</�f��t�BP��wk��sG�U����1I�|�Si�l	m���{��*��^��4����fc�ϠX��{o_���J��*V!q��ն�H�N!��Z�5��Eia��"�&�v2�wt�am����Z��@����^C�۪��U�:0E���Qkw�w)�Y�g4�9scx������8�έ,�֨�h���!���xz��:o�3��(�{�!�5�{�c/�83�d��T�ʡW�glW�c8��ڤ�J
�0�y#���ް�v~�KnVtp�{H=��E5�F��C0�7�����;*��)#��4ZAx x �4
}�3���Ӕ�+���Z�r�mN�Х��p����"ZIդ{m�f����em)b膎N�*�j�+2���M�z�M��T�������lfJw��Ɋ5֎ .c��q^c{���؆����Z����t�P]\����5����Zd܊˒�ޅ�=��f����j�ˉP Z$�9�b]���<x䗜@�jcֺ��8��8:�c^�e��e��##p�wN+�����-K�ty����p����V�-8��]z�����^S�2}���t���UWm.Cv��C^*|�����y�N��J�G[�=mެ�s	�5܆CՔ�j��i�K��0����>��K��56r<1]t��V��ъ����9��Ɲ��/�1J�&[�r�2.�5AR-Q�07S���ut(fi�7R5��.��{�8�\xںq~!g9��ς�,���4�<�����3!��]x  `-fV�Sv��Uu��'=k%��kl�mc��Ϥ+:*��v�<� �����Cu������΢�瑶k���YZn��N(�UeH�[���I�)���)%�.Z8����^l'���ӥ�P�&c��y���$+���m�J5g���������k0u�@j�����wr����H�̍*�A�S��� �Ks�l�6�КK�]/��%3i�H��+�'*�bաjƢ��g�~O�����T(v��"L�0-����ޠ�4��ڊ�Z^84�W�T�js��:���V��ć!Ҡ�sQv�t���*@:��1\(�KR�T�v����W�qL��֩}��Z�6�T}|Ɗ�}�������I(��r��g^��j�Ӊ۬9"�65n]�c-q�M�kw�-d{��뗚���3��av�r�kkGU�E�r���ʍ;� ٍ�+3���."�N.�����*":�a嬣���qu/b�Cw��#�j���ҍ�ڝ�w�` B.���>��wYz���+��� Xj;=RrcٲVk�%�s�]��{Z�𱢚��mܥ�tD\������9�.�*-}!�L!����Y�p�瓡˕c����rc��srR�O+zN�n�n�%�N��7t�#��k�/��%�q休gL}B�˭Q>�u]�Y��t���V��)��i+�k���J�q)��8iS�� �tp����#��AJ��0�T�o"p�pwY��k�Uv2�_^X�5xn��N��H�s�b�gh�o1�H��ή�&u�s��'3c��g��B�&������Q9T�Ĺ�Jq��T7����r�R�;�2Y���n����m��gCx�C��Ѵ-E%��,ZTI7���TrJw5�l��J������4�:�F�y0��Ӗ�E�k� /�����!K�[��A	1�;�����z6(���#�
��<�#7���X�* ��*�ȍ�\��C;8����цql*��No��d���ҏ��M������pN�����)����4-�S�m])j�݋�蓷����4h���S�b�R��K)��V���*��iUI����UV�ZZ�i+�U�UP��[S��ER�T��c���'��EUd���n��η��jJ��QV�<��Ǭ��g�x��t�V�F��^\�jռ��mZ�Z�O.�����W��Ej�.�-o]�,��nIZ�t�E���N����VWGUJS�Ҫj�R�Z�t��$���6���=�)V�|w>g���|��v�)�):�V�Z�D�+Q�y���u��u�.�םZ���5j�nY]l�<����|O/4I�+Y,V�%t�ܻ����.�\�rղ��y��VՕ�>-�R��Չ{�j
�ݕiZ���!���u�=���룮�jNݝd�yxV��J��en�jV��SI����ڳ��<����Jgz��ެ�Uwn�j׮�՝y+)]w�n�e54���{�����s˭�J��QAT�#�E������+Vޮ����os�g��{3}����}���1雽���N�򇯊j�N�9�t!��v�֒<�	iG��Fu'�C��Fp�JVP�ɽ"eM׊�����Ϥ��D� ��~ ����lͱ-�#s�����\*H ��Pb�5&u~��xw:dc��S��S�Zh_A�_N�qn���{�DS��p%�<]�퇄�z<P,�4�.;P��GOa��N7 (����[�#�깱��i(�{�]�?��A��	PH���ҝ�����n?4`�����w�z�H�y���M�X���}�j�֘Jި|�b2=���銡�͌g�k�{������z�J����%�M�M�4s��K��5CT��J�zx1�a�z<u�����J�Ѩ"a�̈���v�{�MCbtC��dگ��&~��EK��OW�d)�!{�z�ml��
��X�;����ս��܅�^�@ft�p�r~
�7,��}?k�$�Kڄ���P�s�4��������ᩈG�����'�{��Uk e�P���)��)\�]R��M��P#7�udQ��	F%K��kٺ\�t�s��7%?/�'�S�iOՙH�j�|w�=��KW�'Gu�c�M=[��{�ub�;�5���iچ/!��{o_��N5	r���ܳG��k~�%�&%�#o"�SD����튇�}�ګ6���M�;�ۭ�����1Z���pw�n�F��2��e��w��g�H�!;�V���hᏤFpE��\ͣ�>��Ҝ���iui�ŐB��*��k9.���7�ʔ���m�V�w���!�#m��ͱ�< �ؕ}�ZA�V���)���y��T��C5�nV}ke]ȑ�Z�r�h ��<�wU��4t��p����8�u=��IՏ2�e����4��g���#N�R��,����n�\�=jvq��n�/)�����I���9�S.�r�,<o�B��1���<�-5��N�k�]ӫ����B`s��<�;uE��O8�6��ZFK#�����ϭz��n
���4�������E0��+_�!Bc/���6.�*���Ǵ���7U����F�J���~����y�ct\�TDr��ZA%���3�ح�eQ�[�8�+e*=s�w])�3zb�kw��Cz<E� �拃2��7��r�ȃ�!@8��G!�"��M�����O���>�nk��CVL��Aқ.,r�k��\юfc��Cq^�H�^O�D�;7�Vm.���zߎ{:���ui�	��x���$;
�= �z�0-�|U�j.Zs�>�؏nKTf=e�N���nu!�d��E�mC�̅�C�
w/a�J�nE�)�(�2k�z*�:��^>�@f���P�ZeK�ua����qt�s�O�ݮʏU#G�����kL?s:�p�u���kaP��aK��p}��c�v4g���=[y��p�b��F��[zΑ�t�f���0�5��%��{��wѾ�+(:�KNS��V�\v&Ev濏ō�5�ic�cic$m�m��2[0� ��e,BNT����-�Aa>��
Qg"��ηX�mj�%��d��%��Z�?)1�{E�_+�<�%t�$�3]C����_�t�pk翤�����^!	���E�0r�Fֺ����ʌh���:xv��ٰ�����}pHq<˃�n}��&�d��x�ݺԅ���\Ļ�q,r��I����yB�d�-w�r��a�a&�Z��/Vi��plMS�z$�͗��HX.�26�z�
�1	��*����]6�V���
rr�F)���Gzޣ��X/��R�B'|kys�@Z�c��ATk���tKL�7R��%V�r?T��2�XV���4�6+1Okq��2[�p���8�����B��i�����7O�cTsv2Ø:8�����=��W���҅���KB>�(��>��q,g݊��>8LP�Ury�`�A����Ôr��J�~�B硦-���jJ�$��1�G��o�d��2��75�|��5<;�'`��T�^�V��N����qxf��`�*l7HyB8��4s��F�\I�m��}��6+���� C�?V������N�0�}����{�S�*Ǽ	�+>�֔�W|^��h,�W4��ݙ+v���t�O�=�d�6\8��ܓs�tY̹@v��-�z����h-`TYǝF�CQ�uq��ي�]�uZ����>|��z߉�ߊd���6���Ͷ$12[m��D�%����|�}�>��KT.no�N���Ȫ-�5Ig����C�38hw�{�O$,�ސ��&L3u���w���<�)�GSj��vF>�̪���`>�E�.�B��#O�!�0#�w�볶ڮ&lew7��F�;�����^'ɾ�ˤY|�.S��7Ц�����h�&�_'��Y6�"�G0�|�q�˹�BP�q^������h����P�^V+z�Ջ�h�����P���b
�����	c(�
�Cb�~3��C˖}����7��m� �(�N��ܶ"'2��(oJ#�	�JkF�K(�~W�z៓�ʹ�d�-�G���;׹Q&`�>˭ahF��=�<O���^�W4�c�"@yQ5R^�P������wA�"e�cƫ��Y���m!LuT�O VU���Z�vd�-D�l�Vݷ`W:��#Рߐ:���t�����/g��zFTD�'��@���P�j��[�M=V1�5ֶE6ג�ǽ��%GL]��I*5�[e0B=ྡ���}<��q���t���/
{�����wR�]y��o���=�&�FT>���l���ݏ�>W��G��Gھ��sP
�O�t!cw{�=g��,�{�|�>M���:�m���]��8�.��չ3r��l7�R̝�u҅UҦ�Y��oF���*�,X�o���L��L�M�,ZCilm��m&٢ٴ�I��������=� ��Ɉͳ�L�a��հ�J�-�?�u�1����.��BY R��~����W��{�.J�����0�"���q�K�W#�܇n!��ht�A�t��PY�dc��n%�8v/GD��Rk��v���{f0�7���Ru% �a��H��.�t���+���[W�����]��L�ż���Py��&��o�K����,h�|�lZH��`$VV���B�	��b��y�xC�=K�:/t�� t�w�U&kg�е��8�����[?��wl3��b�gγ;l3��F���\3ƥ��2�:x��x�.9�Vu5���Fi������Q�<ذc�H�� #�f�M��Bv���׻x� ��}5��m��ӽ��)W]��I�tL��>�'��H���d�Z��Q����N7N�<�}rM��fQ�X�Vԗ���:�L޿���e��K:	�o����tx��R�u(�U�.p�~�cz��S���l����v����ț��A�.�k���&[�"����{?���3��"a�Wk,�ָ�H�R�f�.iʔ�*)(���S�j�~�qe�6 �
�߯����67�oIWJ�lᗐU�[��q��]���&X�MҦ���E��쩛v�{j���彑���U�^W>;��jNnnP���}_}�}�Fl��2Fa�����ǟ?zj�">��熜qM��#��3G�B���B�������Q�w�bx��j�e��E�O���Ѧ�j�e������<�/W���^qMg��
��ݭ��|"2��ʩ���sKX[q�xt1\���YWP��>�)T��꺜:�C>87�2��f�ri8��F2n�Q�ܨ7o�,�{`#Y�.�mC	��mT�m�m� ��f�S�Z��g.ֳ�O�ם��wǙx���	O�m�נ���,���X��h��^C�y{��l�'��b/WZ�v�a�K�3J=$���I� �)�?`*}�Hݍ��|��?6S�x�c��Tx�nU�Aj�a���#ώjbW�U�jzڐ���EoT��_�Բ��؝;_s�hW�cJJ��4`��ǵQ��c�����R�o�B��w��j��o"��q^�j�����G��x���7��[��y���<U���PHkؘ�~j����۟sxgJ�.1{Rj[���Pq�x�ٮ�3�ơ��s��b�j�ȃ�!@�i���j��ƻ¢�����Ӥ�w�m����"�9%����	q��<��R�I�����F�ӣ��lh[�a�M�[[�V���4ѫ���9�pC�XUjb�y��vأ��Г:.r��<F��Z|��f�l�WOb�Kh.�}�6(W(����6�t����j�:՝�7/w����߿Z�z�����}ߖf��M�i�xx ����ᓏ\w�(���/�2_!c��.���TW,�Aޕ �;��ȟ@}k�Ӓ�{��q�p�(uom�܇)ӄ>բ�w���yp��y�����V<�9�D#����V������\_S��T��&D�㳗��R�n�z�T;�x���g�A��lIX��C����w���������dDʒ�PY(���m{j�ҍܞir�'��T4Ssd3��t�N�Y�2<<������k�������^�t�o����&�97F��=�j��A�*E��.���ŕz,oUn���1�vդ�~�DƘF�Plj���'X�Gc��ߤO����3�o7��O��ɇ�!�ީ�c�_<�P��V|��|j�+��s,r��l�ٚ��J���z��/�p�l�)�ư��O�1M2�k�@��~��@��u�_�ԥEڗ��=����ئ�7��N훷}^�4egE{����L��e�u��?G���Ȯ�~1�gi�ڎ����%�*]��0w=ta�B9S���-2=�n���n�v���- St��+VG��QU�`*OӤ���4e��3�ҡc�*Zs5��Է�Y�����a܇�o�m�B,Rbt��|e�ǐ_*3������ͦ;d��ʨ��~�^�J�н�&ݮ-<Gm�`�+����LWV.��h���c;9bPue�WMl��7r��5ɒ�;���"�����L��P4��K� :5y�jҬT�/�N-�|��#��kT��&�/��M�q~4����)?2:�k�j�q~�\^�Κ�Pֽ}+��j���8
��DCXhN�Ŵ.$�������y%i�*�]��s.�-�ok�W�)��Yӭ>�� [����$�d��C��"�D3�1.��{ޝ�x_DDNl��l{77%ٳ���p-8��ӯ"��xjQ��`�?��!��H�Yi7����p���k���&�u�+���ӭe��J����j~{U����{�(�db��sf}��W�B��NFj�(�_����9W&SU.gx�=�D��2�h55��r���0v��m��ͅ�7=8�� Y���
_+&�gێ���:��K�u��#C��㫇��8�em��ؘw��� {�Q�W2T|�3&C��{�]�o�2�;�r�e�^W7�}�͙�/%�gL��fыb�<bG���}�*ޤ�}�TF�ڇ�a�Mޚ�cw�����L�K�j.��|E���h��i��x��J#�~�vh*R����J��
l!G�Z�fs�PM,��T�Gʺ�ot\x�-�8y'q���AfN̵����)�5rYs�:��މ�_^�����Q����1}%a=7d�b%5�mu|>��}]�s�Hl�Bgv�
u�b�[{+`��쨞��݈/1��G:�^U�6��m��}ݼ��L�n���E_����x{���8M�I�d�����������Z���澮�'T�9d��Q'�1�"$���.�_=�����捕2��{��!J�m� �����ú%k��A�P�ɰ��lҲ��Ʃ�xn��	��	rF����lG�ȺYIO�4��zbN=��Rt_����H��Do�E쉸}�x'��=_"C�?~����M�	�(�^O7ѤHZ�������<��^����瓘s�c]����n��ܨ���U�J,���ގ��yi62��~������lpV���rײ.�=�����E�)�����H܍�k(;*n�}^1�P�TN�ʮs�ar�۳���j��7��L� {6l����N����lF�����`�D"��Gz�Ĉv��t��n��;���-7�-m��;�z���О�����s���<��	L�Ht�=�^^IPe/�Yֺ�l_�[yXd�`��>	y�%��q|���
�óc�Sе����i'��&y��l��~��f����[1L�sr���a�iO�<hu�3��犰[���/ڻ��1���b}֦��5u����A�x��k���ye�Q�)�3j�Xy�d�u��1VQ R�c��R!���en҉�)��\�H��NY駫��c4gVv��ggN�#�;�t�ҍ^�X�;����o�bډ��һ��yR�K��m�Ԑ[6�}���}U�W�W� :�.��&g�B�SZ�����^�ȃ�&��H�V�		����su��VZ��È�W����fh����o���N�t#�܅tP��CT��A@8�A�6/�&(g�:���',"���oKղl��_W�o���z/��h�������s�'}tU=/�l?I��~TqP���+���rB��ܘ�b>��&�\�P�i�kXZM��"�>�$�l|q�V��mqCz;T^�"�OJ�%�Q�����R���`�U�q���$�s䖿�艙��X�)?n�r�(;.�F;�劑Uf�e�u����	�*���1��򜮰���2}��SS�n���鯤��+�fȒ�eʅ#j�b���w���ؔ���j�u8waC>��{�2xN#Zo�R3�7�xsh�]���y��*悫���շ+�u4[z �m8��3�ܳU�⦾�����1V~ �|����w�-񉟓��S���ؽu�r7��J񴄞
�D��*��0�tY�~�Ly��`�h9���_/d������(���Iͱ�c�p%>��X�=u�p�Ϗ���@�XJ��29�x���j�ѩ��sQN�z�9O���XhΚ��ک	�mU���%,��}�e�TN�HǛ�/G�������~ 7���;H��x��P�IB�cɎ,t ���Ծ�r�՜yv�pU�)�O�isGY�8�VGmࢻ�T�G�_U��N�6fS���Q:X�������%��J�%n�6�C&D��O�wdWei;t�Biя�jU�����(�nV5\Un �mʹ�m��O����'�T�s�]�$��	�ʛy��w&f�h%�Xe�u9]��S��vX!\*踫O'% ��̧o6�`�XK����|h3�v��̫�"��Zjow-�5�@r$6�.ǣ�U�+-a7"V����
}Q�͔q��V�LEX\6lrCqKN����@K�[�&��U� {/v%{E�2��zU�]e.RȟtT��>B�m�Ʃ-7�L�X�/�e �kɑa'X��^�J�V���2_3oB���ն���3"�M��Ɛ+Y�s GU_-��	b��B�ש|��sx�r�'��]ނ�kO�t;۫���܋(﫨�͡M�P��gѠ�6/�8���,�ڥ(���a���.���S;/�ei�yo�4��eۛ�j�Q��n�2�v�+�+�,qv=s3X����tw}�0�:rHt��]��X]�VN\�>dW\�{��sY�IJ]�q>��t��ں1��6[�M`��䓗�@��t�LaB�);n�s���w)Q��M}��w��ܞ�v�|k����	�4��K�f%� ��e���<ǻz�Z�Nu}7��n�̬�bL�=FY�dEywH��>̹tCԸ4������a`�u9z�ǰ�]8g�瀜�a�4t� ؞�A@ta����W<�iR뽔r$��4���x��{&Eyn΂�rQ��E\Aa�-��Z6��{F���5KO��6�Ŗ� 1���m�������mqOz�O���1Mz-S[����뱹�.Wmf���j@8����G�4:񄲘ݨ��aN�7w�G����{�심Jq�P=��N�m�y]����ś���M�V��@l�������|Rn�`�޼['��$!��l�y�L6��7�"4�S-Wu��]�[i�)���5�Ի	ٜmn��Q��@(7�ص���an����\Ny9��u�u���'gm�g9�@	�1Ûk�cy�nj�*���w.�����qH��V����U�$$ٺ�c7ec(���Bڣao̻0�*J��<8�����{pu��e�PdpG5� ��Nj�q�C��y�WU���\��1�q�`_b=�ys�K5����k)�xk��	DR�ܮ776V:��CD4Hw�-]9�i,H�j���Y��^�mě)*̾��.��Y�[�\v欹S/K�ΒA^�I߄|[�gM*n��KT��y7��o-��W�֪V����N�{�ʪ{��[H�ry�5f�Y&+m*�
l��N����[>�Օ�����Q��o��6�}��e6�R�����մ�VR�UKo*�Uu�ktVSV�K4��]���G��G����e}�uJ��MV���smTV�յ*��*Շ�����ϵ������:*�n��d��55bMM��$�MU%5V;���jǻ�ψ�QZ��g|Wc��[+<��Em[QJQ-[U�R�G����Ef�U^����J+k�t��mIg����ݝ%[U����u����R�A&�}�=�|���I��L���۝v��qJzn�<zq�ًu�R�ݼ�+t������Y��{\U�(he�֯z�Y�w�����N5����[�?7'��qz�|;�yxm0�f�T�=�lN��ܻAEϱR�w�J�y�ۧ�$�^��J"˯�G�0���V�T���ESv2�ʎa�K���3��H��^�*Q�!O�<�_f��{aQ\j�}h31��������)���� vq�w����B�Ǯ����I:���OfnZ��tkB���(cgMȃ�*+H&q��5��E}6���3׷��3^��M�▛�|zY�t��֢b�ʮD�
Q��,	���}�������Z6����Fi�uU�Aɜ��1g˺tǗL��q�	�հ	�S�x�����	��}ّ�Z��'g1A:��ۧqV��Y��Y��%]&�	���{?c9ރ;n$�����~`���E��#��7s�xb8��ÅcvL^èA���H�V.��qԬ�����_t�V��X��$�\��+��X���X���6��aio����C�%��w]����a�$NP]X�|LdWY#=�m��ŉx׃F�$��=�U{W�^��m��O<�Њ����9�%���?�%�v{������t�J�M�����AML�4��@�vT�Z���H���>���4�f|-��97xo�.�zy]L�P)�mM�v�Y�^"�U��-�y��B�fw0?�_W��0a�x{�]Iͣ�F���.Z9�L���O.�)�IY��|g忳��f���'���u��
g�0�o7��[���\ı*�mD���7��=��Wu/�n�O�_Ĥm%���.�p�;ݝc"ȶӯK�w�#�@�:|,,bS
�S:�q*�\�<�m���u�(�=c�ܾ�1T$^�j��.L'~h��n���iz�28퀯���9^�-2�gsCu�NK��Re36��s������͛�A��R��#zQ�;��3o��;�O��E:�)��Pa�)��������
m�Z���(V��C�V�z���~�����[B�ON�`���J�u���MUu�{�����q#uP��j㨫�d
z�T��L���Q�e��=�^����ܺ�[XZUKZq��'��0��O��r�9���]��7������nn{4N��ST�f�QG�FlѠ3q�Nw������5Z�	.ƌ0ncr�q7���&K��������ak�!Iq���GU�V���;#�l�Ycz~�*��D_LO�lW�|t=��ߥ`�&��(��C*�N�������L�]L�ӱ���R)�\�[�f��gò=�`�� �u�F�&�+	�	g_�2��1�Q �Y]�̗Wm
�Z(k*�X��ij�0ӷj���x�y��
���W��>�'CJ���ާ�����c��<��p��f�6�����-H����"ae�
���Y6� ���Ð��rq�,�񞪷�qw4&��]^�1�cC>�-*�D#}_(&�.0hK��@J�+�F���*�{�!�Z;h��åUcG����;��?s�4�Rj�JXe(7 �j�2㚉V{�j�xg�%o3�b����e�Q�j�(`�҈� c���5CU%���8��37���i�W�z"m,t&��w�5ds�h�#�ݱ��|�5k��Q�gb�oV�\�a�Nө�,DF�E��`GM�0,��P�{�OU�Lf�H�Sݘ�݈o�eԀ�����ܟv5 4ϯvf�B��@�A>>���EЈ�H����Mf�4;jh��yNK��_�T4f.�T4���~�����kj;7�mb׬>dY�����F9�7�\h;n4�Z��=Q�绹}�踴�Hq)��2�ˠ�Z~%�&���5�2���g�"Ds3��-g���XS���i��ً�1�f6*\[ǔϗ@|��8�Y��v�}�ë��PŲ.j"�� ��{�*���_��6���ed�œ��mn=�	_zn��p�6���[olZm���0�b�^wm���8�f8Ou2�~M��g��%:��Я��iq/{�B��	Vv`�"�SjS�=�C��P�/gTΨ�7�����ޗ���#�"�� f�簘�5���o�6^]��8Է�]�=ˢ��3�<�_�yIԐ8F��\浩�(\Lث{�{ll���c����Dꟶ܊5�L�Y�M	�#%�������e�j�"1�t���wlB ����a!E壝�Sּ�Ӧ��%Ra�c��Z��߂����vr�7^2����!�]��Š����58���_n��<FD�鮴:�Wx�i�l�C�W��B���{W�ń��A�ipVjD�q���9�d{��wI�X���T�wf�}�C
���.�����ash����^RΥ �-dFG�[�g��T9�uޯu����.k��f-�v}��;��aw�d�Ρ�])��)gR�8���|��V�{��LC��"DLx�^��J2=��P���ڭb<O:�W�O�w{����m�kF��{5y�!y�e�*���Z���l�Cv�ܽ��P� ʼ��lٞr�(f���Uгn�	��]�{��Z8v��*����U��ԕ>"ۇ�@������L��:��ߢ�ۿݬ�3z�|�ܮ�=Hp�2�;�-v5�Dm�
�=��\ݬ؟o+�tp%���I��YTݚJݛ���(wS�Bƥx�*g��w&F�͘;��=n��j����D�[�9Q}n�<b澬X]����o�{�����w� �� uW���觕v��Ӷ/�M����/#��;�f]����&��5?Vg��Z��=�D\(xӬ�Kr�m[Y=R�����\���anP��Y�.�mC	��e�-�m���L�3oa��s.�T�l���u�ׇ*M�B:M��E�<
�.6���ׂ��k��T�HI�����;�ϴ�����4緕&%`/+�����K!>\�.(�[a��F�O��=�7q[ȧ)ul:F(�;��ts�Dx�����-��o��;}L��,�Vu,������Ь�{��Uz�;^�s��3|����ѭ����;ź���/��(^:�ڮa�V2�i��w��;��b���x���Xhj�T��ƎD�፯~>�k�]��S{��:�L��sh�o���*�$|�0�7P����Z���!���	����Bf1����O<豀D#̈��u�dl�M���(��Pv��湡*����^�.���|�Pސ�.����-ŋ�^M��m0B�#Y�m̶�Զ��+�c[�&�Ū����DA��\���g!�Mz/����8I�"�AH*r�m��͏F��l��?R�X���+�l9uiwq1����Tj�{�^5>�x��R�a�Crjm�g" ����I(^�4r��9dM����!	5��˯j�Ӝ�3fR������.魻c-�6f�������  �F6p�2��H�z~�p�+>�<?�؟�א3G����o�S/��`[3��?fz/��=�i2�1�%r�d odD�.o����k	�2n�/�sK�k��ѥv{�v_����ѧ>��.6���h�U�M#�V
���DO~T��E�n��͆*�Ѳ�Z���!��k�[ЃmM"n��V�R�Ԉ���W�$ܕ�x�]J��4�m�?<{*s���x|��j����	M-HM�UЪ�}X�*���(R=��ȥ��aV,w��>sc��'6���~�Ud׵�A�bT1}^�4��ŷ�J��x�b}o���oN��誆������'NZ������`O�P�8�fS-Je���m�-]cr�8���8�b��&��h����&m��v��4�?2<���
�]>?�CL�Գ�fc'�\�s��iۃ��b�헋�	x�s�pƄ���f6�HR7z�!K'7 ��Uֻ�̗��ѣg��򨦲)�>ѧk��]�>u�R�`+��������dz$���=%j�q�Y�!t5QVV�zɾ3f���}~��s�+Z:��(QM��3:�yϩ�㫲�	3�d;n�cm��M���F�J�3�)Y���`QVɚ����^�>��lfi���/�����ItWn��7ԮF��&���/��!���ߧ)��\����/o��a|?�}U�R�����l�c�F��K{��}"�䫚-w'�Nhn�d�Y�,IA�$��uK�0.��B d�S�!U��e�=l(�S*�%����j�]E���-�,5(�lse@�S#��Ϋ2^ꇸq��1;��x�Ð�,1�㝣�s�m�s�]u�5/��������\?#�(s1����fv�x�B�[����#�x�/�U���	Tz�C'��_z�9�2Z,�T��ʎ�k)�:�̽/�{Pax��#��E|�����_�_>3c��T8Y���Z�*dGlIW�q����{(X���*�bH�ڂr<�CL����¢��3m�-�ǉ�3^~��X%�{��r�sx@��)��Gz�U�R� %���>\s\ϑ�9���{U����_3_��;��e�̪����F[��}(���!H}�Mi���u�� �X�Qع-ʸ�r�Р�ɨ�x��iU��C'��3Үh�?J!ڥ��;7��';���[�R�,��{T����{���\Ԏ�ؗ�ò,לIf��d���e��\���{vٱ$�OLP@(q#��Z�gop%B�sZ;���޷9_��#ގS�Wb��9�^�$qE�i�l���e�JYV�j��k��uc��rݗ6K�N�J�U΁�=Z���p�{DڼhJٻF� �����U�x�m���Mg��Ld<7��1�{k�W#+�IS��}un(w�GZ�覞��(��䞶�T�u�[�V��Wo�)�H����<��W��:/�tR^5-�9kA��<�v��N�d״l��|n��*��p�D�-|	E��]B��ʶ�	��z;˯3�0�@)�� �'���%^�5��_nԳJ�gi�Dܵ��EEQE�p��ZYC�*�v�t�h�pwM���^L�-n��<ᰨ~���gz)�sz�����������P��$M�{?A◺Zޕ�?�A>=2���pK�?��ӊ��0�(ܦ��	2Yix�t�ks�kw�d@Q]��lc+w���#�`4�ito*�T�|�J�O�u��au)�XQ���y�n0Õ�����tS�<��|W���<�7�����L�`24� ��9�4%�����ޡ�jR/����h�������E����m*��_7
j�"��"nY��[�5��Z��K\��dj��Tm6O����[cy�nH�\z����,2�l��b��z�IGVH��� ���>��[p=�	�|/H��r�XֻJ�]qB���I�0L��n�'IeĠľ��6��'n��w3�͹��?c�L9�Ϟ[�o��s7�$:uT��RnGϛŜ�.��݁���V��\�;��$SX���_���*���n��k��f�B�C�����VQC�o� A�w�߲N�K}��J���#�����6a�j�������I���^��]��zX�G��,$Dű/~������>͎,�PI�_k�dw;�+Ӧ*FFz�t�v���.cc��$FE%>�\sR%]�l�v�]ʪ��A��N�g�b��7&E�y��,A���$��s��idG� b�U�7.�����V%+�s&�����Q���n�0����T�Ej�o]
�s�$�yr�O�P��1f�R���R�9��1�ۛ�j:�X�'o;��nN�>ᗫ���{���ZB���H�όx�gx͙N�tG7��U�J�>y��rg�A��%����W�k��%Rm�J��͡X����啲�1�ޘUU�'F��"D�ٴk�uK���wr�0`��L������[N�9�E��G����+6Ѽ�YZ�V��,�D6�ߕ|�,�&{T�񆽗�B�/�0�ƥ7c0�՜��;+{E��#�#*B賙�y��C�o�l�B�LD�Yj�E���C;_LG���j���U���_6�G`~�@l��@z��}�c�Td�Kd��j(�1����'
S�5lثw�Y�xG���@%�n.���qK;�-�3r����3�|��`ػl�EJ����3fTu��֗U�[v���� ���!�ӱsE05��Ai�^wM��2d���co�P�<я?S�=)���a b��}j��g�Bɂ���b���ϳ��֒+�Ͻ��^��UA[�yM(J�D٧�ө�dn�~ns��=VD�P0@i�	F�ᑙ1�U�M���V��]���x��E2��-��uXҠ���#�.��Ƈ^��|]W������=�j��tje��=Q�L!�`@Z}��ǫw��l1�㋖��MsF=I�-F(L1Lr4)�ۚ�Omn��O���')1⏓r"e��E�#��팷Xkb�Z9q[�Q7Y�ד���93gtS�艷������$�N�>�6�D�.o��5s�xVA�$]Å#w'�\���x-�ML�FmEug��.A����> �t�MP0�:�"[d6Aa0��
y��7/cZ�ʹ}���J�@���{�j:6^�,oF
���r�|dM��V�R�Ԉ�����{j��ou��oc>l�!78�U�׌�v�����)	�U"m�[@�q�+�'�&:����:3���t�v���;,���ʿ�ЦڽD�d�4��'ͷ�|U�����{��(��0�\[݂���s�[�W�ou���=��(�Ւ��$��u�{Ad^^���Չ���H�].�D H<܎�������Q|���v*KDHս�O�r7�#���a
1.n%5Y���z9�eg%����}�!�K�jN{V�s[�}FS\���;��>�Ӳ�.�=����__jݕűZ X�陜�_9}\�*�2��ɧL��P�� ���'���^�Bh�ࣔ�Z���mM�ѻ���=V���ڰ�F��Ph8��Q�
��[F1���U���?=�������o��� nZ���96N�Z4pr�P�T���	u��Щ���o�k�-Ǳ���������kT�[r-��}�����n�aΆ*\6�s(�w���m#�o+fଳ����-a@�r����w��n�-ݻt֝���"X�CtP�Jf��j����Sx�Sn|��Ҕ��e��!j)�k�KQ�.�s.�*^�8��C�Pł��-"��l���374�[���jkT|T�����7i=v�h�.g'���i'X����o'7&�C�����w�-6����A��ӊ��i��	�n�S�q��Bui)�%6�����ɫ-S���̛QTP݁k��)��%��L���ޑm)�]�^���axSf�����C��E�u�S����J��")��V���̫I)���Nk���@�4b�9I�v�A���<���-�2���]ڦeҮ�Q�;lͱXR��]�n�q'Us So1����
:�뽭�=1�*:R�U̽3gp�3i�O#G@nNR4u�G��E�eD�`�cy$V�?��yGԚ=���� >Z�[]���-V��L�upir��%Q�ig)
�Ю�p7A��=ofe�-�>7�k�U��T���^�$�e�Pp	lf��v�vsxCKAen��=�/KL��y�3���b��.����u���[r�rdxl0�����y6��&��׮	�!z��9�o��ܨ
�qEV�r��N�Eż�r6�5�'�G8n͑�e�=I&��K���O&�:<��ޫ��րo2��j�N�ɻIN×�5�ےj� ���V��٭�������w��Fѝ]
=m]��V7�q9P��
إv���S�:R�2^(e�;,�;3�f`Y�^6:1-��D5�,�\��ƺ�5e����2ekv9����rB��]k[I,S6n�gRۮǐx�Yo�Jh�c\�9u��Q�e���hE���t����.
"jۻ
�*��w:r��#�fuf̶������M��V�+ݨ3Fa���It-��vM��AsX M�]]\^�n�	0n�\�<���]���q�bX�PU�|���$����Dj���U�@�A{�h����Ƣ9$1�k�C%3W�p�ik��s�S�_f�e�5j�Ay��#F��ʑ�{ltRW��c��˵JЭ�փV���R�ޒG��\��&�q��U���}_1k(��V�F��Ujt�E���oV����U��y:�H���:%Tڮ��m�ij4���䢷[�W[u��**�KS[��Z�9jQJ�Y���St��g�[�ó�]��52����ج�t�F�����ֳ��jح���5l�c�Q��b�Q�n���E��+u��g�vg�u��mO&7[�:�PV��u�Q��:��}Y�
�m�f��f:ov:��Q�՝]3�XHح� �"��$``��B 0�������c����5�������61ީ���ȥ�7�q��u	L=1�M��k0�c�7�9�3�Ι�K�6H�F�]:������ զO��Ü�ׯ�ze�R�Y�h���!఑�e1X�S.s�.�n��^X�I<'aynل�u�oy�2`U�?\3cX7��t&��p;w�A/9z�䡦A�r1���wJv�Y��!S^�mB̝}��V��P��Q�BtC;_\{�yA9�d{;1��VD]���Kk�8���}�u�~Zt|�"�l
���""�Av��jsK��-{�PúuKb�CzM��⧓�~������Cx�U�#���C�����3*ec���2�0@DG27S-�s����J����kN��c��5(�}�	͜Y1�����6��ݲǁ;�.;J�\jT�3���Y��Z�q�{�w_#R���j���8��*�zd[u�h�I�^��Hɐ�X!��E�M-����i�{m��j�6��=���ba�������a3_�sN@.8�����Z6�w�ի�ܽp��"���u���cB���b,"r!�
	�J����P�8�mZ��Iy�A��i�u����n�V껋���{N�5�☹`9��`K���p!�S��3���ЩNTnZ�S9\!͌���
*���T[�|bKT���\�ԷԥX��č�^�:�p� ֡���h�V�M3fwr��d�ϡ�ȡ'e:|�ʩ��.S��=�3^���p�7X`�X@��M�����xY:2�����ld}G��1�z��-N��iD�7�.~f��`�����n�;�#�~��!K��x���X�n�(f�rs�������by5�(�l<Q/�5�6���>��,^k����aTK^�J";���GdZ����Q�'j�+�?.r<���̫��-��p�(bוG*E&ڬzG_����n���M�ܲ�I�x����L����	�H�_�~hkh�$���f�p������=��� �E�۫�eڸY�_��!�)�ڽ%K����*8�z�,��~RF��T�:&�_�T�{	DZ�k˨_,�a��&�%��{.�<c	SO��tF���Kz�m��,}������x���QE�p�$�+��ȶ4`u�CXj��ͼ+��+���%C�R�2<���R�}z�}��|����{ٌmH����*���ݐ��r�z�T�,������T%K[���N��M�2�jB~�FN:`��\��5M.­S����*磻���/��=���^�!�i�6�~c]{a7;;�P�N�ks�V��۲�tC`�Qw�s�y3.�n��	S���oa*@0���y=;\���u->��ѣ��ņ�&b	벟Aqh����9|�3���W�����?��Yh�u�;7;�fO���/<�Q���w�t*���h�ۙ�������L�S��|�C�l�g��%�%��p~>�ᨺ*�4{n�J��}G=��v3}jn}�Y�;�4�"�HZk<vº�z�Q��=`t�D�������||�'�krb�ף^393��vs%��y����kok�h�Ԗ|;�L�B:}�WE	�U�R�(vMn�w�K6�;ԯ#=D{����L���F�W�r~�贳���:<|:�mtx��t��[19n�|�W��%�ҧ���I���SMA�3,/��'����i�kXZL^`N�p�F��4��;}�I��ܬ����_�zD�z���3X�ڽ�l�h��tk�����|�.r�ZKy��"�Ԍ�l��n�$�M�:#gΏЏ~U�~��N��R57��a\&С��z���uMS�Lr�^�5-_?H�ᮬ�/=
����b���~ty2}QK�=2On%���?n�]��j���bK[M��֢��ۑY�%Y�.�jۆ��kg�d.p�5T�8˃�����%��u�R>�8G�w�c)���%��l�當j�'���;(n�`�@�
���ۥ���>��Y����[��:��RM%WI@w(Tݗ\j�L��k���}��)�뤳q(�;��\)�{ۦ����iSV�Jf�u���f�}�����뙾�yA���K�g��}f��X�h�x��8%>\l%�3��VL���e�F]�ݱ)Vѿ[��-]ȟ��Pt5�.} ��r�x.�m;.(�[a��UO�7|�|�������=�ߣ٤j���D�*�+0�/T�x�#�)j~��!H��dV�K<���c���+x��ނ���n'��r�JJ�ȿ$����ݘ�=y�;ȡ҆XuCB6��0�\ݮ�q�E����GO0�P�ϭC�{]x($a4%ô
8��L����+:���x��[[�׳;
R ����qt�O�1x�+��.V��Aޕ V�Ml�j9��0Е>>c4�e늫w)�����QL��=E�@q:�n�K�XO��?:�6k�貵W"��©�+^���E�r��L.�?4c�L��zh���~\u_�xjWw��3ˁ�/5��&m��'5����X�!ldg������iB}"#"�\��7b,�ÃbYY�v�Q{ld^�d5����;,i;�6_��J[CbJ��}�7�"e����5�G���
����q�sr� DW���'+Y�<�r�ŧ�7�K�[Z=٫v���Ԛ�����.<wk��X�fÄ�u��rj��r�e"���ƫ��ʙ��76��	ޏ)Õ��;dZ����R0����)gWX�;%J�}J�a+z�O%�O���.��u6׸��`��gO]0�4��7D¾p*o�}�r��;������K�{Z�Tnښ��(r�[�ZD�9�A>�Dd${�$��W5�������[��U,y;�w��q�T�i�4���3�q�9��b��r*�](S���~��V�\G)�J���'� `#;{W��:�W�R����]kk�E^X�<4��8�YUL��;�^��:�r^���]
����}%�h<+z��q�mn��y��K2�l�i�x�u����[;*m��Q���P��5��z�A��Fdp3���K��ʡ�]W�Iɹʺ���F��.��	�m�f�j��'�=6nUr5 ���btC;W��z q�K.]%י�>��W+��Y�r�<�jyYx�N��]@�T�yU��
�������*���e��S�qCi^�z�6>�lK)��-��v�W\�k�<jbcx�\u$1}�q�̅��p�ay�1�*0��;�S''-���O418��a�Ⱦ��/J8@��q��Ox^]TKw� ���Z�t�9>P�rO7�j�Vf�&��∅w����M橕��@���P޿������^�	]m�O�y�2����	�ΛM��r��%�{e�Y���NS�Ҝ�/jW3�e�c�&PIa'�&O�՗�ч�w(�*Ϗ}!��K��ymm���n�V���-�^Y^�}�-y���j���jf���������zW����>PN���5흑&��[V�OmTg_��s3��vp�i��V΁;"0�O�Í�C��ֆK�A��?B��!��3���Ѻ�x����TN�!�X��[�Ө�J��Ϛ��#���ޔM���"VIe�-K�&�j��}u\ �%/ٖ�����C��D
�9�A.�MX��J�jJ��N�m{M�b����^1�ژQe߅�������Fh7,��J#�Gk�AWã�E5���+G�9�{�;Km��O)	��������}욲7�����ܲqW��4n��F��	��LFU_��J�Ǖ8�s�(��J1[c�{�@��@�Y0
|���O:�n��@�3���"��\]����GϺ�xw��I��"��ho�т1��	\@��Rh�[@��ޙ�׸�7�{N�V�ݢ]x���{TR~��)���ǻ*u�^����^}L;��N�LW"���ü�=�f*�f���;:�>��i�s)]F��;�㓠\/c������RZ|�UߝO �%��OJ���]�v��	����
�C0ż).��������鴪�Km��&��p�¦�?ti-�]����2c�Kbt��v<e>�����M��q�7���1�>~�%Ń���Qi���_Rʶ�M�c�쏮��ȵC���%:����T�p�i0#`�u��r�`���q<���W,��w*���=�H$kʩAB+�[��c1�� �J��������F��Ԛޗ��.>ױ�u:v�e]1�2ӊ�=�/�x�ԓie<��*;���VЮz�KH�2e���hO��v�b*��Z�X-V#(�C�v���GT�ӿ��d���F���>\)�˼o�^��ԫT���yL�Ķ7R\U�z��s{**�0�L���-l��O6���O�#�R�F-*�C<jP��͞1��J!t�d)׽=ۭ���`c�e���ll-�5�T�5C�I#�lԍ.�E���Ec(#9���Yt�!kN���dv��`���cmމ�a�l�/"#��R�w�qЙ��!�f`����y5��7�HL�P̢s˽����ih>��$�29�Y�r�֝TO���58+�Ku��B��%�11�z��b����oL�/��b�\/mO�ד�͖C�my�2����N3}���U|�Ѻ�ܡ�Q����I�m;˃�nIQ�6�����x�{��)��Ƴ�7�ea�g���C`�˩�ī�¥��[�<R��T�ι`E����m���:%��P�{�۽���c�!��ˈ�/%%usU=J?�չ�u���:>�o�];<�TۿWG�TO�<��{2.����ؽq�x�A��J��7�=�v�s�]u!}�y�2!����l�j�q�y�3n���|s^��ǘ�^��p2�Q��|����� [���Y���Ce��%cU�/`v����R}�
ʯs�k�"��*�6��Y�+����S
A��5��3!�Wj�:��A�Q͍\a2籊)>ߖ��*�\]�[P�}yڸ�������QM\5���o4��!~\L��F�WtL����搶�������]�Ը�oV����Qޕ����*�B�
Ձ)���Go�>�t�{�l|�jK՘[��3�`,��V*�QΦ���Ӗ9zc {����(�3��BW��Ե?m�ECzY���*�Q�l���暋�
��L{|�$s��:��1U�Qv��ghL�^��<�$��T���uRׄ���A�ۈB�]=&���	2Y'�H|R4:A�ic��7.ق�#*&n� j�&"V�e���TyB�'c*e������u�_��.+P�~za�9�2A��M@�;cf[�3ٵ���/.v����J��6��Q���';��_lb���6sr�}���>^�_��H���8�c� �_c14�Lv:�'���{b���Ś�dȻev�����GU85jO����ر�O7i�^<K\4X��|�7ϯ��ȿ7����f���&`����қ�N*���G4]*�mj&1����b'�����ut�g'-�i�n�ᐁ��Mz��j0v����kS׉�l��ym��W�S)�[�㲢��:(L�����T�@�W����㷶�l@�+g��B�N�ř}����tz�J����:ؒ�u}�@��H�����k1Tn�淛M�[F7z��"�6i�[�u,G��lk<'[� �蒚��V�l��bl*��w�1�d����b��omQ�C�z}�8���_���
_z�:a�<Kf��z���h����Tq��B+x`Zn��۬iUM�~���&�]
ǽX�*�ܡ�<��]�ʕ�=��ͩ�KJ���Ʃ��+�:9s_q��ug��k:��{�U�����`kt�7b�����]7�� V�C;;�rn�2{�4��܎~��Q�<E|3fS-�s��g/����k�U�}+[5����Wz��kޘ⥬�B�ޔn�/U��o�� N�KC�yz2a�$�;�%]HeaJh�Fm���l�eH���g.Q���%�������=S_LӷYS�{apݴ�-��.��7mr�����p�q��G��u��]}�L5�:b����n]s{}=!���e�v
*�?��l#�����ͤ����&,�=uh��r����uM7M)8�s�f�W!�A/�r�������D�-Yl���u_jǏD�G��b�o#�Z��i�����@<��+(r���������~^�f٧����-;xe����>�&(E*�=���D��y�1��r�_'�i�78)n.�����#ͥ�^��&������-F���Q����n4�ȿ��SY�Q�\�S���~i�L�Ol��B�Ѽ�ƦlJ��~�ͯ�:��9��om��eeO[�������fq����K�t����'!�u_,�MM�m+�5_B荭�y���|ޣ��3������.7�\~�#�>N9��ၒay���.�n�E<7m�M�J�3k���Q}8C�Z�K[�(9�3~JPB��Fp d��G���܌gN����d},�.3>�݆�������ڶ��0-�q8O��i�Ѓt��]���<�y��Sۅ��.~P_��t�	�IX�\s.ș��B�/P�]�P/�[Hw� (  =�[c|����h�FLHc�vn���74]�In��y���'�$wq��N	9�<}[M��]p���݈󷠉*���wJ�XB��ʾ��)ueBw�e�
��s����i&�āNS鹝W�r�-P9�.���� �3ne������+iR�HV����B�d�^
�k�r����*�G.�����jV���n��(��f����u�3�]���ޫ�1�8^��]���4q9�l��N+@�B���%Cr[{C8��ɷ���3����&�m����X���9m�;+R��P�ֱ��FM���{��?���J�?s镆����GB������m9*����&{�WPY>�KMňҤ�7,"p�Η��J�`����ّZ%>C��/r*Oo6V��zL3��t�,Ϥɱܙ���8�U����2�J/�b�Gu���T�{���ؑdW�b˷1��;�/\]4mu��Ԋ�o���=/�Jda6���`EUf2rVQ(�<�mƊ��H��r�������VP�����{pi����׫S��SsR��Z��p�������ˤg-��^��U���Sv���K��v7F��d[��@˧\�d�yb���ZW}����Y��%�b<72}�cq2JJ��빴)hV�7Oq�"H�E.���K��+��'�rdmފS%)�V�ۤe Ui�I����uЬ�MN�l�[j���/�h�*۸�^��ag�Г��:�`��y���ia����TuIZ���&���2?Y�h��6L�T�J���O��:J����P,V�ّq��<�����|���ɹΛ���h;�K8�g��5'P��j�+�|k�Lk(�^˳*���.���#�+��̠9,?��3{��&���򖶸]�v70F��f��'�o��D���y\Ԯg�	�5��z��0��[ml"Eyƿ�8Gw7��P��ԮT	<�r�z�̗����wc+�>����r��(⧸�̡f��1��+�X9�������w�޾�mJ����?]07k��S�~�u��ۥ:Cb �7q�o{��;�Y�2�yu�έ�(�E���E�:����ͬ�WG�]G�gh��:�SJ7����n��,���j\5Բ�[�(A�gsh��O�4v�����of�TD�T�(�[������%:#v�Y�3N�o�����깝��-��e�n��A"�fvT�;UZ���H����$�t�fڟ@��Lv�33/��S�ͻC�%�GU�w}͍gm�^�Mj��}F��]���S�I�N=��얹�|�gocH��2FK}�4>�/�9긠������]h����HM+������j�p��p��f�Ƈk�&�hwm)KZ��a��Lu�[0s�:��]����KH?��O;�۶��%7E�＊�^���?}���$ Py׫��y�y6ެ<�[PPj�[ycy7[o-��X�t�U�n���κ<�M�uYy�t�����+[ic���]W������Vڳ���;=�MG��:�3��Jg���:f�u��Z�����l���3�7Z�c�wCȭ�el^s:�ζ鳦�7Y�N�wc+ɼ�^��P����ycɼ�:ٺ:�B�}L�o-Y�ۣ�n��|Y��yU�����; ����7��BjmˉӘ*�p�[z�]p'*-��6�U�0hN.hݼ���znS5>�������t{P�t��߳�x�>|�M E���MG�ھ�U����{�h�q��7퓹5=vMY��5UƘ�#��$�x��{OB1�ʑt#$S,��SϮ����xX�-�^y�PW��1к�D��V��si���	c��F�Ч��Q0EC�V:��d��p���c��LϹ>R#u��96�?�F�V������ �E��^+�u1�]P_��ɃR����w߼�n�^��Jv+��^���(���'��Z~T?�^���ռr���c�g���a���U��kޮ�����lu��/j
3������3:��·r���m(�1|�F�����95{���� �T렖�l�q�P��C����3�K�Z������.�{8R�a��/���@��Wp��n<�+�����ᑬ��d�
�R%K[�"qNۑGo��{��c��:Z3p\�n����Ac��X�)]�i#�"08�[��N��ԫ]:~c_H�W�ry��.�H����g�\/�u?j��]��?m���4�H�#J��Z��U݆{��vg��=޳�k�gv�:�[ېta��F�P�Y���p���z���fn�<����L��\��e�9[t;���˝u�nl[I�a��d��v>��Rn���[�W�6���|n�=ŀtèRy[.�ɵ�Q��dD��gPf`�����%l��}���i/��=C���N7
41����Mi��X)��:a"o���vk'�%��Zb+S�H��8`��q��㡭�m���۽x��Pfˊ��+�����o��[L(��1�ڠ<�\�g��+���N��_%��)m�C��rZ����!}*k�|� �Ae�~�"�O�����/k���wy�7��x��c��z7��X��Fv������Y�>]t�����VG�TH�:�{�z�ܶ�UZhe��ٻw�{�쪻�u޷enƾI���Tۖ��A�[��K��8Jz����^���=j�W��3<io�K]���R����:�t0vy�5��"o��(�yr�Hڂ?u������D*�_�B1Zfŵ�d�����B��Y_��Kc_��e�`b�O��(^�J��fs�ahSm���S3��+�֏s0���l�ҷ��Y����p��	>�J|�[B��Vr7*q����Y�[�x�"��^�>��3�"7�Z�\ڹ}��	��\�{s2��켠{�o�@j���s�/+��ί�R�m)�r;Ź��m&?.��|�1���"W��)�B��^����.�Ubq>Og.�4���{�8s$[�"!�P��:�.!����f�u�e�rF5/�����m����}�C�Uvʹw�E�n��V�W���00o���6���[�`8o]?���}�o*�|r�C�Dsw=s��>�L�WҸ�f���Al_0�'g����=��$�"�Z�����2�x�� �X��4��dU�
"�Ԩgaw���ls۽�iI��3{�5N?v�	@�Q�f�q���:��n����BBɀ\`����ʑ�mż�۩�v�^���c���������N�T��ө�dw8��rǌi�A��PIӅ�Z:d'�=�4��� �]��L�jr�������u]x6�(��r�[�T�ٝ#��������w�cޗEJcQvT� M�Rr>�zh��;��|�=�Pލ>z��3�l�8:e�Y��h.��NR"�68��‟D�S�|��E�a7-�CT�F�=��������c��x/p�+|r�\D���T�ڂ�j
��{862���������w��L�}�bE���χF S�h�K�X��@n|A��Y�PצabiA��#}Z���5�� �θ�Qۑrvu������e��c�0r�k�X��
C�R"v�`� :��]ȕ�5���c(��,'�T-=��V�5���=��lK}u����H{���[�'��+��Ó��,:w�3+��9Q��͝^{9+$�z�Dg��-1�����3�٭��-��w�vV�DYf�΍����im�Z2�E0��/*�'-ǝ��ﾡ6.��{�c�g<���Z&�ٚd{�]1k�!6թ����`jƑB�8oP�^wůo��MBa�I�K��Ss�P���^0
i����Um�C���-���z:�e�5��5�i�ENwwM:���yb��}vu��õ�t4~Fǿ����[@�tIas��-���p�MucV��<ר%T˜�H�1���
��x�	�G�0z�Z�T�YO��]�D�Ѽ�Q5�8n��JdhԳ�������]bb��a�M�G9�ҮY�U����:ϱ/�T�?=�|�)s�pN)�>�v�9v���EO�`g��	�y뽙9��
C\n�H�j"�F�s��K����LH�*t�u����^����iul4I��6j�ު\��*��G(V���\A,��Tɼ�<h��n����ƀ�i�q{V�����}R|���w2_������!@�`�!]�"��4-[�	���ߏSN��|F���E�콳U���ҟ3L�ƠH�Gk���� a;�*�a����|�e�"����{m!��WZ>.�W�u���
�gkq�{1Q�Q��k�+���9l��a�=�����l��h�In掇�!)G�"�*j}�Yy�K��u�٫�4�:�s��2j)�����u�z�^۾�ڔ�T��N(��Dz���s�m7S��xz'z�[{�����LW>}����g�Q��n�uތ#��Di�HL����`=�t0R�L]�鯮�s~2>?ya��~���˟��c������F��PMϳ��A\1��Ѽ��صق��Κ�P��_Z&�w6ô��n�0mq,H*m8z��N�y~g.ţK�M'P��*��o��N���pe�bL$�/�o ��4�۸kI�b[��rH�ȡN꺝)~�0�P�_Za7�KUr������Q��z5���׏�j�����[��m��Q��/2T����8r"�3s��k�]��$�[�O�R^�ڰ����
��H���vһ�[^�Pqٯ�:�O=t�:r���k��N��a���7
�/b�K����Du;��aׇ�]<�/� ɭ�#P��=#LI����QI��["�k�M��Q��ۛʨ4z����Ff���G�Ii�죗��ྍ"B�t���j�n����Ӻ�{�=)�%�eO�u+/֮����[�G"3���k(F����cy*-a�T&���%H�v�U)f~�����O���5�EΤ�a5Q�^�A��]��6��7�8ػ��{�/��6���t�%�L�E�܊U�;��q{��ĕ"�B�9!����*�;���ֵt�`N=:�eZ�L.ȹ��Ѧ�
�/��s_C�����y�eM�����o�� <n4E[u��C>U��7�/���K��_J�D
ZY�e�o\Y���|�gl%R�%����ƅ�u���?6.G,|��J>+�^@��uW�T���:��H�Y��Ӑ.������ŧ..�K�������p�� X�.�^��wm���q�L8�U*u>W���15�ގ�.��[��N�~ZM��c�Sе��/:zҢ��M��d�ZVG8�6���M�1�����C&=���b����J2<s^u�3:�^	3��!�7O$wi��a��e��c�
�H���rZ�/g�>�2N�{B_i:�1Kj�g
�Yd�l]�ݟ2���ژ�)v�/4 �^��!3ήI���3�PތKj��x������\�������﷊��p/��N��ڥ(���}g�.l�g�}?J���Y�~�mnM�T��;ba֔�i6�xǉ��Ԋ�������eiFyTuK��/A
��WGi�9��5�
�Q�1���(�Cׯ!�6�/�����)}>J��B�_	4�`;0�Fvڋ����6�[w�G\�[�i�X�1�*��Ӻ��c%mfR��n��w&���Z�P�]�C� ܁]��f�;���k\�)Nd����g)!�\��Yq�e��b�5֎����/*��.������u��Ӡ��nCE<S����� p���=y�
�'܁��O𻩶
2y� ��7�R}+$M���ȣ_<�P�j'O<��|�r+��j�;Y��� ���W�'�]N�lJlk�	�=�R}���Vk��0G{|xE�**���㩴����P96~�\LY�2�R�_\��F�WQr�d��ˋ+pەf2�"�N��r7b���\Ŭ��$$�Wr'��#�j�.G}!�}ܥ�����]Ǻc*#�R�5e�L����%>���~�9��͖�#��^�<ꟼ�����11�+�X�t�e�ةL'�=�"�Գ�X	Բ���q��HcJJB��TE����i� L=�}��sY��E���<��P'l�J�w�i�WأH����Vk��!d��+��Ӏdˬ��ŗ���X��t�&`�W�t{���%J�ke˥���,%:\jς�3k�[�j�_�vȳ�C��2	���3˼*(���-����⧞⼲9�{qMN�Ъ륙���z,O����a��cv,�Uȃ�P8�-�
NC!�+�4Y�u����>�^GN��hOJ���D�S�Z�E��3C!������X�o��AmR�eCY��F��1y{�y�/%�"����!;��M�Q��ri�I��-�R����`�������~Ku>�a�%{�O[�O�`̛/d켟:N&؛�Gh7�sr�Y?��͋B߾�R¦OF�b��B1������߽{Yc��Nr�‟H����_	E�"~�e�Փ���2�V�<���#y���_#��<Ꙡ��Rz��]�#��"��7�g�S-�WY�0�ӳ9����Z��л��[��Z�N9_k<� ���E5��'�s�,����[>�Ռ��b��p�6]E��6^�V{Ə�q�R>�_>2&�c�H)}�D;��f
��Q|��D�����U�J�8+*���*��)�SMZ��ht+*�ʍQ���]�[�*|���wzT&�%f|�mm>t�ڄ8�g�
S��~-}
m�ĩb���m�h��l���ʃv��,�l>�������yZX�7h�/�%6��*�S����+-���RkX�z�A��yݢ�xq�,w<�S.r�)����aEFd���b�$�0�)+03�(�L^���훂*���C�{��zD���e켧DPn���׎��ű��^7�x̀b ��o��~b�a�m���u9�#��OM�2n�1!�༩���6_Z�Ӳ9�Z�� ��|}�%`�m�牀����ind�Ks��(mw���;P>?4$;��<���$:�P^��q�Q�o�W1ػ.�S�W�DSLwu7������J{Il�Z�GW'�U���K�=�0ۖH����cz�p_f*��r��݌)���ڻfΟ{=�����3ǔ�F��	�msY�@��r��^h�K�s����ˎ]&=*��{]�;�]��ƮI@=����F��g6�d����7��IdZq�yg�>Ʌ�xH;7��\o���P���71��G,nHEl�
݀��bgCB�V���F�����/w���(�?j���z_��Q�mV�.Q�� �䩁=tPw��j��W����[_���޸�U݂[�㮝��^tg��8�m��@��TWӽ�0�ބR�PV|�"�Ƶ>ʅSv����Kj`)�c�?HZhm {�a|�'�o�x8�k�#���d(���,��P	`��G^߄���t�[��h�����Ln��;��4�q/<�Y�v8�"��̜��'���	�CK����,ɏ�3*��כԌ�nX9[C��}�J�bʯ���Y��m�4��
q����Ic��N����"���{��f��^�5�R�.kp�9j����}O��=|
�ע���I�@k�ѿwH�yQe/r��3|��Y�ez��h�C��x��3�&r���XaٙʫAZ���so�0ձ]�����5Iz�N�p�8�H�lzR��H����%������
�{e7]����%5��m��C��$Q��o1��.�\:T�5jn#��R���CHۙr�^`̩�}�G#9�+��V�<�ӣ����͏;�]��7�u�� ɨQ,����({n��\�MS���P���H=f��k>��zc6O�ٹ��#����rF��1.׳b�|���>k� I�mյva�R�'㹬j}�Sy�r޷�pЦ��=�Z���'+� �s�W�\�Câ]<W��6׿mr������a�[p�=�_�vw+��M�}~���[�>M�=NfmIG[�<�ޏT�dd��*�i}Y�OV�n��n��[N��c��������>����qM�߭�p:>ݕ'\�3۪�(7G������[���IG��"���*7UJ���YB��I�Z`\��t1D#��3�o)��K_V��8כ����D��	^/$�dF8�&o*�n�!'ӳ]rƇב�5캧��	�XJ��ml�Bz����;�~�c+�4�����W$}�ܝ���Jee�4%n*�5?l���Y�C�euc`-4#kʪ��%���R{�ow�Y+��qZ�w�=D���~wf[	�C�sY�=��sߌ����c��a� @p ���0�6�4��ƀ�����xq��
� �Kז��X�1V%@�c�b���:R��:�+�zz�.@ūV��3(ӻ��?wT���.�]$���qV:p����o'sOk�{�	T+x6�H-:͂�mwC�{C���Fn�:�w���^���!��qqV�	\���5}y}�`�Ki�ip=��m�=�R=4Ξh&�����
Kۧ�����ܗ�l ��ߵuM����yPyVhA��#:���.�_�7A�X��g��؏���n �Mh_S��kP�y�5nv�hoN�wo�O�h����u7oQ�������l�tu9]���[Pf�(W���pQD�p�//�5��tS�iʆ��b���0����Z�,n\������s���9�s����#�Wk�z�u���0u`�̑Ll^n��9�.�IZ�����%�\�K��h�0\�ZΎl=�/;����Shq�ppN5�3�[�\s 
h�(�w�w�E%Թ�ol�ݱ�H!Y�yc(6fܵ��ӗ{M�i��p�lRKE(��"7Ԩ-�-�Q�WB�F{�h�Ygv�\��X�ۈ|�hᵜANcUf�GoKbf;����id�q%3]A�<��96�t�'x���*��4��K\���zm����� �BVQ��Ͷ:8�q�F�������ի�d�iU�r�Qô��Ư�j'����嶷��a^�V�4�n��4�W.�EdCs0���Z�@�J�z�����f�\��i��N�U�N���,Ih�z�;h꾎�Hu������I�[��7�;�ڽ$q�w���%�l����Owab��n�BZw��}��S��4����X.X��.	��6t}Y���6Nt�c̛�!���fI�r)]���݈�9���HRl�!a���q]�ӱ��4��Ȩؽ�9�q^Y��(�L_���d����ꮦ\� �qX�m�56���{��K�Z�ɶD�y6��L,됛S�ފg���0�K�2���-m�|��6�}K$�D���{K2���}r��;��n�'�S�o�wWN7-�sm,m���9#s�r��
��ݹ�-���}�b-v��&���'���(�Hz=ѥ����u��"��
��JY�r�_E��%���속�;+��58���)Z��N�9���N�����]�F%q�ܰ�t�9s+�k���#yswe������*U�@T�L����ٓh�5B�]GmG`��تW8�Rʨep���\o1�걁�ƅ�d.+����)�w�77����2q����hRz[�����qs��v&��	���n��n`�ܺ���si��5�NW��.o��^��,��ϓ֫�b䲲�iIR����<���x���)'ӺP�X�ۙ�[�cspܢy� P8�+I5eiq��w �zs8k B5�בM���uo_�Ca���҃���h�lK�1X�x�܌`��s��4|�f����o����ѷ��Vn�z��ڙ�ۣj��=[t��<�3t�-����57�o*c�V�M���jWwyo&t���uT�峭��/v�g�=M���۬Q�Su��[��7��mCS����V��Y�^����t�t�l��n���yT�]m�ՇM�o&�6�mO,t��[tճ��ҞLtu�ZU�鼇;��=y��ϙ��l�g��>,=Y�&�]u�u��j�G�����x�h磏a<}{�U���*=���s���ѽ�U��PD�}IZ([XS���[t�)�����=; �F�j�[R��֛%��U
UD@�g�� 0��X�sufC��	�E���P�/��dx�
��7C�߳�o@`׷g�ݦ�߷�9�d��r�jU�&L:���$�g��Ƃ��Mi���h��.��z)�&���e�ac��Կ8�;��鵻;���iCZ�|�D�?Rg��ۺ����!�^|�d\d�P��hC�Vd�ǫ]
�ƱZ����F�^ˠz�p�t�n�{>��>�%@څ�hDz��T�e�����h�I��BP�J�e��o>�7X���=Y�C׷���~�7C]Yi�ʉS��i��&�]���}=���X<��~ty2n���R+��è�h�ކ[^�[�k<]a��.���q7�<�{��k����@��#֑��?@�3f�s(H��r���̚-~xR�uO��O �{;r�/�����V/^�e�������o32.U������G} �X�FG���U;�ݯUėO�ՆQLu� �����=�e�iF���~�k�����'|�ҵY�h�i޾ƳxeM�:�y^u�f����s�9����,L�$�4�2��W�Ž6)�N>:�;�%]_�l�fj�T1m�\6�Ԥ���K���-±ː�9�}1�� ,nX]MZ��o���	öf�wu<�`{���.���q�}�ԙ���y��9�A�Ͳ
8v������p��,�.�ƱZ�6��'��������+�)S_���`E�c�u��N�F\P�y֑��O��:F����~�h��#��}��(K�P��dh��+w�la,�6�w/����\ب�G�g`�J\m��t�Gs�J0���w��s'W��n;��5i�D���@pH%pY�ac]^��R:v�{��C
�{��ϒ�1[�i&��xK������9����9x�X9w�-�
~9��@X}����=_N�����D֗�iY���N�ַ�kLZ���c������)�X�_`�� �VFu�_e�����ݱ�f#�y]�g3�l���[��/���'��'�
Ok�#�o�D����x㤮x]�S�ne5�|�1B>��p�vK���,�zG��> �颚��X��U�8 �|e���7�»|{bu8<�F"=�SQf��cZ���ZE�0�8�A��9!c��	�<��-ō����������Ţ��C0� ߁Z׍E�yP��R=���n ��1c��3��Gj�+T�:ޭ�g�P��#�"���x~j��iw����fڡ�S=��R+&�Z�t���U�U�~��/�W��h5�.�}���%q��3��ZEAE�߰�X�6���zl!�QяB5]����Wؖ�}�V>;zg*�v�A��<���Ke���u.��5j�����9cW*{�s�-��m޳�W�n�U�/��$\��O�y�=xk�E-������PJ�Eڱ+�W@��N�?ua��=׌��G�����I�m̱/��m�j�P*3&�uqA���l�W�r�(�������ψY������_F�>^-2<u,�޷�=���]
�B��	Ž7Ę��0*��`��'�e^B:xK�k���tHW�/���u��)j͵�;��Z}ҷ@[q��)y���}��"�
�V�Q���G�Az6�A�~��[ε�PK�*��f.�4���ˡ��-�W���$��:�ңH�"!��
���1Ijc��S��ޛ��.Ft5����wG�-�q�����	͟���A��J�Lԩ8z4�9�!J����� ֑ů*�U7ϰ0���!��5?>��]���::zD@�-�
~9��H�":��5�z�f_�Y�T���k�T�nw��xώ3�8dFW�M{�CC����4�� /r�=�6&��SD�����p�2	ʮ�Z�p7 =�,�V�Η{FE�
f��1z.ڸ�%�~�<DUy=|(I���g���x9�z�=��[=��=�OYO�.��k+5^э�����F ��h�����bl2���orn�rdW�}w5��%�V��k:��!��7�!��������A�ǅ�w��LZ�۱Ӎ���j�O�����M�Ѱ=b\/��^�k	�H����l�<�l�8j9�c����cն�s�<�PN;ԵWܥ,2�����^�~-;��ľᵓ�Uoy���/Kh軸d:�\��A�,��m!��9BW�K������f��ʚ� $`�ғ���X�'x��=����s���mc~�7�wH�#�"uR^�Bڐ�H�2E2�f��퉕4�7�՞�m$�e�Ke_T1}�]���O���6U{�=j���5?]�`<�����ʃC�5���ѹ�CIu����ߨ=�弥����5�״<u��7�l�f%��K���yךюf>[�Ix���9B�A�������<:%��ڦ�y�i�{�D����[��{�Qc}3t����f���@��~:�p
���;���\"����UD�t���ÕnLB���IPE�֖P�
������E,5��(z��P��,����F�A�jə���Ƶ�w�YxZ��u�������Li���;�IԐ8E�H�!n�0���$���2b��Tj���i���ۭ7�Mr�\HǤ�Ԩ�m_\�H>(n/��ײ�[�]�gyu�W����[�k�}Ѫ�@�����ǃ�u�D��Ky�#�t�����tJ�,O�)r��C�ӈ��b+0��'�}0�������0$��[����N���~��q�%(�����S���H�9�e��nSB{�FN:���X�)]�h����#��fsu4믏���Un�1*u>^�\�7�U�:de�Қ�<����t��E}�B8��#�+���Ѹ���a�e�����⤸:�����-�<��M�&u8��thcr0�*��.trK%S����E6�c�i�K	I$�ċW�Ƅ�|!�ّ�v�t4��>\v1��z��K��Q��Ϻ�Q�&5��+�r����R�J�	�F##ڨHL�rM��̯���x�1;������|���E�T�I�<����Љ�iT��9�I��E?�Pw��7 33W)���m�]���=5�5�$%���<L��"���䞯�8�bO�X����<^��/bc�x��}�+exB��1��wh+�j��A��y(A�ׁt�;�Fm�����$�5U7�#*Hد�>e2)ߧ ^
�O9�u�9:���e0�^S�W"O)��ױ��9fEo���.P��"�nd#�?/�tJ^��iM\���{��j��;'<����Ye5P�z^���r���jN�umj�:�ni��g��}��vKq�\w�u;���Uo�t�b1."�[ƨ��u�x�ܢ�B�F�Y�Z�.A�pYʘέ��+�&���tdu��)�::3��
�+/��ƴ���	�+K�"ŉ���o>�r�qӿ����5�ߴ�C	��;��m�6э��?3��di�:ş�MCW8J�m�U����ӣ�Pm]o�%>(��X�����%`��
&��s�j��m}p8=9�
�������	�5:A��A��F�@��i���l7?m>��默�Zoʄ���,���[�c�$?�n���/�>Lr���yʂ��dHީgyX]R���bt�s�hS�Ғ��/�j_>��[wx�N��Xܥ����%��y�v'�T/�qVmW0�2Y1<�qCS>�m+�pvS����h�/g^��S	&Ʋ�r�eJcb���o޻'��qٽ:��Gs�o	��)ꂺ�y�'��3�E�bt\�U�Ds� �N3U}3��E2�����qP̲w��~�ِ�k��}�s'/C�󙓆����ڐ+�b��!I�dO�m��ws{�Z�pE�@B�'%��㞫d����+Y򡮴Ū���C������$N*	�ɾX�G�O�r�(����gV�&[�����a[@��EPށ�g�S'�
N�&�B����޽+<��.o!�K����Pɝ�4�2�T�m9�X�;�&��+���n�4	������ơ���l�Ǖ|ܗYܟ�E���h�m&�M�E\4�f��n@��2\�ڛaE%"�uI͑��B�4A�ܩڜ��ٟ�y=��d����I��9�3c�3%C׻��r���9Zď	n|A�M�V�"�q��4aד6����"OH7D�V����X̌;��&N�q�]����țyD�26�=�'6�G�e�[ڐLs>�D�����.h�+3k���CMH��߅��̜;|ĳ������+�Ѩb��E1'��i���*oی�_qd�TL#ߔq<�^
SY5�ϘҘ��u���غ[��×2�˖O׊i�b�of���[��T|�ž��R)�I���#lD<�R}|���PѮ�^��,���)��UL��.�n�j�QQ��/��%d�S�
Ȯ�.gّ��e�;��ph���?;�~`L��6M�Kmz��mt[[DY2."��!{5x���mMM>����\�O�h�/!��\_�R�է�c�;�� ��S'aR��o���5�+,:���D$'<
��b!�5;�ݚc�-���&(G<��2�!�,B�>�U�;��<��P;��<c}��C�^u��^9���M�b�[dn*-m�"ʺ�}���;�J����"��N�����%P����N��VM�V�=�Z�>ξ�[V�}�͵���:H��L� F�v�ۙ��St=���zm��}\�6��i�HQ/5�F �r���D�:�U��gz.�}�0iwd�%�f|�����xWtw��u�j����+ڔ�+�a�,i�l���y�hf��?2�Κ��ޙ���%Vsنǭ�[[ztշq�lX���r�P�Lεx���h��.�Z�~2��*�{w�.}�Y�Uf���_�x�c�t��&՜�_L�Lm1x�=�4��2�mW�7��{�aq��#���o��Rˌ�،�����)�Ô�W�ta}�mt�#�1�C�;�w����m=�S�i���0ܗ�w1,����j	��4'�xԡ|Ⅲo�ng�;����=�?Oz�o6Me+�z;l�	�/���뇯A�~7œ���?������n�d�p[��p�*���w�z6�|7��Mrv���>�G�:0��ꤱ�P'���֢W�S��#f`�{Aq�%��%�����ר�/5�3k�W4�z���~ۆ�WL�vs
>��x~��<��5�<cu��]օ5����m���s�Ƨ9(1k/�謪ciek]�S����nT=�n��cX`:�mti׽*��������f��Z���LIǱ�):/������M�E[���2��%9�V'�����gf�����Z���F�U'�J}����LW�k0���e{l�d�^��g���IkٱT��z1kut�����ٴ{of�g9&L��t4g-�w*^����s���|5on���\�'�z7�љS$��ܮ��Nʉ��h�z�"j��y�����?3l����W�>Y�Ix�8G2�As�:D�c�,Ry����۴.�1onqdu^�;<�f,5m���w*�>G�����U�S[f@��,�>�Q�U���t}ԧ'����]݇�%u���#���C,��~c:G��!��σQ�ý��A�x�GM��˯��Q��l<�46�e��fA���s���i+�R��.��W|fU�E�'(���ycKd޸wm��a�ӓq�]vO��w�?qQ��z<65U{��[�s(��Ǻ���6�i]9�ިf*�Y�����>~v`��	��h� tq�c�r�򾰴�C􆾶i���suY�g��e�g����b� Y�=��ͧQ�I�9���f��L6���[umz���Ca���w��R,\������&b���Y��yon��7�<E�m������;�,t@��\�g^]fMϕMJ
����=��=Bwf�7��u�R�܆�l4Tb�c�2�qpX����]��7|���r�6鱍q"��.��7��mm�(m2�ޔ�Y��Һ���CX�θ��B�3ʧM�:��wm^9�1O����M�mɹ��n�&+'4}�w�o�I���ЎtL=��c8��<3�઱z̳K�s�eU�:��wLM��æ�ܥ��0O�Qhyu�#,��-أْ�N;FaՄ���c����W5U5��.�0��iI��r���[��]Ľ�l����������Ͻ ��dԀ_9�^��W�R���i�c[�/�Wg��{n�������eQ�o�3��:B��C�mi��
L�@�N��6��_^�����xJEf�*���yxƥ�!�lr��m����[Zx}2�֏�y��߄�]kx�yH�c��%v�G6���j,3�5귗F�㍙��~�Y;lm��sڽ�M�G�˶�%�i%���9J9�a}̟]�7R��ȷ��aκ<o#�֪g��z*�jK�.}�(�շ�)���-lX�wl)��3�YoO����zg%(��� 0��,��C��1>Ͱ K�����K���r�ֲ�|�E{u`�Qf[VoYz.�q;e�b�\�Bp8õ���)޺ޘSQe��j�M�Y�P����b[����(�e��T�
��7���dV�y����[ڔ[o�Q��T�D�RK,�>�1ا{��n�G�j�K��gu�N�RC��@�Z��e�G����*����z#͘��wS�T���cp��D����um0���9lzTO1w4F����\��yS�(�$�U���g-p���b���x㬼�/���p��u�*�+�yw�krkMf-���.��S3g^�KNN����[�*�L�J���c�SE�R�x��k�6n��e�YPk{Dwe�l��+h�V�fŰ�Y��j�eu���*�DuZ�^4���YQ�!�*��	�)�A��0����״9v06�Oj�k���h�ɚ�Ʋ:�7I�^Ws�x�Ǌ�9ln�"��Y:��R��t$Rh��5���5ʱn�Wyy�'(�؄��ow�.�=����ԯ{q��$n�0ɓY�2K�X�Σ�.Ѵ�%�<������s�4�t�A�:?�3��&MC��u;VP�MfD9�e��t�sy�qj/1�YY��]��UKM%ǠB'XE� �9t����+	��vf+7}C����:�v��^VVqP�R�
qҟ;Z���sW!�3��vc��V��)GC�n�!m�M$��ά�K5)���r��h��jkM�g�mDK,��xd7�5x�аE�����.I�,:���Mܩ�2����4���m�9��(�dcP�����d��S8V]�xb��&�#A�.�N�.x�Z�Kz�����.�R����1��k�`�{�����v�]1��<�λ��U/�R�"z����jR�r��X����,N�KA�Dv�Ԥu2������b�S��G2�WC��U��RhT�Y����K�����\�v�F�ulq>�{�M+7i��v�++Cȳ_r�Yn�8V�ъ(����S�'�Xsf1ȧ��W]�qR�|6��b�:4ՎS��ʂ�tf���m����{]�ĵ��L�m'"�W����9`A�׊Ԉ��0M3H`� ��:��k[@�V0�_c���em:����7�����{mp�9�T4VN���o�b5F<9{|�e���W<��)���)r{���K�	`d�������K��+k��ûu���pK�r\v�;�:��p\D�3(�ӽާ��u4��kp��p����n΋ۭi�$����Z�7\���$D�K��ѣ#�bR�z/��f��Ѣ��H�ͻ��]EQ�yӰC���>Pwil��n�uK���`h��>��K10~V�V��4�"-�����A�(�W۠��G��z���B�gÌ����P���:�p+���!e�Kq�j��Ӭ���M|Ȩ�ځT͹j�M�0~�N��]m��u�7�r�m�l˗�Ҹ��3W�����MėV�w���� M�J�!�7G3lS$�ټ�A7+' �t�#�����3�ݠ���R�յ��rۡ����jj�Օ���m��g�빺�%6����핳��ګ�W�qY�^�t�m%2��ӻ=��ج�3ݞYMT�V�b��M����
:t�Z�m[U��)��X��n��ڲ��{�56���ɫj5��(�n�>�Gŷ�x�I"��aF��QZ��/}��[n�o.�V���ʪ��+��;/ޘ�M۝2d�ع3E)]�Ȃ�B���.2������zwA�T�K杨fDW �����S%�c�~��"�.��~���5n����-�y�̷�Dj5镯�L%��׷a]M��A����U;�ԁ�z����׏�ǃ�v��ؔ�}=3U�1$�U�|�Z��d{5����������|}��~���ˍpȹP0f��3������kre���;c���[�6�0JK�Nv���S4�t+{V�܀OϘ6]�VM�=#14wƼˆj	�ý0�f^�1UG�ӣ;�wZ����|"l�����47��)��7�[$D���=M:{m�L����ϔ�T��i���Ua��5���`m��q�Fُ�y���\�+�K�j��aǉ��/wʚ�Z�"�ML��m�(O?+�W7���ib���Z��,��fUb�xl�Z�u,}Ȍv\V[v��;����3-�y����G* �*�R�-��4�d�S�%X�!mS�qune�&�c�N�3�j��V��P�U���!7	�8��wM��_���m�*Ww���j�i}֯%
�i�H�*D�2��q�6|Y�A�x��EXI���X*�e1-�����Z͆0�S.����ח����,�QVQ���PO����B����]�Σ��k����0u�-�v�K�I*Z���K�j���Z��?4c^�vvݴ�U�k��[f;7˰�_u�l4. ��.��6b��a*���k�ά�Ɛ�R"���h͑���5ӷ�
~S%�T�L��353���'l���*�� �
U��~!������f�y�u";W3�יoSݻ��Iw+O�cKd�Y͟�Z4����`����YZ�U��ʈ:�5���N��<� ڈ�FvI�~�avLUZ	��6�)���''Z�_�ܜv,�Q����X�یs���gr{��h���wM~�xr+�%<�Yb���+6,�b�݅�JF���aR���W%�y�Ч��T��nB�d��w���ʗ��!T~A�V;V�74f�F�e޹;��lm�Gݵ�B�/�j0_;��&�U��Ng/'�4(��W���G��W�q�.��.`eK^xi�v�����2��bݵ2��4�i�ْ�Z�;�2PE�F�'Y�ia�)��=+"ҝ[e)��e��-�6�x�Wm�3�qrV�̧z�8^�*�ڣ�9���g���J9�n<c�.,����t�*S�(8�f7�0`���F{Y縑���Ϋf�#L�å�Hx��Y��_'�h"#����zMɝ�yy�V��M�� �2AU7X���m��-f^�E�D�mG/o����fHr�r�\f�iv���j�W9I,۱�ג����.ݕ�y�mk��l��̀�W/��!�)��}Ѳr��d��r#�t� ������[���Z�w��2&񺥓馼�)�rÍ���Б����3��]�hx�y��7�qws�{��P�[$ى;���~r��["�?�3������Uo	K�NU���'o;���2�l�>�oLRr:��υ�k���ѹ�T��hvY!���1��G���葽G��]��>삍��l���{�i@����3yu6���L=��#��2�͕ل���b�%�s�+hk��m��˪�ZTCU��[�m����LGX��Tr+o2�[�u�g�	"%BfLoX��T��kT�>����/%­�4�+@�7���ݶ�u��uϰqXKƁ˝բk(}�+5uM��NV�!}���mV�3��ob۫���)��;���.��4�# l(�R�XK.�题ڴi-�!P�b��W��5�:7o�cz�q�/�l�ݿ�$���a����x���W\ua6��l�����g�8��|��B)��f���³6p��]Y�dN^��6s�Hk��8���Uh�G���l2c�I�F�H���u7J����=Zn�U���l�����|č���W
���e�G�Y�3�Yz�BS��i�=�����6��y9^ԛ���<�!l��QZ��~IH��R���:*��O76e��f&�W��|zbmrO<��u�t]������ݹ{7*1Qxx^���<2���ǃr�{5t'��UV�bK������\�K���]���3�}�߷c��<��pk��Z�"��;<aZ��g�a��]�ڇsNo�k��Kr�«�4��# 5�6�0Sd�#�C�[�:�C���|�vE�[s�9���R�kkdR���,Ȑ��bF$����A�*�/������c��8#GI��(�WB�bo8��=S�'�9�1v���m9����҃��0+r��=E�A�\oR�y�kmq�>��[��3�7K�n�jY7v��lswp��x�n�s�4��P����
�m@�}�R�p�����\�T���R����{���(�t�1��J��#�Pn�)S'�l}����P�;�w��=7
:˶�%��"�������mlMB�4��.���\fj��a��r�Ը�޴�tO=t�\'�����f���_m�!�)����3�z�>􈂍zOG����%(Ɇ�
	�k��^��&w/_�y������XG8����+H-Z��7���ͮ��ɮ��W����k����]���w�5�n,1%�#p�2 ���R;[�`mI���;���\r�A%�`ɞy��q�#(�ũ�0��st^Fu��Щ.��w�mŔ/�n-�~:����q�U"��a�0�H�nMl�~>F��bN��6V���OC�C.F�@�wEA�C8��}�1i�F�g����!���*bl��������3 \�p��l	�\�V��w�))|D��B"����+��ǒ#��<kiņ�.fZܐwd�{���Y�y"��"��k�U�-�_Jc%N������Vm:�*.�_me+��c��EvyZ�ɪF�&c�u����\�t4��3������~�.g2���l6�a/;�:��NLUd�N�D[�iX��y��c�oi������ɡ��eߊ��}ҽ�:�W���l5�Pp^[�����e�+	sY�(�|/C�ZU��Ŏ�V�e��­V��;�A�;�&;.w�*;[$5��8��'��%�����ȣV��fD�L@�UM���1\�-o͇;y��b���>�ǫu�i}K���J��-�	V���BKs@gWq�}��3,�:�$t��Ŷ}�,�]�q}�nZ���
��̯�V�D���HI_(%�vW;�v[~��g�Z6ӛw:������=��~Iǹ�,����=�t���Q���6��L������"�D{J�K�W>;}��^���U��mm�K<;�bs�-����>����a�c-0��Ԣ�t������W�N�oVrՖu�}֞���"X�:����غ�=�NI'Xw�&:L���|����{�.D�r��e�m�8�o#��+�%��5���5K�ZJב���ljc{�u��1�d�a<�S>�9	4�[t�'j�
O��NX"�ع������NWT�`O5P�Udl��Pa��Y�7gK���,:�춓}�o7�0���@e�"Z�r�|/hĎ�[^�ۍ@�>H3;W��R-�[7g��������c�Dn��lY��O=�Q�X���Tl�H�T��e���]:������`��!Y�8U{w��֜O�� Jɓ�3��i��E��5��2���ϔ�����Ma� Ȼ�jxpq�y��å��R+��j!�"�HW:��4�<;;����|d�t��]�fD������齴#V]Y�U�&Mx�'�!�LU�R+��Us�k�Z�G�����wp��� 7u7B��F'&�k����@��+(�r�W��TͶ1f�c�˽Ehg���3:���dS�Ħ�������O�����N�s���ލ|5't�i��]��d�{B��4�~��f�8�Zk�"LgU��ޝƼ��u��������֛��M�H;�t�<�3\�ǫ� `�?2��������vs<�x��ҁg?��!S��dw��t��M�-����7
R7ĸ�M���Үw�,	t(΂w錻ۦ��	��S�QC��.���r�ΙB�󂔝��/fg}�q�cRQ�ȭƎ�jb:���Z�^�rM�{M7$U���|����}�E� �fC>y��V~A����T�%D˽=�%�T��h��Ҹ��S�ս��l�c��wn��%8+�A��� C�O�7��6�ʮ�c��uJ�q��mo��P����k���n��N;G�������F��G�'M�*ȵ��
;���=[�Q�my��6ZfH���A���!���0{{%GG�=�"<��y�+S�=Oh�:�b5�1���-����@Vf��R�MCͽ��Sۚ��;_�fām�o7��gC!��T2�s#���M�eO��@
=�:y���{��������*��~�����VS��g�~d(
���ٟh���+���GS��O�=�^fR���C�B �D��Ϩ��m����8t�&�A�騴�D�^�Ú�Z$�0�p/Y�I��l���m��Ɩ,�J��m�k�v=;[l����^_+oG�dv㉈B.�j�����^�ᬱ�=�^Ka��_'p|NӤ�W1V��&�9C5�M�fh�v-FƝ�޽��D+���([�h��� N�ŧ�
̗q����E�v�P�λ/L�����\25!��ק� ������e��ڈ�ɡ�{�v*��=s�z�-�|-���t��§Ȩ��흢�O7���V�,P���ﴂQ]`b�Բ�(yXm���Hk��m�ٵݭ�b�P����źo=�����z��ܼ����r���0[09,l6Fc�np�+[D��x�i1���X۾MC�2^V-���.���(ɼ��l-���3�ɨ�3�VY���Qú��A��Iq����#0��ΚV����^�gR7m�d�ss�W���V����`-�UZ�bv]��o"5���U����/���6��fk��C��tAF/���i|j3��\wd���ѹ��Sw�G��Ƴ��un�}����Z-�}DT5���dv]�H����{��e�{0a�Gr�40c��V_���d&����U��[�ˊ�&V�J��oW"��,Ut0u�Q|Ґ�3y-T��㵝M8,C�A��XzW'�@}����"^�c=P���gv� ��Jw+�n�l�&ɽ���z�-�I$���b���A�pr�Ggk��NbͰV��DS��N�JQ͸�����{����3���9)��twC5o����C������~�ژO���N=_??{��P=ǻ�[e�s���F{v?n�1�i��)['��P�4N��l_nA�F��P,tC����б{3��)�D`&i�ٞ�k�9ls���h���j����Cj�<d5�>�*bl���|��``F���|s�Ѭ*eo�p��偽�$k1�<�v�{��X-�H�Q������P���"]��2��ӵ}>�)u�����g���/wʳ@�ܴ G]�f�f�o�l�+��ݪ|.3��o ��ꣷ���j�ڴU�&�Ku��_��fc�7���G����C����c�q���*\sgc�k�Q�D����FF��a�W�����>�m�a<'�O=rGAxE#+5��g�oke�7o*����=/W2���"8-����@�(� �� 4@�Y���-�P���n��_��d�Nn�C�"�{�������JӢ���HX;X:ѕ�o�����SY��AkS� W)2�e�j�(�N�E��X��W�z��3Q�`Ȱr�sP�X�%�*W+�����D��MU�K�1-? #�z�#\x �������G݋��F�yx)汰ճ��}�J�T�ie^�bYxR{GvWK�#�
�_�i�'������s.�SŶ�p�j,�v!��g!\n7ӄ���[r΅qj�g��5��sZ�7J�gB6B3Kԁ�{fW�D��ǌ�;���'L����aWrΖ�=Z�����4Eس�4N6��r�ާ{z��E�Ϻ�B1�\kC�&�wZ��}��|�Qʂ��wq���	��`r!�g���Ꙧ��[h�nK5zgtx�J�@�&A���e�U��j��z�����9�k2@ר.�wB�7q�����[t�*�(�4t�$x�hM�\I'��@��#�Xܮ9��s��#�;12�6]�L�sf�K�������>�1���Q��EAy;�]F��]]j������^�������3���Z��ý[�G]{���G9fbڽ�j�B�jU�-�؇=\���i����xc>^�t�����7�"���3뢖��!-硬M�,��G-�V�N45h�E�)���	��Xz-�����J^.kN�q]gU㮽�:�oE̉��9�j���5�Gx��~����/;�g�dh+4�a�N��,��ok.��2�!@�֪�C����1��yJ�ݮ-�  iǻρ����\�M�ܭ�s��<{'c�$o[aPc��[�^�8.�P�z�U���s�< �F�5�uu k�+�C#[ r��e�P�*W7;f�\��
��q�R��xD��]i�I�IX�9G��>Υ$v g�s��݆�uQ�[i[ʼr�<�tV'Hς�W{
&Ơp�,0��v��cu��l��RgS�4
(�h��T��5��gS9t��&r���֖�z��o��[|��XQSz�[x'6T=1�e����9�)�pҲ�3���y0հhj{E�|�	�$n�-��[��@�'�6þw�X�xèž�ז�19g��f�x�ʰ��j�o ������ft�yS��ݼ���
��Su{�P���5t�hg6u�Q�ԗ5륪�QL4�i����D��MA�pK2��`���,�W�9]G+��꺂V��s���GbVX婎��ɹ���Z��̈LОl: �ޭ�����IÎ��5�@��d����2���t���r���}���0�C9�-v�Yr�[�Rb���ݺ��*sB%�śl�����tL��;ԺG��|;3z��+�ˏK3��3Ύj���J�f�Y|�� �����0��Fܣq@AcSS���W�d����S(Q�U�}���jڶ�QX���Y��+/�ܳV��S^w��H�Jիg���M�w2�V(�\��V�QJj2�!,V�6:(��i5*��~/}�ER��Z�[�s�ݪ�Su�Q))[U�*SZZ�ǫtws��jjVT�󳒵)TSS)JQ�/Vy�Lꚵj|ۢ�����UemD�JUZiQ����'Z��m]m�K��%UK��ZN��IV�K���)5s�]��t��v�պ���ջ���TZ�Wr���u���j��]�V��YZ���J��[����|���P�T(W���{��Բ��kT\=�F^�[Ѿ�4�����%E0Ҳ�:4b���E$v%��ϧe
ۺ�]"lv��\���9q�p��(|�"	� " 9V
�u�i"�À�@��[c��W���]�Iv�C�X3Α��uo<����6T�׻�*(���of�R#��
�>e�M�ݓ���3�۾ZlC�#R-ġ1��X�V�<�|�'�/��0�Uv(�uI�kpfM���l���IlF���?f��T6eq~�-�dDiU靍�޻�-Y@Yֹ�O\cp�LV��Φ][��w�Ӟ�!��n-�.:�\��Ӵ��s�e7�4sjZ�Pt;vw]si��Kz�����q�ȗ�9��0a��y����selHn�g,����:6$��G��2��:\c�E�YseX�.%���n:eX��ֻ���]=Tw[)�v�$i��2�lX���Њ��m�".jVt�̮L4`���Ģwv_JgGG!�+�����.vM��E�Pw�:c��s[*+Z��_�!���t,�i���C�"��T�~.C� T<ݤ{�A��LZܘ��S��c�z������ބ8��i�ã�np���ܺ���?3>�IlJ�W睸����S�}��fӡ��!j]��Ϋ�bY|�׹'%�c��%����ǽЗ.��y)2�.��Ϛ��8��n�=��
��+fȇgf�w���ø��l���L��&����yXy��5s�/rm>�%�oFP��9]�S�{��,�m�)1�wa�v���V���W@M��7Z�'���')��z��h�ʶ���*�=�n�{L����W�Y�W��d�4.k���s}��{h���VI�[\�"Aݩ��k�!m�.X����3r�YVv���|k����%A��W�����V�(ocÌS���ngjֵ���n�1����@V]�m�oJ�a�K�Go#E���Q�˽�u'nsZb�V�ܓ�+���o�iUv�4�%�z�B�2F�U�rǶm�HƦ�7�����؀8oC�dN���U܊��̺��z���c�~��u��;�?ۊ�����lH8�q�r�od�B�쥂�1岳�M�WQ��ai}��y*=�[ߐ�6|�n��Y�Q��[�y���R�����ώS^������C ���U��=�*�]�1ϴ`�嵙��#�h�wF9X�,4���8(B}�ɵ�a�39G�s��oF9;n�E5v����q��+k�#)�Jd�,3�1Wm�
�J�l��V���-T)���s�M���uֱrɀN�N�#ޒ�-�w���o�����g�?W�`�-���q��u����۹S���pU2`�hV�j�8�Ca��dr�̪F�6�}Q[%U,5���qh��:��(�Sg�`ɁvZ3x��rHmt
��'����f'1����r6��l�������VӱY���m<��-��'3x�Xx'�}w�z!��V۲�M���CMf_�'&��%��\�C�WE��a>�[��ꛠ0ڥ�ϝ-�x]σ���!�J�le\D��9S�4��/��t�ܽIu�I]YU�8�}x˥��m,Y[t���qoj���:e�C����d�G	Ky���ʶ$U���OSo&��ެ5Z�[ͼ�}�6C�s95H��*�f�%t�9��Ժ��%��yǛ^*�ɬ��Lz�H�B�_�˶�%��"����+�B�d�%��J��R��V7���ӻ(T�,����>3fы[-)n���L��<�b�Y��$,1��㫩��%�S%�36��%�siE�v�;j��'/;; 90�<���2���M���2�m�oW3��c�o��J��o��Rn���w��M�^28Cl��;��#V�fɛU�z�X��5ag�����	.�U�φ�����J7b͟�d �=��^���&�n�DjwW�2��TA=�7e��;�--25n�F�y�?�K@e�=S�hݳJ��|��UW�D{�\qZ+����c�,����O2��g�ГYgM�+{��ѱ��ŷS���&<��F��6;Oci>�뢥�u�̒�jԣmw��?�h��ڙ_X����_j��>v͠�/צZy������nz:b/p�\55�Yl���qeH��n-�)�w��6���cz{��آ0��m5e�]���ܪ�~�nyM��͓^���R�8[��
Ө���\-�h���e���C)��[Raq,�Ə^�f��3��<���	�V���Khs��� [���>����q�|z�WJ�_��X\s]�1'��3 %��7X�2Wa��w����]�z]�V��4��x�^[�ȗ���K�Ns�.���E�D��va�Uw\Ď�O\�Q���oN���Qw�5��5yf�Z��7�X�˹w�3��emڼǵk� �s��Wڝ�𱕬M���ή���ґP[�g�K��]N�T�a��YC�
|)B�Y|��Z���n�Ƶ�F�;�������'�����s條�,��ޖ�w��6Cz�����I����~���LN,<�
\�P8����h�mK����o�8���[bWGyi�Wy�����%�����_,�𿌯�_�Џ?w��g�8��r�5'���2mX+��]�Kn��qf|�lp�N�`��0�u[��d�lY=���#����ϙ�Tq9�`2҅���f��nt�z�<*2��9��ݵ�>�):��~p��>�f�U��>����x'��s�����BK���Ϩ������ݪ�,��u� SLq��=%h��`�(Nf�l���F��C�	56��f�V��ܯ{�٩��m��k2^��^�(�r��T���xQ�;pș���5�nEف����9'��1����0<��$<��9O4�ݽ�P�(�|r�W�����e����^~u~k�%��}�v�&�lגL���7�p�ֽ��1n�y�rSWs�S��N�� ���߅�Y�ԮNV)��;�ǯs��k���u����b!g7�#r�3�A���B�0�l����������Ng��z�X�q;|7[��E*��ƙN�[�\�R��}oc/uF�+��]�pQw��J ��y�2D^xi
�l��0�}�˺������'w�_�b��d���V�n>ӈ�
(�R�3��4���,��EO�Z�E�+ �pT�jR� �M���K;�}jV0xb_jp�c�.t�oK�?N�i���w�jc�}��@��������w~%UJz]j��kx��#�+�3v��*�x�[-����[��=\�|���׸�=5���&f�Q�h���H���t��^Aݜ��k�'��F�^�d�J�ɻ����3���䑿2�o�j�������c��0d����C5Yo�s���%ᣕL(��m�X��6����^�
���|3�/`�\ѭG$�_]DJK�����9�X�j��֎��&��ӆ���x2�.�Tb�D;���ޛ�G+r�� _D��O33�=[k��%�Yut���#7,sފl�{2k8-��m�yZd�>mn�۬���̘z���"�V�@�����g&�]$���ӯ���|��~�n<�c�D9��ȸ�m*�ۤ�z�)	n���O�B�<�����z[/#���ZYO���͸���B'��Mg"���,�M��LmtUkb3-$�W@��M����3�⺀��rY<��M4c��^s��z��� ��:���}�B�JX��ja����y�qL\�沌7g���V���<��,��H�t��o`ْ���c��ꌫ�PFx,�4.��{�ˍ̘�+|2ё�u��- B#m r�B�>������<�G$� N�@���uc.��#Q#E�9v�)߻`+���6�g�"�n�Y�L���`�xYOwUy�z�~�ʝ��
��H���b�����e?Q*r�۴i����,1T��G�L�Ml^�����;W����v�	�^E�8�������t�Ľ<y��KT�q�c^��sXY�9Y�U�x��+k�:�[b��D+����F��;�
���7k]�R�x.]�n����y����<�������X���`{>U����Ee*j�etc;��s�o7O8���u�,�;h��l~���乻N~��R��^57�8�ot���CT���S�m�(�[V�b��c�����gUy��zJ\mml�U|���I�ivY���m���dS^��l�;C��- �F��T���O�x�����1B�*�����=��cj��]:�=C�v�H�P,�Ff�_oS�;�Xx�	UR
Qd����h���>'�Q��7&�����{�[SN��p�fFe�O��i��f&����@,D��~�M���3����Y���ڍS�TEu7E��Ӌq*��K����뼕�-�Aa��v��ӳ��.e0�X��_n��ʂ"4�G@��T7��(�r��=9ܭ����r�X��jg;��,:Ӎ��e$��[���@㧏����~�;\����L�R��FɏK�vFl�VpX����}��z��8�N�;�9�����P*yAL.x�GQ��e��Ś��[��t��fe%��:��N���+g�4fuç,繰�_�I��Z����{�큾G/ܻܥl����L�r���F!9Fݍ�$�B��x����:��Ew�3�R[�;�N���0�n���e��	������p����=�5��_��!a���X�������42�o�_�.ͯf��9�wg�P��e�e���Wu�EH6m�[��h�9��D_T��b_6y�M�0�f���P�>���E��&������؃q���1r�\�ue�YSwՆш�W!�\�)~Σޒ�&��r�,k���{�(,����NYF*,�t,��I�`&��.�eN�ۓ��j۾ڛIp��>.�9My�i@�� >��.�p*R�ӻ�Fb�F���lד{��Ϙ}}V�%o����"�MLkyW�}��[�hC�^�|c1�f:�����D�v��+�M��ژ�S7�j��x���{�Y}�wqp2�퇪W��6����O7�S��@�b:t5��ݙz�pZ16�c<�=�b��L�B��P�7YZ�y�[�i ê�˨�'�����M�v��'*�%�_]�1 9���v�YCi���q}3reg+���F�C��e]7��rT�}��'(t�8H��'�Y�44t�"�ok9GO����qk� 
�Pei��)��{�k�T���e�e�&&��i�4#��}I�{��W��LF��"6 �S:�zx�\�9fԄ5ފzxiv��2N����Mּ��ä]�,�����W�?%���im��~�R�ɐ��i ��j�u��`��ϣ��/�n�F�o���׺%v���v�uY٧��U�G_$��{���]���d@XnҞ���iͺx��X5�2�?.��:ZAF�A�����gc�A�*Ҧ�!�� ���f�U��ן�Cp���h��v�"�JX�)�lR<񜞔�U)�� �7j�c��t��;V������,�x�+���e�U�_	�]�$qi�;�Ch������Ǣ�Ջ:�)4,�^|� ��w�$�C�WT�̛�oXȄ�� 2ײ�቙z�Y~��o;�^Z��]2|�Q��Z�n����f�����z>�����i��T���5�&W(���#�`` @  j*w�M)��8\���i�pY�bܶ�Ҁ�M���o�Fq�k^mnd�Nr���د);�)�n�6�b�G*B"�'��J7E5��0�]tuz�3��eA�n�O��Pۈi@�֮;�0�A�K����!��t�H�j(Ev�`�[�+φ5��U��F�#�+$�fQ%E�������y�v,�ä��
:��l��/�#L[��X��aui��A�����']n��L����0�t��l����p@���Wf�\����Yn�
]|�!)-�}Nm�b��L&�J���+
(>�K�k�k{.=I�*cۥ*���Mʺ/w.��r��ۅ1��Kv&�/oL��oykY4^��>B.�oZ=zL����4�s�5��
Z��83��2��uϡ��)xd�T2��"�L�2�U�ֺ�C�%�e,Qt���7e���������.��g'w�T��͊_͹�ŃY���>�s�6`�*^��+kz�.�}�*qh%$��
_�n�y�M�5Ǧ��N�>֝���a�Y��T�b�"��vA�o `nugR��Q�WH8�V&'mnP�R�>�Y�Ōm�XՃGMm@T2�{W�$���l�.+�rk$��+.���v�I㘪��ƕ���Q��oA�1�V6��̬T魺�j�T�0�s��o��YX��������;�@�E��8��d���UԢQ�xt�dro{
K�C^a���օWZ�֒4�j�i	�C2R@j���TQP볹�)��ٍ�$��qP�	���_Ӏ���T�+R�ݤ��|��n��x�$ԡ�[S�F`SoVk��:7W���y�Y'1�ܼ�� ĝG])�]|�ˀ��R�O� �X�J���E��o���O��s��.���U��-W'�E���w��y��a���-�Q3���´�;L*�n^�#lZq�����v���φ�������Ѭ�*$�V�*��ʠ�cx���ҟs`�;VԚ��əZ�2���;�,��1E��s~;x�9v_Lꩫ�me*F�{���aI�9�:d^�e���&�h�K�U�V-��s� ��>��|�L糒v��:�.
�v�[�vJ�*ڭ��۵�gQؚ�(ڮ��q���̾.d��Y�1��c�����k*U��19����J>u���K0f27
��tm̀.��5M}�8X��E�Y����W+g��[�sʜK*<�}��4۩��0��q����t�EQ6Ȱ����ms���J6a�BU�Ҕ��;����.cۜ��[��xr�y���o^-,���f��,��Cc��uC-2 �2�Rʥ/j��v�nt�j>�}�� �K�e�Ź�FP��Cdj=��]n� �\�2^�֒/��*�|n�Ӭ?a��9݆j���p��i3���}v��&���
*��j�p<�eL��f�g@ں�Q˩n�O:3'@��)L���ު�P-ݻB����5U-U�%ԥJ�T�E�ҪɪX��v�-�J��V�������*H�VR�iVV(���YZ�J�h�jb�Z��W�v�kTR)JUT�㬵J�i�J{��V�<��j��+-m�R�R��Z֔Qb���Z�V�QIIKK�U�u+I[ZR��%-)U�m|��Ej�Y,�ժJ�-T�j���*ڥU��)Z�����R���VV�U�,��ԪT�,���ZK�E+e������j����^���YK+V�%eeR��*��ݥR%�EjթIZ��ISIZV҉)�L� ��Ď�I�]0�^E;���bț���-�z.���Qvn��v�Q�ٽq%���D�����Gv�qxU]'XiG4i-{q%'��{��{;?��U�����n1�Mw�)�o4�6�"b�9ѻ��(�R;��^�)oQ��r�G+|�
/�-�����r���.Z�w��2^�$^��7R�nI �f�vm�O�'�H�i�����e��=�i�����s%H������H��� �Z��_�g��:sg���^J'}��x8���O��3r�:}�D.3q���S#�Eګ~
Ն��9��׻�����2����(�C٭~�%�޷Ʒ3}'750z��m�՚��ej�Ǜ��ւs��[l��ހ���s��g��NN%-���7L�{�l��3�<w,q�}aiؑ
:R���|�
YA��{����m�y��Q�&j�5�= ��;%���z�)<�Y�56��g��6�xwS�v��mN��o�E
F@�����4��JD��l���| �HҚ�̓ĜL'���*>^{�wOH����ݔ"�d��ءt����ʅ��iT[F{���{������Vڂ����5�%��oi-;'��6Z�a�U|��%�c6ЪU�X�ſf�v��+)�--�e���J9������v��~�������&V }�?w�}��Z����;!�H��R��n��Qc�s=�Ur:��N3�C��f�S]u�z�(ح�ץ�LĪ���	eG��V��Fс�'��؇�[3��sί���}�*l��/��wێ�G�SYA=��S�㶪��g���j��s)�k�.�[^a��R�w	����7\�V�f����]S��U���g����zsf�;���4F�u���FM�}����I�s�d�����)U���swu�˳0�u٦rr8ʧ͙Ų}	l�6����F�Δ�8s�qƪ����;�q8�d3���Q)��u������}M�˶�%<(u��Х�\cꃳ�"-�_wu��6I���Dҕ'��O�h�g1�u���ޡ�k�d�1���^\nV;t��5��q�w�:�$J�������J��І3c�1�r�Ir5�?
�{S30A
Z+�5��՜N𺇮Sr�[א�d�����A�Z�%�_EN�5�E���������y�<�⮕�������pѼZ�`��vf։�i@�u��<�r�Yk��s{��,=��#14��q�������劌t���X�B��ȭ����M�B�s��J:�1�wVX���C�㏂XM�W)v��o�܍�rd������o���/t��No+rv^�twq
���7���6�hj�F�H�Q�Փ�����w�ˁ;��uΈ5��vim�*w�A�F��>q��ǟl�fE���[>��<P�ot���*��[�t�kr��=�!׋�l���I�*�������TDD��LՉ{���t��n'k��q�ҍ�������a1�+��ܳ����fY1Wxs!�Q��Hl�Z�-�c����l20*ꌞ��A7����(�s�'f����Ҧz��R�\�j�����nޜw�h�1��8�{zE�o���j�s�^bT�a�ݲ�� J��M��ܙ�t�im������5�d�@���Tu��܁�۫q5��ޮ2�܍ťo�h3�z���YT��;w�&a��*O�N�-v��G�����[���L|�����;�S6���YK�KX�+7�C[h��ʽ�<Y�RL�����p�K+o:��cfq7]��r¬��Q�;�zGGϳ�a˓Uj:s��v���9�|$�̈����&mH*�/;2�"9-��;KK抳�
OoR�=�����-�	VҬ�w]��{�)��,ʘ̙om�r�����o�@%�Џ\�1�h��)_R��_�V�g��$��̖�cٺ��8�O^#����ַ7�T@+�XN�f��|3usJ��"�4���ñ�7�r�!oT��ٙk���In�J73�j�鍶���k���F�=/��.c��5*����w�\��9�fբ�̜i��񹳹���~��>wU��̀�o51F}fnTli�o�Y�]-�T��)��O��Gt+��f"�q��}��ݗt�#0�W�hwby��O7���u�i��;RB�jHʊS�z���.1�dݑ͕1P��8���[�G۟P�l��^@�m�O^x ~��L�a�a�ϓ�}��9蟤�]}�n�Vlf0�

����1�?���L��˝�}x�T�qǓ�6W��*�.�IS���F��Ww4v�����]��R״�B��w/���]��+L�U_��XJ��O��� �\�;�����p<���g���5�Ǡ��B����7�o����'�߉��a3�H�TZ���C��}��jC��T�Eb����Rws:@ժ��
B��r�����Ɗf��m�S)&��WS:�⩫�f
����
�K���e�Z�m��릾��~����3�\�V�UJ��S".��n���/�Ѝ�Y����r�v��N�"���'�̜�qV׊��c��(���]Y�{��,��̞��mx�r��&��Yi�x���yv`qF,���`�5պ��'#w-| n�ÒH���Ҳ��UN�][_4C����u�nS�k�2�a0*�v���}�+�)b}�u-5WH�����^�L����h�ɻ�u��\z�cm*��LEO3��b���m��:��GM���/��fM��|�H�3es靛����e��Ƽ����1
r]@�ɸ`�͟�ve<.���,,/�P��}^:��Ӳ��n0�u�����C��־���u���=���܆%7R���j_IΤ���ⴙ�{!��w<�K��Խ��Qm�C@������7-�����M��Dث�y�7�������@�3�py>r�*����;���C��o�L�kܾ�4��wRboOj�ygZ��>�=>���jasP̜�d���|�"�	��l���B["�l�Ǽz����Z4p��*leн����*����-:�{ @*
��	�hWaLoZA43Z�U\{r�*^W�F)g��z����7��}�D+3��X2�����ݵɐ~�K^a��"rZ��;���^a��#�h��8����֓����Ũ�g���q}��|l�i��#I��\�M���@�k2� 1U>{5��@�;�}+B�h��5���)��P/4�H�Stv�P[l�:[EPٍ��y��M���9V��5 ���[{��Rڵ)PYy%U�Y�[�Cc	�P%�l�sټ�ű@4q��e��kM�27��J\mmmD@�m��20��Q�f�ضtǼڹ�<�O^�\���&�"��]ڭl���um*wH� >���ZUs��q����sY�����s´����?��i�u�ݬ[�:l�ٸ@�W;�jf�_Uַ�Y���=`�A9
4B�7�+��'4����WA/�F�u���� ��M��Ow���D�_�z�'�m��e�\��m�s8�rFAxJ�#4#��Ѧ�!�T�MY��6sk�\OEG�����t�]e�{[��	�ܞ�;y[[}7ܰ�q^e+)`7g���1�ɹ �%�Ǜ�s�2o���;w�,�{_�7�����]�_�wb�ܔ�J������8#� ly�cͤ�W7G��z��F{7�'�%[۫,7�8��|v���Y�FW����W�=�u���Iغ����wC��H�{�\M\��t�T�l�忢�����f.@���C9L�̧ս~9a�,no#�a���]�M;�s�٘���wR�"�e£B����f���0�wA��*����d���;�(����Ȼ�7V�����w4ӓ��֋H�^}��@29>�(@�I���T;�7����׻�S�I�q�c1�S��>��b�;ME����X������b�l��m9ajV2e%z6��R�o9�aɤ�����!����T�� l������3������s�n
�M��;�WU;���r�|�Ɵ=(r�`ۮSz�<�����Z�6ѻ��'�-,`l �)�ћv�m�fs�}}�u|b�&$f��I!�j���=L�e��)�-vѨ�۳��Y�bc�����Jf�m�>ևF���*�+U��ʚ��hW����v]��r�H�����\��SD��]q@ȥ�M�빋c�wG$�h���n��z��Z��j;�Bo���d�q���qj�k b&8ì��yW�i��ގ�㓒8բ�⭔�dj��m����g��z���\���1��9��~J��%[�Y��$q��3�9��Wb�=����3۴&��Xi����uƆ9�� ]����Rݶa��vJ!�&+,�}���8���U������B�i��J��,YtOKdŘ����ޭfi��������U���r]�r�'.E����p;���r��#����<ǋ��D����w%x�Z�15f%��6�J8U�;Q&�'ӭ�[-�T��.���ub���n��x���s���Y��M�}/����򦳮����x'γiP ��1��ܢC�+n��{Sz�d{���ʽݢ^�N����ػan�/!��2e��V�<�Sԍ3�	���kvSo4y�/f.S�oTm>�8踞��O]l�y�Inղo_�F��}�[���Y�KV�D�}�6!n�M<q���v��[���>�	�3A���=��	��7��ٕɜ�I��Ջ�/���1#�~�T�n7�t�ƼH�R�1�V2��s/Y�ze��;z��������r�=�/9��H��i
�[�u4�V�����f=�ף��@jU1|�D�Le��	A�����L�E=�ض��m���rU@�Ll��/���5�q *�w�Z�\)L�S\�4�]n]����B� �����.���K]�T��Uqʸ�0�ܭ��sN���Gg�&�v�&��[E^U��W���f�	P�_C�ykU酖ƴ?�k�[�g��$���@���e�(yUي�{�q��Ct=S����Ψ���k���4@5��Ք�-���uve��ܺ$���J����f��œ��sǣ.joZM-]�^2ru�׵m�v4��1t�ǵ����ι���4�K�[e!��fX��W��+��9A��5bN��������7{;ܸd���#A������q]-�#ld��[A��3=Q��~����.��3i�2��|�9["�7
=�=>��t-1��G��G�d�b�{lFE��G藛�8W�����Y��]gh�\�q�iL�ι�Z�8ӱXI�x�������=
Ɩ��f�b��C�S[SLn��Md��3p��+s˙@U�t;�����`����p�u3A�BM8Ol�gflue9��P%?+{q�zV��Q֕1����;�Q��1'�n��X�b��|)$��.j�NSH�7>��j�c��t�5�M��u�;Vm�@1�2�`��e󄪅tu�#��u1��Becblh��)
z�sY�p������m3Q��ȅfDM��ˑ��� �=N�S��*HƉ����$ij8��c@al3���������~������������m�n����m�M�����pmX6�6����y��y���y޷�<a�;&�gM�n �-�"��m�L���c�l��LoV3n&�"ق-�"���,�m��M�LO��q E�D�D��<�������&�� �`"�m�XXyg0 E�D��,,;�< �6�E�DM��<���D�D�4M�CE��m�Y�M�y�Ǆ��&�&�&�-�[mmmmYʹC��9��{�������ٍ��)g��g}�����������ٟ��6�W�-���]�������������'�������/�d���~�F�.U�������/���[���������f�����y�����llͷ���Ksc��w����3�9��o�^��[��g���ٶ����~[6z߿;����4;������Ϲ�9�������oY���W�Y�foV�fm���	�X�m�&c,m`5�L 	��e�B�m�,C�m�� ��� kL0{i���m��ً��-&͞���ݳg�}���fj(l�����o[6~{~,�����?_�l���������~�/�;�6l��0m�n�}����v�^����;�s������o���>���m�~������������6f���l�v���������������m66f�����<�(�a��v[8����?���Ǚ�wy�}�������s�}��zg��m~{�l������l�~��53��}���?������?�>�o��.�?-��l�|~����D¶ڌQ�̦ځ[f�cS6�����(�+6°2����+6ئ�+1�3mX�C6�5�6�S6��LaC��P�[SP+6¶0��

cmA���`���
�
�(�ՙ��lVm�M�Vͅ3aY�m�l٩��
6S2��m���V�S
̣V�Q�6��CS5m�Q��Y�S(elj͔7��{6{ٲ��<��[~��{���ߵ�gٿ����W���m��φ�}�o���l�{ϝ��V������6�i��>�����?��������8����~�����3ߍ��������G�?vv��߳������PVI��J��׀RGw��X���y�l���^��� UPT�@J�Ҩ��J����Z�T*�"�E)�+Z֥A��i*��ݶ�5�U�TF͙��iK�4wq�%�,���T�0ɭ�Th�V��e�ְ@(�:�mX�e����k�DL�� ٙm��6fVU�h�֫m��6&��V�Y�Qi���6���򙶬�� =Vٯ\�m�s�m�:��5�6�Jiv�h[P�Nu�k���Vݢ�8����`Gs��U];%H��Gf�VF� ��(� � ������զ��ǦZrM�EqA*�����Vݺے�L��u]fvp�:���Ĳb���� �=z�n�s5�ӝ��R�;r\��`��J�5N��Ww:�۵4ήZ�b�-mZ�f� ��/��]�N5 ��ga�
��]*-����JYn�p�#�Q��ZY�m���j�x�y�q+�q[����Y��,*l��V��s���wMZDӵ�ئ]�3I�K6�����Z�[���r�KG9��ۙs��u�$�-$]��5e�3k�:�n�cLmZ��j�k6��g��j�B��)���t�[n��hTkMXZ*NΜ �Z���n� 5ֶز�h�UY�� n�
 vw: ���: ��p s�������p
���� ;U�(YţR�f�m����� 3�� �� ]� ڰ�s� ��� �  q
U;��P�@ 6�٬6ţVm�� ���^�e���΀۷��۸ tMY�H�� 6��@Xt j��      E? 2��j�C �ɀ	�h�S�R��ʁ�      Od�JT�� F&	� �@ɓO�4JU*0 L�  10 S�&�F��I�@ @   �I $&�2d&&��M�Ѧ4��RHZر���
��1�q���3&��J1 @��47vk^y�'�B$������r}� $�=��X�	HI�I d_����HIy����8���,�މ�?�;QF@$��Xs x��	$C �h��khR�1$ �@�'����|m��3�>_�_S���6M&���)�e_g����i�ӫ�7���_��C���c��q�����Z�mq��f�e���m5gU��� ��0Vn��-^2l�Q��T�W.���E�L��`����nlb�Lȭ��: �\�����<j6��սi�)HJ%��`c "�XɊ��x�<u����:�!n��Z��ۍj���Gk�i�M���')�u�g�h��1?�z��{�G���݌�l� �in�����EkÝ{MPZ��1��l��gv�ӹ��f���K6L�i��)LduNS�����͈�wI�t�Q��X��WX�R�Jش�?:�p��bnb(ZÎ�1Z4���*�@O6�O5���B��ȋ�bḏSX��cɃi����y�~�f���ʉ��_ n�mKj�֓���9Zh٨��+��K����yw4t�Mu,LjX���;��n��(lm*�z2�2��0��B7l����>J�T�!V��"��-�-���T՘!y��W�-�{��r�*;���J��J�D��ʲTi6���m��R��5�n�i�uS��KS7%��t�FC�nZ�wRn�N��PI�yʳZ�*��k����u�]aiۭ߉��2�ё}���Pf�V�Ad,�8mP�VEĬ$�#^�f.�ܻ)�CIYP;��ԫU��E��GZ�q</u�ۧ,U�َR��[zr�M��L��JI�䳪l���jM4�+Zi��n���{��V�f�eV�*�c4;:��fPc[@�t`v^f�E�`�~�&M��lSDLT�ݪ�A[C.��kb�N�,^@W�*�p�N4��M����)h۫�v·�i؉M�b�P���[OZ���:3��K�[h(�����<�U�P[5�4��
�.fր1�x��M��E�L�9Qf�拫֚�Ƈ$�z~6,+U4�S�wwj�ׄ����b�YƉ�&�mͩ[�Z5`U�M�}g ���C%�Yw�V��8�[�gH������īC���zvV��QɁ:�t(eՑN�mb'/\������޽ %O2�,*͡W�6cHL؜�aڻ��VS�1ͧ��4���Z�ɩ�VYt�1����^Srn����S��\ِ�YR�K�����9�xۃpP���X�ڷW��a�S�l&�oZ]�.����X�T(c�up�,�Ͷ$&��2.\[X.�:9�H��d}gr���҅��u���z&DF
v@������(����:�z�T�1k��떙�����{f��A*N�7I�{2ݍ�S݋^TD:r�
�ߦ�k[/1�n5���7��z6b1�$,�i�L�n�T&��G`�˴oK�[�T�a��e�����\��%61�S(n\ѵg�r�5���Ӛu}�o2�f⛚�M�yO6	)ݩ���q53y�kXm8�Wv�΂e��)�@^Ĭ�ݍs&�9�Z"�ˁ�-���+%Ѵ@��Mqt���*����8�hۢԈ毜*��LԔЖ7e(6v��#�y�#��œ`�,Tɬ*�u��R��ź�A�� �kn�	I�l_]L�AB@�9MD�� ۣ��;"y� :(b*I��f������mz�Xke������ŏN⠊��S�%h��pU�+v�Ztf��	�:���U�.��jYo2����GA�~�ʶY��m[p�CJn�k#(M׈f�P6��)n��L2�k.R2�OZ:�1��K�Nкrd���gc�n`ĩQ��x�.`��m�-6S�J��#rA� �j��!��aI��X�@�7����NE����#�աhMʒxn�'�s~XXR�m,ImQis��
҈:�(�%cEJ��F�ٖ�j�t'J�\z�hg�ͺo%��R�bbޗ"������V2��A���a�n��$cD]!�M�ݭT�'b�we)y���a�-�,� ڛ,�wP@�F*�k�u��ЦP��JnЈ��dj�LR`'DKX��$��������ǹ���-�Ҵ'yz#�N��ZU46��1:�v�l�.f��rۭ�l�#t�C�m8�ud3F9w�p�EM{�>{F�k��2�
csNSY��m:]��u�����6�23Eh�(4���r�-�r�4��`��Ս���T6/�?�V�y��AQKiVg0ۼ�GQѨ4s]Ě���U��l�!�F�[:J�1��,���� �V�f� %*��5���XF�s�4��9�j-�u�Gס����1��Z���2��9������z�#R����^3r��6HEV�V��k�@�Ȗآ��$}�[�D%� X�=��+%@�͐��.��w�m�������*�R�<+ʙ"GMn�W���h��J��G@�r
�G��$�r.�2��m��h��{1e��P�NFT5��KQ�)�5��k,
�(�;Me��V�\����X��b��K�;�Jyt��X�n�-V����H��@��7�6=�3L�oT,�[��LLir:��4�+rje�mX��P5���C.�l��CQ�Ӹ,.�"u!b��R�w[��h:�Ihv)�F��Чvp4�f`�W�Ք+m�X{�əi�B�m܀)�t䲔T�"���J�S�ܹ�f�5��A���F�̘�D�R�GL�y�#����&�1e,��1V̔���[̗r��zك2nBb+�F��,���s5���a�f�sr��C퇺h�fee��2+�N��5�V���:�I���k��#539b���v��JP�ї��
I�~��g#�w�h4�L��&� #i��_:���N�lM����Ae�e���ؠS�.Ԕ4(��β/�6��$�E���3W�Y��b:ք(Y����n�v��Z��Ռ����:���Yv��W���J� w�U�6br��(5, ���H�.�	��J� c�n���K_�j�5�]c�Iॣ4Z��e�8J&�m�tm��i�W�3X��p;�2��2�۔>��V��T�sU �U�ɫ��ec�A�f�@6X��S�ِ�{�e��ٕ�4:�n���Z�&�:S$V�&.���4He�z�ø��dy�b3l
�kTU1b�,�"��Z�Nxt�1r��u�E�ѓ�H��b�
ͻs4,V@��b�� ����"����)T���3tiXծY���L� -���� �wjԚ�Z�6��+d:�4�2u�E�e]���I۷b�ln��b���F�бC[^n��5Jt��6�h*���D� Cv�ݥ7A�i�ܬ+	6*����&uS.�1R�i,�,a����ј�����`1-� ɮn����ѧK,�T��Q[QX3f彷D0�7N`b\;dʘ�ǐ�]�8Q�GK�!�d8/�)���z6��������V���`���b�Ub�J��S��\��b{|�z��v&�rbR�B�b<���s���Uub˰�@qͦ�wH6^bz���Yx��@��V��)�M�+�N#se���`(���0���h�Ɓ�[���Ct�,�P8�PG�����]>��+H��w;�m���!ݲ�� �b�z���C2Z@XbT�v]JЬ�Z��]��ȑ�SY�P"bWd��+SImm�h+m�5{D6��Yr������T�P�.S�k^��J�95*�p[C4��EZE�.���e���Oi�9LJɌRH�A���1[�J�\�m��̗�� �+f�����3�kl�o+n�;x*�J�������,�x�D#n�9��3,����v ��j�����% )�U��ʊeM���"d�w� ��y�%6�T�S���Ua�40��
y]E�}֋�-;*M�ݨ��K\��b�X��Ǫ0�(�f��^2�5��k:nʱB�M��zM��f��W��1h�N$��Cj������U��4fV��ݒi����[�G��t�ֺ�`�X+s�Yv��.�k��������M�iFSՙ���ٮ�W���KѤKr����U��%v�1�E0�e[p<ض�4�ͩ'��������#��Zَ���T��2cy��)ati��2m^�e��j�UՎ���R���f>�5���`��r�ȇW{���M6�cMͥ��+ȳ6a��V9�f+�(<��B��t���mB�;*�l����XJ�55,p��Kp�dZ`:��/�`Q����V"6��	��iͱO[�lX״/�GM'�0�;I[A榆�W.kň��򑙤+N^ɦ��|J:ن����$Q#qKv5�f�ƌ�Ra�FK�)�R�YW���Y����]$�t������*���-�ޡX����-BS{�:���֭�̣��T*�7V�:@�^�Z4��V)��I{��ᔰ�������*���Vޟ���:�n	�ײ��r��3�ȝ���j�eo�Q��_ޝ+i�V��M���XIYk��i��6��tT�µ�5wXa3J�������^�V�P��MH;�=MbiN\y�o^Y�]Q�X�gD���n�>6懚��X��H6/s:�Om���(q���08�:Ή�l���3-�� 5bY��ݮ-�1+y*�K�Z.���A�[��f�8sK�V�X�ۗ�N5��y���)R6��d��t4�W���j��<�����{����qH��-��eл]��S��L�t7%	�'m%��ݏ�,̒���6vy���V�����5�'\����:��xit�ƪ��ӉNTy���Q��2�d�T (�n;;98��4�w͋{��̄�Om���hϖJ.������C��Tא�(�[YCkb�]3Wc4r*i�Jltq� z�=����e�Vl {T�u��n��%nE�ڗԁ��Uֳ1jZ$ё��u�%��B^F� UipS.Z
K4�Av����;U��+�5r����88n�u���f�&�h��wzt_#iF{�yeYbJ)({g �om`�"�q��I�)y��ɯ��9��"�ݡwݡP��S��1�6<3wẽ*��w��B�eD�0]�րtV��$�XtC��=6V4v������fN�]I�����4k�$�R���y0����PuY�J\�R�:#7��9vRɣ��][����)Q�)�z*D@�ܽ�;���<���`��E��CYڇ"�4��9&���%n�=�i��m���HzNF[�U֓���x��a�uً����ۈ����<��8���grY:����4׏LR������F�+��4��7%A��OX�Q� w!������z6�+�3����S�2dΛ�ͯ��	���\�MW͌<8��v>��(�`��;�vK�윅%��rD�*�V�F����4}��J����a��;�6m���v
�m���fX�#ν&gVٕc�E�sm��άۖ>O~͟7�0V�ԫ��hm��ԫ/v��n�N|};4�V-�y����Y��s}���vTl
���j�V����8��|5w�ɭ-��ɋ8L���E��\��B�=B͘�T�	�3U]'p�_������� ���%#6�XA������{49oyp���Z�t%�La����������W}��s��zړ���z�0%-;ݮSC��)[{�O�4�\��'��������N��̱"Z�}�/*:w�2,:�ڛp��7+3D�{,GǓ9.�(�E>���ɟM�{���'M��e;"�V(W�r��ntk�MwW�ӟJ�{yi�lǕ�C^��%����������vS�rw!T�9,�֮���V�(x��F��)��̣
�0�Fܤ!�^�`[�*�-�L�tr����`��PF�̙Z��&;�ux�\��*f�fKD��`��ڼlq�N뀕�u�7�qi+m;45;8�(�9��E�n[H\`�A_oDEI:4����IGE7�v��ݗ��9�[Wb�U޾��k�_������^�Eٿ+�n�w�����2��B�X����+�ޔ�'k36Lٚj���-E���Qڱ��co8q�GQ/s��Э�V���=:󓧒��K�q�X�Q=�յs]��{ټ�8Vv8ck{-��,�uǡ��Yyְd>�J�Geћ��8��� �V��r�fm�,7��0��)�$��)�V��׹kb���N��Q�wo(TF�8P-�q���Vs��2��t�L05k�z��\fTX�!���G!���;N#�ƅ��X��k-̙Ї��oJ�JF�3�����U
<�K�g��ߎ��ip�*q�D����\0ƈ���fe�E�We�טsWs�9��=�D6zo<���-cDA�e��;g�łfou�n�&�th��f�c�T�Y�H�͓H�[N<%���x��B�&F=Ω_�b��ҵG��C�Axb�۶ %��&��p�VG��V{}�w��6OU�޻�
쬠��5�X+��7ۆ���G�4�퍜y�]᏶i���IwC������n�En<��o�[%�U	%��y�ӫںQ5�;�*\����;4�	\�]78<�[N�Wv�m�+�1d��3�{|�Z׸7x��y��4a�r��f<��PJS519c���� �:�s4d��P�&�3�<�G/��ƗM��š�;  t��W^��J��F���A���z����o� �]�b��պc7���B�_v�hNt2��QN��uh���Yig
�!���"�p����\�X�R�`ᨷ�k��B�-۫Lr�Ӿ
[�ec��f��)z�a�n�ǯm[����j)�2������$h����r���NC�\'[����R՝{zK�u�v��k�$a��5�q���e^>����w-�֧y�flm-��.Y���ڵ�yWZ^V=:z�+����������N�uؑ��Njp��E�r�<�/E��=�� v�ef`��j�e^ۯp���D����.�D�m
�s(�kt��uk ��k۵.�Sd{S,δVf����퍖�{l9@��N;ޗ��3aX�
�LJ��GAQ��B�9�:�
{t,�C^J��Ŵ����b����#ok4�f.P�4��.��ҝ���:\���9�5���U��C	e�e�[����+��n��P��wX�cŰ9n���kr�ox�����Qar���Ӹ�����9w!��e]<T�U"hN\��y"	r�'ƻ�Nȶ�T��[+h9�,|nt�E��Q�O�2��Z����$ U��%�f��\pP�KM
��Tb��̂��ٽ�<Y�F1��zd��2�%Wm1ɥ��N���)�@XO^��Ϝu6լ�\�[�
��cF=� ���6^nj�Q��$wJ���-�Lp�S�)�c����h�U�*�X���6$�c-��	�u������Ǽi٧�W��i������v�Mҹ>����f2�b<�<��Ȟ��Ҭ�)L�m_2H�w�.�7o�Z���*�8T�XGf�*��택>d�|��f	�����-��ڹ�9�DVv�F�H�l�|k��D���2���]�Fg]sz��p+ڗ�Ji5�^N��y���|�3�֩�o������;L�Z�<��
fL*�Ҹ�T�ɭ�J�����T�|�8�4pm��΄Y��
�@�"��J��� �[O-l���%�R@����p1�2�Z���H<K"PK����H��y��*2\�6�ܒ��[����bi��7�:��]�+{�8@2�8 �j�nAǩж�\I�(���k�ҩ�+��c�����c-�$T��u��pձpq�|t-�\l��݂Rh��� �\^`CEm)n����8n�����4�L�]���*�T/8a�*��M�� .WKEE{�������
�q���D�b�r��uY��,[h��32�ذ.[T{����;�%>���>�ٕ�^,�i�܉ԝ�5��u,S(Yz��V��t��� M��Q�鄆�Si��fI�`�i��t�1Nv\t��ƱN�vz-���WM4(l<��il�:�ٮ�勥jfQ�fWX����Z�95�3D�b���V�"wQZ����O^���-�6�	<Fna+#��mjx5+�b���C�!�0������X�q�k��u�؂H,:U�C�ũ�'vF��)B`�9�H�Z�SF�艻\������Ǣ�7B�sw�]Ơ��6<�pW��6��%՘��rp��;�"s�/�<�.��յ���G]d�J��n���5;#O�g.9>�:��Y�S���jqk@���n��v�̝]l�Q�2�] �M�� f�f
�9��x�x'u�C�Ry��fu��s�=w�W]u���]��0�8	lm5a@j�t�[�3[�X��r���N�Y$�u�./�����+VY���18��zr����x9]C���b�����E�K8v�S�\tJ�;u=��f�ev5Άvvl����PSb�ڙ�M���,�n��taB�n�	�j{��ՓJX��g��%���]C�^ɏr� y�l(-5�DMf�t֮[i3 �4̮̻{���5(TyN#�+�U�ݧ;�S�ٔ�����4b�vB��p͘E�O�I���!M�n�*1u+[�ڗ�`�y�$�̭$�݇�.����.�wG',�J,�)��;p�K:�x�k(����f��-��7�c$]��s0��ܜV@�f�	W�a��_jܭ&��Hw50T.���C&5zifk�@���G,0zٝ���RHےI$�I$�I$�I$�;�3'by	uN�έݜ���r�����M%R�PLU���G�}�c�Cycfx�:h��53)t�d�Z�O�o!=�|P�ͽL,�3��GN�,�w*Y�,�W�/��
�u`�JO�o���<u�T����'��I!$�?_�&�8�_/^	  !�ﬄ	�������@���H ���x<w���=}ν��f��t��qV.�3��ŹȬ���RH^e���o@��뵢�g%��/���bqy��L�����}�o������Wkimg7��a����0S��<���#����������/<�,5��S�� 0��F�9r<7�h��H�8���j�8�����}���2��|�������n�0�j�'_!A�����t���a�u��R�zұ,.ycJ���+��FU���
�*+�B腷�e*4Hq�
H��q�_=0�Ѭy�V�H��w}].�]6!��U���l4y�t���]>қ�������Z����ȱ�.0w!�:��[[��g!�m�\�v�-�u�\z�V�C*�o�u0����0nq�#�W�ORM�Yo7�#h��.��
���[:+zGр2���[ɏE-؜��)��pͱh�=�����q Z�W�=�!ө8�l���of��[�:��
��4��u�æas��E��6�vV� �֍�WGln�. Gh�+;X����i^����|���ll�,�T�`S�{�k*�3zs�]��[$J�"ټ����H="�S�cR�f���pu�u	��S[]i��4D7.���B2m���q>�����/��[���E��l[��j�cl�VG�qmb<����M6�8��׷Ě�b���+-6�7�e;)����ht������E��������'k 8�鋩��ف����f�ie�"u�KU�e�ýJ�f�O�,:�H  ˽׹MQ����{�9�_^�G�aTb�}ɤ�A�D�
�N����������;D����9��z��K���:U��`+�B�����;�=lU���o���Q�W�
7WH����D��ky��j��p�bk��óbYb�b2ݚn���pʼ�3�R�<cnk�R��R�1�� ���ib2},� R/��c�we����I�QZ�*Y�Ç�n�GU�M���/j��h:����OM�\�3tP����;W"2�HT2��0�4z�#�
�����c�n-��}
���2bSw�tw�=͕��� ��Ap�N30�X�r�;�ź<��F�U�l��t����#ݚu���_1:Mm2��"`Bu
}���ˮ7�NX!Q��&N4(cg��l�S�(O.�4y�o]��6����ub:*�ӳ����gu�F��ζ��ޮE�l���1�ُK\	��w�B�t�G`%�`���T�+[*��t�����b1�w/s������h�֔/5r����7(+֍��׎Q�l��/�c+��!C���nTWۊ7���y)��ے�$C��	D�nNIŶic�A��|�:Dn*�} �,���	o����u]"�b\�R�Hˬ��W�۵�§!�un�Ӻ[Ơ[����}γswi�pK�l��%�Q�g:-��ʭƟEN�]ƞ���V�m���J���cZo�I���3oB��V���T�7�\}i5S�˩6�H�m����L��4umFs_AN����t-6��g���J�Tm����H�)���9�X�LI[�����p\�>���;d�	4�󦼳)Z�t:���-#	`\���[��H�ʷa���p�Ӕ��1;zt��Q��-��p�Q�7}�⃟|Tt&L��tEzޞ
W>�Ont8�#������Ҷ����n�P����c���71Y�&��NVᵪ݊�{�]�Mǋ���^[�hgFt?r;���N��!�󸊁m�FsǪ��Qt�I9�f���م�����[�
��]��\�*�-ѫ� 8)SwYƳ9��U� 7o5�``�I���`Q%��P��Of���ʮx/��W���6�Yuxec�#�t(&Q�ُGu^�{B6h'�'e)��#|Ӽ%+�� �� M��{t�u���V�eԹN
;�ڷ++ �[,��ٰ���w"�W'w�`�o����JE^G�(�Ĉ6��'W����Ğ�:��Y�+��O&U�y���XO�$�8��䘃t.���rk�Fp�R��b���6r�����3pԾ�{-�&��Sc���GQ�V������av��:H�חًvY�Ŝ���@G��,���^�zb�u��NX�S�7Y
�2�v�"��K��Y�˱ݻ.c�rI��:b��t�N9pV�%�ϳ,Iԍr�W%��u��D���S�H�%����n�q�c��ip��� ��b��70�}�.SMr��va�[c�W��I��*;�&ޗ[R����p�3�VKv�^m�Ya���w-��O.u�Z���G��f����+5�P�h졆�p]7f3�\��u�[m+W�~[|	���-�	�ݼ�yZ&��V�,l]n�}"��]q^@rmզnR�{����Z�WFhhͼ�U�g��	�F@��2̓va�!',�3vn]�f9I�r��_3Ǫ��ت�a+v;� {�sC����@OV�\wz��2UCɳ_C	���
7N�z�ur�<�]
g���v,5�]1���B�bRZ���%J�����3:��B�L;aa�2N�<�:�;`m��gHKn��5�FXk���`�h6�|�.�*+e�M/��nL/�B�ħ_m%�ihF����(݆]fժ���ڵ���u���5�=N�s�k�q�Z4J�e�;}xh�=�r�tB�M�K�g�V���uj$�W+Ό��I	t!��!o�7���"T�f�ů�s�Q˦fgd!v��[۬�	�\ӕ<T\λ��]u�;�wb��u�fc�/�dǬ��5	�O�
��-��,�W��v록]\����h��[t-��hK:f��g��֞��OU���Qj���!��XwN�Ӗ1��n�f�mV49�{27�Ս�3��+.dٺ�	lʱbN2j��wŤ챇�6r����nRണ�<yWY���8�Î�i�PV"WW��η������6�oh"�&��D�*�p�[7U�N*�Z�h6~�aѳb-�2�}�;ګ�79��躜8-֎�ҳ)1NX���>�fk����r��!܊#����e9����ܲ�^puX��sՠ�.S��r��9ӝl!׷lom<AG%��]6Z+RYLe���1�F�T�����Pɳ����k�@Pe$�F�߻�`6�av�����C�'� ��\��՗�NV"^�V����޳yq�g8l`\�o�_9ã�W]�멊�<ٵǯ+S�0��$Y�1�ݚ�������N&x��8��VR�s�����z�h`�����<�|rV�-��zrl-�!�A\�N��:��j��-�Ǖ%���wږ[[�R�Jg6��n��������nt��T�8�f��Z\"C!u�ٹ�F��2�]�J�v=蚺+1b�f�����&u����mP���Vj�h�Bp�)˷�$�k{�<W��:�tA�nvR���@%��J��o����u8vGgFh���^<+V�����ۑ�DP#i�i�)������ �������Ok�٧4���Gt�/�X7&��swi$�`YM�̠��j���B9�����(t�jq�B�PCw;��ש�7ۘ�m�֤��*����X�G�Gqps���BJ����9�����9��Xݬ��԰�J��%�wV[9�Xqg\Ł�N�0p�.vb��L�����I��&�&��7���&w��-���Am0�y��c5�/n���t'�Gh��6ؾ���A0DNʳ�Y+:رXt��-����.����S}���'y]C�;B��]"��:j�j�Qc64'�;y�4ŏ����=Au�ˬ�.�"y� �W6�eI��5}�Q5
7C`��B]�<��!��#!�,㮂����1p�������[�ض��Rǉb�p��yD;��9�]�lҲ!L�T�}́1Bwg�5[���0[廋s�k��I��hB2F���_Rye-���SJ�st���B���owb;IR��]����f�������� �hY9[�\�N-�x�0͆E��T�*7���Ջe�͹xG],W��P��%��f��K�A��B�}�L!�>g��E����u۵�uw)�4�ͳgjn����Uƫ��]e�vc��B���
wt��;q�,���*���;��OD�Ui�yM�ec��������gZwk��sV>ZuoC!<*�̩�.�;�ݾ���	��4�G;wu��q��n[zpʽ�N2F��'�*J����3^r��Ù���:'���]a{,m���]u�*�P�v�(�߯��2!�����aRUs�����V�c�h���*�\�l�L�6��V-��f�{�eym$ ]���ˬ<2��&�)�����e]�b
�GK��YW/���u��:_u���XV�vSJ�>��Y�>�/����j�����_L-Rv�N����
r�-���NW����_��@A����9!d|m�qI�>�?{4_�Wߪ�Y�&t(�4z�T`��#���v�f���k����+ג�-�*>ʚ���)|��(�N��s�U�be4�C0����&�+%q5twj��4cw݅�l�����v��{��{���ǎ5���)�����t��MQ�7��#2���휻Q���Ɯ��.ݑ��![o�IX��W�����ƕt�2#��;|.s��mVo�=�jn*Nj�%���i�������#�3Yp#�/.�qI��)\��Y��>�|o��_�-��Í�u�N�ofQL��@�V���Btow�}���i�d�:���O��7v����v�6.�Q9��t����Pͫǹt�e�գ��3]X��]J�:!�]*ؙB��r�f�CzibV��-L�綄�S��ˊ�oٴ�����+y ��������W݅ő����
��-e�cͩݨ�j�(�UH����QeX���"��F"��PD�6.3,YLeD`ŭ"
��VD��U٬Y�V)X"(�b�
�EP�D��
��-��%��V�mcR�Q�U�aZ1�!�QĶ��j�b4f��U-*-v��AT�+c6�l����ٮ#CI�ت��BԭSW2��V�u�TE�\�I��֋mm��(�2b,h�ªU���.��\LDUuj�r�ծָ�EUEaZ��hl�e+J�TZ4a���"���X��H���㇞��f���Y�l�kd����o�����u�Z �5��'h�}]��3���A�}T��ɽ��W��N�d��
��
�T*
��LA`��*w��6������ت'椀>�hwy��xi��
��_txիM�W��qrbp�64D���kA_EW�&�/��Y�w�癇Q�i��z��~4`��*�Z�� �]�p�C���c\�e��k�j.������D#��S�
u8*Zj=��K�}'{۹Pz�A�ˇ¹�Z��i�\�QP�,4e��nov�+-�i�=u�P��=�6+��
���:���u�H�۱Q�r{x�޷���(~���Ώb_[5~.��RwΦ��4�!N�r,.s�.���B0p�zfc�J2b�c8��%49��B�C�hѐ�UC\�V�}l�a!��0	�S�g�E+/�B[�:
�[l�_1G��%����q�y�$添V-�	/vճ�=�9i9R@��]��4��RY�kUv��k�[x^E��u�*�ca/w^ig��irR[�Nw��w�[8b9��1�.�&@�4����.�Ls�;1��Y������c�^si�ҙ�G�r��{ۣ�Ƨ���i!H���ׇ;U��h�lxX�0h��(2�Ou�&�v�]��*�J� �'t���C��'�E��?��w�vp6�4D�c�eI����M��
N�]vH�|��]Η���8�HȆ����p���'E*�c�,;,ڙ=9ͧ�PO�b���͕F��!���ݘ4
�N�&��)��63�w�2��b(A�:6��1�)�n~C�aL9��*>f�1oo�c�x��C��U�>b�a�m��J�5Ui�k����z���(�[�Gؚ�x��x� ���m޽�+<aו��m؆��O�U'J�(�*v3��)���5���&�J��d�71�h���	�FjN��m���ZjK��3���OV�9 ��Y��6P�F�*�ێ¤؈�l ��Cgk�{����!��Flt��uf�"po�ÖzyV��Lv@n�jS��K�u
0Ei�~1�6
c�.��;��i����v
cC't��=����8A��]9�*tkD�o5j�[X����	&@T�1Vc���h���8GG�`B}mrP�&/�@��?p�g�Y����l�E�|2�
��h��v�Y��86g��t�]�H*�^�R���,����������W�ʠ�`���PT�D�,D��;ż�W���I-��d�u"�1'��!���#�Lj�)�n<���{2��\&� }x��F�u���OiG��W�h�Y�)����/�a���H3���&V�觴���N
�����n-/\�*2��㵆��=,��֫+/A,^�|�ֻ����v��V�H��yt�E�������k��n�YYK�׵ttU;��72�M��+@�ʶ�,\�B�㧄�J�]GT���
���aR+���@s�7f�l�mR�ej��B A�� HAQ��1�b�1��CdB�ox7���Y¾uQ4�<�ˌh8!!I��~(x�}vdڼ����oC�䣮� �
�9pxx�_iY�.܇N�U^��H�+K�7�	�b4hC�q���a �PZ@�{�'�=(ea�\U���d: �<)i���Gm�Q�)l��5�+X&,D��RU�XCBi_��ą7W����^�ֳуW�{f��}�pp��Frh�����L�t�[�}�;
��=�.���>�>���T��}n �*�<��	��2��5��({e�3ݱy���ի�ͺx��}K+z��R��}�[�X�W���x��7]/y�[���-ve�'��6��[���9%������#ͦ�Jn��5A�;z9�՞�2����\pR�YZr*�	�֭ �V���m�\c�8��э؋�1WF�xK��6����>jsky�l�n�d�1P���c$��a��S������)D�\`�%=+M+X�n~! v�<D<�"b�G
��[�K�,%w�72���FtX��;���4(w&�eاt|%��Ƶdn!�6���;��V �S�o����[���x�a�4\�i�g&�.t@��UC ���� 5�b�!V�}�gbꂢ��Ǚ�X�ٞ����f%9b��u1� B�Oi��V*��r/����0=<>��@��vc���и�T3���1]?u97��6�E � ц$P�4���Z��Fx�U˗�x}��iY^x���`���{�;j���q�]eAbM��f�ym-h��8�V��R�7؃y����Eb�%es�39ĕ����i���Ƨ�u�b�����5�ͅ�5��ӟ�f�u�����*#4�_nM��Y/ijK8G#B?�	����!�ݍ�����EI�G{.3�5Wܛ�� ���P��ؠo�xh:�2���\�f����з��yefUp"���\4�֍�4���
���I@��S�3==�p�}iV�/��4gÃNqp��kE;���P�s8���z{����R5 
��_�`��E�҅��+��c�np��i���c�¨�I�k����lun�)���z�T�l�uj{)i�t �Rr��c�u[�փwᶾ@���ku6���+�vb�Cr�V:�� �)�&�JT0��=6:�B�FYO/39��*���hpJD��R�1��Lv�xD�y�.a�0��5�̫����o�k5D�<L�����*�q�[�Y�1`�&n�'����gp�����:��r7@3�ި�:�
mu͙���L�ǥ�ز�N���G޶�.M�Q���s;Xo��&0E��-W�t�6n�n�j�w8�1R�"����cS��}�� ��Z3[���@�ש�����j�S���i�Sk9ZUT�w<T!���1�$>:0��3���jb�	�g�Y�'E����R�p#@��d��U��5��z*��r

���^��11t�>������j0wf2I(P�'S8���JV���}8���z�1�-5k�|41N�MVP�>7kc�>]�R[��Ō�q�;	���N��]e�NeP�6G�]yr]�ss(ѿ�Ԕ��LT���u
�x�9�����ne�t�V�`x
�c�a���f����4�<�jFjv���@�cl����[����"���+�ݗ��+���rk��]
k�&*ё��(̮-�ޡ��i�V�6�]7S�r�Sջ5e^��N�#�Bq�*�ڴ:��'.u�Ӳ�A��6����C[e�W��-�v��*�pz��I�͝��$j��d�s2�ަf;�w��|k7�A
�#PJ
�L���#o�*Y���X�N2X���eL!!���)*�&.�ş7\�H��cn�]��2P�c�IK�8�R&�Din�� �mr�����U�@��� �ʎe���#��<n	Z���i�\��>���0�	�x�"x�P�c���~l���lÄm�>jP
���,h�.^{M<ٔX��8�>���ߟG�WrGK\ܕF5R���j� �f��^�EgB E^�^�"�i.�۝u�G���>g-�Hh�3J��� �����H����.媂�X���T4-_�wb�|�}3����T}���Kjk�����x���myoV#ܗ�gs���k�K�8?�=Bfb�;�� N���PV��RYZ�g�.P�e�r4����&���T����F���s��یt�W�6gwfysm�t��{1ZMw�!��~9���U<?s��dT�s+!7��?Hq�͡�����)�; V�m�:D������7+�A�;��*h�O��=b�<�:5F��n_�N���%�z��_��J�pcF
��OK�
�@O%G��/��[�Up��:1��s��w���H�r�r$p;!Fܿ��۬l.s��C�^��S��?h�(1IJ�<�}u1�%f9kcs	��@�w��(!_�lp[p@�����nm:�j4?�ѡ�@b~�0bw*Bp��W?V,���sHVo�Z�ր"��/����?An�i!�q�5o����z#T�g�!����ը�͂���E���+�bO���W�6:TgzU�4���l��u
��of�\]�N�19eN[Z�ugQWv(򬴐����z��R�ĸ� �˛���*0?��z�E� s$D F օ7ZY�y��;V��G�+!>ã�W�`3	�1����=��j��\��pAHz�c�W���뼽P��!��JK�\Z�ʘ�'}�;��`cE��������'������	vN�ֹ���Xp$]a����+s��� �<uYo]{����HÁ��E{���D��U���x*ʯ�(ųa������'�W��B�f��U��K��X,X4`;��+�P���WC��u�s݈h�gA��5�KUz~v�
,W��{վ��m%\����\�*�_h���b95�J���^C�ݞrwM]�X�D0C:�}gDK(Fi�t�C�D|��������8�G���h��S�tu������MHr�u�oACU�W�i�+�;ATʺ:���\�-��1N��f�r�.�gͻvk���p�N�t� j����	�N9w��u�	Chq�R�r�Ɔ�b͐�x;�j���_:�$z��a��t�gG��n�LT*��||0�b�2؈
T��֗��'�t�HR�lP���n��5��-�೮�[W�5��֊��CB�]
�֐��f�t��zU�n��ϓ�rTRYCg1Տ�8�ep�Hf��G��lv=��v��)��Ko��f�n�mɯ7K%�x�p��{�f�\4џKg+>[@�Z�J��]\��x�WU�6�\U���f7Id�)�؎�19������W<];�Mz(�u�q�Skc7oo+1:���=��h;�9��Ґ�K�l
{A�,?	w�m�1Լo:u�C9Gfr{�:9�3�5*upX�:�uj���oV:��ܦT&�7Y@��8�m�I���bmGGGG�����ж��{v.P�@� ��;.ʫ�3��˝T)Q�ٚ�oQ�Yc$_p�e����]]��v�����eۈV�֫��C���);b �T����.�[�nf�'h����v:��+��]G��zV�b�Ծ���B�ʂ��}A\�U����a�;7����|a�oS笜{�.;���p�j��7���8}.�qJ����6CFa�f������6f<��u��m�+َ9��1�:��vhk<ؓj;w�L;�t������4)2:_�	��c�תk�&���Y{��}S(�%f�T�Y�M�:=����t!�㽜�C�����Q�0o_JyO��lӘ�U�0��qi]N�-�L���Qes�{c�Z�X�Ԩ��
�����@���m�f6;$ǎ�L�}�[����V>D����T�É#
�m&p�f����=�p��֌έy���ŷO�u4D܂�n
lj:n������*i㍭�˾��	�����g��K��mj4�hcb#Q�`��z�LM%[B�Zԭ����(�2�,̸�*�cmJ�Em*�`ڭB�jJ��
�U12�J�Di�Ӥ5H�b�Tb1b�ƫ���0T,X(��k�1�X���R�D-��T-��TbZ�USV�eE�d�
�,ē�QQdD*��(�+[��\@�Qڣb�Z��Q+
�kJ���Id,AdU����)+EQXVJ+E�J+#
�U�l+&Z���"E�7��]���xۮs��5���돎�5Ս�q���=]�s��s������ ���yβM�����"Nޙ�7����9M�M i*Au2�3�6H(lx��C�
�����A�Ô7t�P:J�s�	6g�"#���ܶ���yz>"#�|@����NЬݒ�偤��u�z�n;�v�[`*���'I�c�Ձ���������Vr�,��H*��W0�9�5��wֻ�Ht�uCR'�6B�<$��� ��J��h��+���ެd�
��W��̋&$k,��*�>������`����]���B@r��
�v�<��i �&�Rt�`o�f��xLa�+�'i�����<w�� �k�1YRT����^���j�
��DPZX�=өΖ�~��׈p��Y)�V�&�c��"�R�<�զ��0ۚkœfbAv<f@D�>��J�`T���
�����阆$�^��~�N�o��x�~6��]g`b��
�����AxCt�H(�������S�@P�%T0��r�{d�3W�x��|;$w�ɌRa�xV��s{3{�����u�=��Z���E1t�h��Y�* �N�y��M����zAH(g:M$�
���X���x�| T��E������#蜏g�ɩ}�+{;ֶ��T�̞&��4�R�膕��\Y��B�m:��-@��:IۏX�U��&�l�I��=���0�6������:���^7������LH(u����+�6i ���bA@�T��t�Xtqa�P*�dޘ��+��{�߻�t�Ι�5ݓfc�f���	��k���|�u`"Mݙ�l
���x��JɩlY�xC� �������Aq���Ad���CVl�w�*$���dĜ1|��>}�3�Dt�`���uoV�p�>�n�Q�錜y���ߘ���j�̙�E�I�k�F�ܘ���恰�󆌰�]�6<�X�W��\g`Ǧ�`}�)��Fo��J��4<ğG�6�KnO���P#��uU��*��n��4�LY��&$�h��d��N.�;J��Wb�6C�bx�Ă��*M��]�T��	�����.ۺ��w���N9I^S�R�f�����
�~�M�&��N(�7N�C�!�C�p�t�(}��#�^�f��̌��y<��� ����LI�ZE铄���@�+%f���bAN7�b��5��E�kȏTp��xpw#|�gubMs=c}�
B���h��O����Q �g<]��-Lv�B䉼7|�V>�B�ń4^j|tդ��?Hh:�᭷�ʳl�E�����`��0���#��&Tڊ�U ���%Q�"�j��z�V�5ځS�P�W�%i�.��ܗ#S����=�.oʍsf�Q�]�1�N�\�����,�����տ�쭙��7 z&�����������T~�~�5��s*�(76�-H1!0'&��J�.��^$><)U�=aSAq��u�О��d$p��E�!��6��ۓ�OyA[mbU�M�R�U�z�+A~��=P����/P��WZd��nI�5ي�-���ݩ���Y��_ BX�(!�:�k�u����s�YX���K���={T1�z��K-�5L|Ю����2�?X���⏷c��s!>��U�x4�?R��`�~сs���N޵�q�6~s(U��@(Sw&��pP�`�_e�}�]i4,0!	����1|@���4��
ZX�c�����M�${狅?XU!뤫|_�
�W�x~��_��8�9���7#�}S���gn�k��@���{�x��H�:si��.F(V������]�͏0����mlo��_z��%�s�V�dT����^�>g��»<�s�ҝ�\q�鸧V,�]N�+���Z�/�s0.���; �='Voť\\�d�Oo����ꙃ
w߫ˇ���
���%y��D�s&z��4U�@���_,	�*��!����y�*���5�>��"�["=�͒�ȣ� �����n��չ�q��v{OV�">iC�v���t�7���2���uq��뼻��M��ku�!p6�6�:�+�4P��='�𺃡3Խr�w+�՝L��r�濤�+o?l��a������R���P��f�];i[�����N�5U6�v庎*%B0�T�}�q���z�t|}������m:���ί
<����i��q��Q8�&k9	�u��F�"vFߦ�z����&�q�����!���Gy#��Թ�^	R�/qD�%ة&�%PH��`�u�a�[(��pO�CP9h��}L؝,�v��ߡH�@�V�r���X2���:�0�vVŻ�����}���a�
�m���
sMeA�[ʣq�M��&�����&2e��~Ȥ�n�r�	ͪ�}K�5�9G������!�yOa{^���Zc[U���o8Wo ��Ū����ܖ�f�j�&1VeN�z�t���Nz�wFm�F9|�_ms2F\]�g4�U_���n����7��~yV��~��b$c~����v9�u�b)(�Hr��Pu7�b��-f�y{X})���C�fC|�V�TUi@SԹ7����iS�u�7U9��ۑwn��o;!��H�ʍfP��~��AKp����N}~�U�ӿI9�"o�A�b��PVy��s[��s���QB9�"ˑ�Zod��wN�T�z�:�"����X�$ p�3"��Q�ر*,��N���b�;ب�ÍZ���Ր�i���|�vF�t��:��W�j�9[9���^�~^�7u$�s���G0�z���I���4׫�#ղ��g��ܑs-�6�;zo�S�6���ż��R�r���Ol���y���9nxb���yZ�iG{:T�9Z�tf�#�Z��ѻ*�^���/�3-_v��M�M��3Ur���l=3�G_&�bN6��L�B���X:ey�2�s�+������E5�!�a��hS�ʎ�A���Ui}Vmg�eo���Y��pIGttu�$%�7/��ޭ�)�Sy�����{MG؎���r	�R�[�WqBgha-R 3w��f%C���{[�O{G{��sZ�T��5~����c����JW^�� Y�1-쭡lj���k/��<��=���6?��_}�bm��������htժ�+Jx�U�fW!62�l��P�1��A�E���
]�Dr�PuqՇ_���Oi/W��>?z{(c�)qҪd��_Z=˧���|=��M�a�D]ɘ���Y�$�~�놚�0"��{�yOJL# ��7-���iiy��_�Maa�+�U��>�Jn�Vj���oTdt%�bi�ԥ�Y�~�7�����;�S�єT
\��~==��[�l����s_����,诵"�o8ؖ�GNm�l��v~j�h�ѽ��S7��0����m���0����'�r���7w�=�I�ꏓ�wb�;�#L��x�m���]Se��O�7�2�BhΈ���m�Đ�b"��XݺiV�������}��U��Ӟ7�R{'����ڻu�{�+\x�<�kwUN!q���v�۩�W;��=��k[e���R��&(��{{u�UO�-���$��c�}W��c~re�#ʲ��\k�5D�a�Gp��GOs�W�[���Mj��5�[���Zhe�����T,�Xt�Q0�2�8經뙽T˷���-��RH�+��Q�v��a���Nոvv�Gjߊ���܄�WJ����E�����k<�Y�ΜkDt(��p�����W�#��"��3|�W�4��^��������Wpմ��l]�F��� r�,����WI��L5�+l��+�Fv���~�"ĭ�Q�~�zs����1��KsU��e_�9c8�����ꯒi>m��H]=Fj���j���\(Zg9��H�ϴ5�=7�L���ރ��5��7��7؁u�޾�t3U1��~΋s�*{6F�J�,��N�����h}xk��9�@է�ոעV�ԋo1����}]}.�+�����ck���W�J�ٚ!����3���$�����OS����:���ӂ�T��u��EL7�5�����9��w���޵�$:��ا���یTt%����M�����n[Utٶ��]�?GU�������ޓ/�2��S��ں7����uߌk�x������R2 �ˍ�}ZFժ��/w�S� ��T)��ǒ]�4�m��wi������vv�����Y/�ho5O��}U_P��9=5�+����h�n8�Hrj�ˋ�6��p��`>�H���9	����r�+��k[}�vNA�1�\C��R�s� �mޤ�FB���/d�c��\Eb
O�ֻm=�F%��W�*�yƮq�q��X=��3�;�"�����
T2��R������zjJ���vC|��~��vz�*b�].f���աMX��^��=���9:�K!R�6>F�;���:/I��c^�t��n�1��Ǆ�,>�D���Li�f׋�����כ'�O�O���K�7Bd~ǧb��}�+ETf�vjYd(�
cz�q*��YG�������\k��u���%���$5�'�kݱE���ⶍ|��9zu�@�D��z�/h���+�c7���c_'����c�,h89f���n^!-�m!��/���Q�/�3��S����Ğy�R��e�ҭ�{�zn��-t=�Ƀ'ܾ}s"�-B�ReY��sFv�$�MmS�@f���;��86���`8C��:I��Omp��F���y9�+'���_g|\Pֆ,�v��i��Ṽq�c�)���Xil�S�5�kuD�Ƹ���
��_p ܵ���cQk�!��:i���@�L��,&5���J��KvJm�QX)Y�E<�8 9�[Vor�W�0W4��U�>M�I3oVS ��}����Z��d�ζ�;w����%v��w�x֢k�$��T��X@���.�Z:�����{B��%���w�]Po�3N}K ��~kt����J�B��wzb����Ћ��6d{�����۴��%H��̎��E��%Yc3����+L]A-ü����A�a�õ��PBby5�?c�\x�"��-���#��V�޾�%׳+��/�$���<ን+I��ۼ�D:���sfhuA�u��n���FFQleIQ�-��일�z�ZPc�0�d��l�-���mҠ��y����(<B����\��CW�,\j�{�w����e�=�T�)�V�L-���ء���ϱ�j��SAX�ǵu��J�%n���O0h�,jNc+d7�ΰC71��8`e�t�՝���w�\i���®��y�f�׽�i�I�Wړ���,��
EH��O:��Ib}OsN��5yl����E��*_r�nӫ��S�][��ga��K,�H*�O���(��&r.��� #.�����[���!  �VE�"1`�-Eb�(��b&����P��*�
*�`�"
�`�2�,E��r�#Qb���X�*�H(��`"娖�ՠ��"�AaR1Qb��DHc*�"�Q�$D"��X�őUIS1����YH�ªE,"�E@�
�Db �*Ŋ����X�("ȤX�Ta��"*��PPP�DV
E���lAV
)DEX�,����Y4���&{��p�E�-�)᝷ZK��	��|��e�[��Ŝ�d|�w�3'�UUW��(�<y���=9A�:�U�8){S7ߝ~O?L���6w&�Y�r{��-�ֶ�:~GE@�c���������j^^�����Ftپ�@w��~]�\I��筩�U��Y5�1��ȇ]tV�G���ź���=}�_�k���[�G��Յ�I�\�x���/�(]ť��V(ÃT�1K�g v������{��K���y#�{s�z9����̧8��nWY�|:-���+��ɩ���s��ֈq��Q�J(�{�z�u����o\m<v�f�K���F���L��{��o�ֳ�:��ݤ1�R�ܽKJ�e��[ժ��(K�s��o>ˮ�77KOL6��G3lL��y[f�pV�@�ЭW;���G�}_}_}T��m���/?/��J���;�R5$87�7'-�h�s�T��I�·�ʍQ�����i�h�=Ld���J���������,Yޞ�12���(�=�ܣ����b�g��^����zN�H'?c~���W3A�!�=�x]m�u<�����K�M����+C٪dA�t�v��2\�_��5���K���K��}��`~O}ȣޞ~�9R���	��������d��M��|�{ʘ����f��yjE3x��68,�k�Шc�'��]/a�SKP�h�[S���<��ʊ���;�Z�Ȏt�kƚ��{��N�{�m��l�Xj �I��)z���[�����
��c��t yn�/�]�M]��0U�)��UU_U|VV������Jw��]n,�8#�Ico�ع�tu�z���l��@-�|kfY^�o�I����'�m�JS�G �q��K��=�n���~3\��D�I��f@����|�G8z2byS����,d����G.�X��9����yڋoereI���
t�̍�oSZ�+�Y��t5�!��+�=^4�`���O�ɞ^��0����oJ��>}�qy�8n��5ɿL��o��5?]��\֣�f8�8�jN��M��y[���!{�_mײ)6[�b��~V���q���j�P�8�â�2 �N�]2�1������tw�3�Yqa�D�8������AueU sEu�Ј\�
b������_W�}��j�7�����b����U��Xow�m^��;���v�|޹���,dc��vT^�����^�k2-�J�j���\�7ܟj=�;�f���:|����r��s����*e	��]O��(�T�J/g?k���f{��/Y�9�rCYMv��J�.��̅<�
dkj�.z3��Q������;��N��#3ܘ�;�НC��Y�O,�novkpb;�<������QZ��FЃ��X����Ox�S�QS���J���\�Wi��=�n{�1�G�W�Hz\j��<��|=w�����h��ee�8��	���U��7m�0���j���}�)ݣۋ�֝#�� ^꽮
�-~��
 �s��Xq-�v�A�sr<s[;����U_}_%�s�)׮�����iS�s=Dj�*�n+_�Mnt��	��o��N��²,6��<oUA����nz�q�x��]*��t+�+�V�Y�|���I�9���.�U�w����s����r=^�kz���4�~��B����6�
�i�o����̙ϝF��mn���2�9�����}�L~oƛi��ϽڃT��S�{^U�N��OL�����b�[�L}��x�܂虜�x�5qv�ܲ`wLΫUCm���;��'Gr���ڌ����k�dƫvE.ۭ����}9kJ3d;�WJ���V>�'�n5]5b��w8�V��N4�MR�����V�[4���̉���ŗtl�\��q#�]}�Kw�QwX�ugj�?}���}_sQ���M���rs��odsP:��U����ƻ��kn�[�G�.q�"��e�<3��2�^'����'qz:b�tQ��#�o O���[5�ju��1����)�J�S��L#����l�f{�^�wP��Ҵ��Q��Q�Ќ([6*%�F�^ok\�?��b�]�q���֨1�nR�Bx��
�>�^Ɛq����b�s����}λ���|�:���2��r�����yQ���|gZ�42�p�g9Ϲ{�ui�w+���]��o�p�����r���{�������Vˎ�R{���2K)Ggp�s6��`�U��7�P���"���=~�>��"���L��}�3�5�M�^�Y��׈��[� ��r� r�[G-No�_}�W�Si� �����#�z,Gy�>w�&�������Z���n���݌Ut�X�b�w�T�>��8"���`Z��M�8���e���?A��ʽ�(AR?����Қ��3{md;��K�<��M\�i(�P7��]�W>mr������\�%�җ��9t>ZL?�coͷ^
�{��&5��S-�:"���v�X���3r<r��5��arS����:{��y<��\��C0��Yx�B�x{3˟�g=�bbY����ܚ�iͨ�����r�U�:���[(e��Vf5��;����y�F�}���(�~t<�|�Kh�������l�{k5�g�Ku�%G�u]����ѽ�WE�w1��e��S��_}U_yԽ=��̛�[��ȓ{�&!��!q`#���t�VM�r��{��,a���}춌S^rx6ɺN�La�W��v�޺�!��U�1�镁^z�Γ�D�}�lf�Ȧ���g;�OL�'�h����h*<�IX8�㝴���*���ۼQֽ�K5����q#�V:��z�t�|���^�`��%�f����z���6��V�k��?��Vbs�]��PJ-ϧ�)���T�p������]�S�e[��d������8J`�ځ��].�C9F���(��.��4�Y��٩�K�@����~mἘ�=s��^�eI���i�]:�w f��<�?]Xhp6��~ô{mm�o7&��*zA@��+��b�1:v��ծ#��>��]��g}�w#�@�|�F�Ӎ�(����)W�{{�&�p���kLO��j�a�Ya����@<���3R�:��]O*��͛����4���]
kB���'.'7y�lg_�[�y4����c��U��H{]u%N����N��f*�jic�tμ��N����vL��X�K�%�d��͓�>��K5��z<[O�+�}� =�˵�єo����s�f��"�/���[_�k��>r3�>n~�1��g�62'�VÁW���q��uU�I7݊��w�:^3���(��b0�~�l��觙Ӓ`e]<�N�Zz#����JM��ё����ם$�mm��v7��>�I�;Z��l	�uq�;%�6Sn>�.��n��0/�Rs�����DDDFL����U�z,�ކ�ɥ}�+��4�*F�������S��G��we��8���|׃�w��$-����ge�������&w/z-�e�u](i����]���Mʾ֍wE��v��|7�GAۧʤ��{hۙ�I:��V"�v�����MU���g�>�7_������I����*dTVZۜ�w���s\�nκ��b+��\�H���\���oR�+��R#�&�y���C��(:�!B�%r�Μ��^��+���a̓��?*��Y��C��n]jF+u��W.��+{Ν�K����F��ޭm�C�	�4�&�Q�@U�����Ǩs΀���4"7x�A�y�L3.K/`�74���SY�Zr��,\��͈$&��rfmp}�g`�zU���c���c޼OL����ۂ��4����R��,fSJ�U>��4�w��V<�'7�Y�a�+Q-a9���<�K���
(�1|�J�g>���`��S��F�w����⻄qq�u\v&B�^�l�w4�Uwʴ��6qʛ�^t�L������ۂ���}4M�b��d�/�����rm֫�ѰL�z�r���b_6�m�.�1�pt�;Ż�:��J���=x#�7Ɲ�¤�Gm�Yԙ�Aq��T�r�">	�Ӆ�3q��pr�o�1�֟e��\˱�)=�u��	*���cd���bl;�-���O�e5oh�(e�:͌���H��;�Ģ�i�ϲ��j=z43�]�֕P�F]��{�����w����y�����:�b-���,Sq��[�-,�λ��6��vI�t6��w.���mjD#gw����E2X�,%�kfs�r�c����1�T ;��V̒f^�񂻉��`_1�Kj�-�-�҂������_}va��G��(.���x2"��箼ۥd��_7��8�v�q�ur�bے��Yʅ��DwT��]�)1���Rʠܨ�e�m�PA�1xiLv�>���(pN��+Q��-4΁�A2�
���8K(��n�5uK�w@�B,E}/M�C��EgC�Y������ԥF�t8�1X�}k�YL�nB�n�j^h���{�z��c-g_<t�ؾY��XHlf �݃�)R�X*\A�jA�L6m�4��ʦ�2h������W��;�]ta�5*n��ţ���ǂ`�D�����$��C���ݿ�{��X�)"�t�%dU%a
�ȫ��H���YD`(�
C-PQH�dPZªH�b��*�YXF�* ���VJ�dD�"�Rc	P@AH,U[AH�YPQa"�V
H�EP�X�EAA`,"��$X���ci Y�hE"�b�`(Aa
��,"ɉ�d�"�F1��>9罹�;��Z��	�\3@?���c�wٴ�\�[n�7���K�I������}�'�����#[כ�*�#����[K�{�3�o��6r��} �����<��t�;�ۋ�u���O
�&��;�5e-"K(L�w(�-���\O;��Y�4��M���%�3��-rs�hP�<=@��7=9�c+[�Y�l���続��u��"J����1�*�<۞��ʚ�Z�۟r���oHӤ�1��*���󬫯>عO]���B�<�p�n@�>���I��65��]���qS��bR�D]�!�;�ji�����|�����\��^��t��B�>̺�~1���P�Ù�j�l�-���.�!Z�B��2���N\s*�$ҏA\�2�=G�=A�
$=�M�5uܴ���ە�7��m_1��x�H�U}_USRl�>S��ޣq�t�uP㜩�k6���g8�!du����[s���3��a��}��q��L��+NLT'.f�?}s�5�x�k&v��c���]�k���)�r=�v�O�:}=HL��QM�z�]�71�1��kg���q+Թ�(|Κy���v�Kޞčt[�{�7�-�?l}g6��Gى(�[��Nc����X�]a����4�:�YZ�6��ٞ��\������{2���g�s���k[���(`��h���QZ��[��v3.+H�\�F��/#��!�m�%;.�A�+�{�hＨQ��i��\f&�r��\�୾R�����<c ���<��Λgp-�=]մ�1��̕�,8�B����9?}U_}���#���ӻ�E<�X<�W'��E�)·����4ݩ���]4��y�܂|����b��ޑkWYne7:CVr���8v\306�7�8���_*��_Xs�J��͍�t��[�IF����;��c�ܮU�P�
uF��Z�B����7�2���'���|[繳kq'*�*�Z��B�����S��FE���u<vj��C�P��o�N�y6`.f�Sz���h2�y�����?t�~q1�U
�k��Vz���t���������w�C:M�{�}*�6��Zl	y�>����U.0���䙒��hA\*W�:��Q
4Ӵ���N���-���\s�}�}��;Rr��r&j�S74��:����X�f���ގg���2kr�ܲ�f3y缐OEk{��Tΐ5�:{�u��/�`�;��'������)��׍�QJ�WLU�<�V��>��^tN�{� ޅ̚V�(v*�"�o&͢�SrR�j��Tǹ���/�<�F�Y��.������D'��jkl�)ȓ ,�.��J�%����#}<5ud:?��G�3ZU��X}¾z[s�]���A�aڕ�O��9�I1&5ծ����zh�Yt2���.ۡخ*�1hJ�X!U�<�)�8�N���i9;�iC�4P��ѥ\�n��f��8�
��H])�x�&�C0Y���3�:`�V1�TL�P�'�f9�Gz`����{��vwC���e�RG�ʯ���{"qϻ���1{S
A����h�Q��ɷ��njrm�����L�W9r���/.�;�7wx�[	��mB���њw����v[���9�U�֑��c��̞����GX�mD��m�a��k��r��4��Ó�f�9O�g\է*	�Y|<��)�3Fg��zf/p�5�����s3��/������U=mf���/el;�]��$��&?NS=���}�={�������#�c1|�9Iy���p��|+��J���I]�Z���X����vm���@�D�}[�ё�{b�����	ě�ۭ>�ʽ��UӹD^��`s
F\U�2�e��lVWE���������~\�oyZj~�!�,p��lՠ�w�������������T���ϱ��=J��k��g,�઎\ϜY'T�l�aI��'��~T�^n��^��}�Nr���Qi�x���ȇ�F^E��u�[�c�f����ԏ�Tw��Cb�,,�֩�I����4qb��q�'�<����޸Tf�^�cZV4�[��e8��\74'R����'z�_BT$�����s��|{��;�CZ����y��Wa�����?R�쥤����JcS�>�ل� ׵��D��F�;�B| �8m?�G,��I��;xif��:��˛��,�߆���zh9r��{Q �/Z���ܥ�w�ep̤0�hQt��83��u+�
�[��9���߫���*6��?voe�ZA��+c�9�F+Ϝ{�B��Ʀh�����Z�ޟ��G��V���lɕ�ft�u���'���#}j��{9v��3���-4����q�޾uF
ǹ���~�t%mo,���{�ry��7�M��
�#��B龾D�� w�;q;|����-�����Va֪�OL�ܒ���ט|)��\k ��
j��Lj-r���c*�%������PR�ۑ��f��������8��MZ��]����VR�����Wx����M�MU��ۈ��ܛ����e7���~}�Tַ�k:��pt��K�pS��Zd��I2pRN޾���c�j�n1�E�U���s^��j:�UU_Ff��=���W=��t�WS7�#����ssZ[�{�%��Vsk@j.�o�vF�ȸ�gi�MM1��
d��]p���
T�f��ɩ��~u�'���r���D�	��*�n�aW�����A��"�T��b�·1����z.�������^xӺ�<�yU�-e>�������Ǒ�KͿL'� ��ռa�$b�X��A7�9�L���h�Dm>Y���QMOhX�X�y{�����(���y{�M:r������Y�'��,q���'v+�O��&�_T�� �!��6s�8/I���t�B�&���)���rq�t���X����S�F��u'ix���eJ�'Vq*�M��e�P����-�ڀ��b�">#&������}�v�s۲���ŷC��|��b�i�uK�;}�yq)q�؄k���wCv���}��/yT��Q�<�br�F�C���p�썴^g<���N�꒱2��=��n�h-\{5y�����v���66C�G:*�%�[q���݇��R��9��}�KC�>��sZ_���>��7P�sS^��w�;�n�5}�+���q�������o2zj��tgʑ\.��|�y0��U��3P�����fڡ.ϥ�m�n�Ryg65Tl�a=F���6���*n� K�A�6�GQ�)t�CCq;���/%iINn�D�����y�X8�s;2]�Ӈe#�]mژ:����+�;��;�ec�dZ��G��ꪝ���{�Ѧ�~ն1���!��C��"�]�<��efz�;�:EZ��o^G�\��ԫew	Z�jo�*j>�P�Ŭ�t���x��S�1�ǤL���w�tg6+�[������4�םq��Rn&��"?*�=P#�7E�zb����5z�%}V����4��5��)V�^^>��SJ~��s�U�_ ���%0�R'�jTV��K��?�R���xƶ����S�7�<�}�Ҍp�C�T���C�w�mB����|�k�[A��Y]ۙ�~S��n����_x��w^��5���qd}h�����i��K]�Wn�ֺŵ0B�p��t[϶���� ۜ�e�sʻs{�L���7!�P��צ�R��Z)2�����k����'���
�]�^G�rչ�B���T;���q����k!��t`�1�S.֨��|����,��a򁼢0gSX@d�E�x4�f���/n��� �t�Qs�VAp2�<Tֺڀt1�T���$ �=b��݈i{�S9ps-����R���ʮ�7od�����.�;9>o�yJ�40Lӆ�;��B�O!�Iº���w7�$�p��Zz�(\��ܾ<��뫦f�\��끶^)+�=#���2����3�y�[E��vwWeШW�՘6�c�+�eӦƨ2�G�8k8�q0��E�v�\�m
ս�۲*�k>�X�,�B!YYZ�W������ۭ���iİV+���-��E={׊Pљ�N;k��WC%��F:<�ꀍ_���"�*�\k��^]Au��d�w D�v�-����Đ�L��w�\���,RMe�ScN1�!ʐ�� �d���=�GF��+T�S�[=�{e����iۦ�9���b\�X�J�6����N�y��m��؟&VH��H�Qf�8��Z�q�},�/N] 켔M��w�M�_��r��;ے�:�{5�e>jƗ��5ٲ�Mܛ���yG��x�d�qsl-����������j��>��"Dӂ@�t��K���>ەw��M���]�A+3Ö��wt��o~X���4x�콭�f�TYk"C����A�v�Wiq�띎�!x`A��QK��p�ԈZ{�<��]���]*gdˢ�i�����{�Hs��ϓjV���s:�����ݥ���˝�����ݔ�X_@.2�����ZU��ᩓ��0!����|�2�,�K�u�k�GX�]�I�
y���jRh���w��d��
Ad�
H�H�R@�&���*�E�`�,�PA`��H,� PD�dP�,�"�(��UT��J�T�-�T,��X�A`j�Ri���U��`�dAE�X�%@Xc* �"�Y��@X�X�2(����ݫ���Ү�|5%`U��{_*P&�4���Z4f�̡RE�p��ƿ���zw4��?�높g��+���q�L��|�w��N�pK�1�*K?)9���)����Y��wOB���y�Ҫ&_˟P�C*VW�o�j�ϵk��evr���_[B��I|�5����\Rȹ�n�v�X����v��=�ц���ܔ{k�=�Z�9[������>�;��,SmЁ�J�,�y0৵ڟ<w�}[�3�Y��/{�0����Z�������CQ�$\�YJ���q��*�ǻ+$��6��~x��n�{}�W=��y�GTw-����Y��<*=P-�����]K����-!�CS-��,��ܺ8�ѡ�2��C�kV�a�Ԟ�F�
5���ޚK�hIw\�C�Î[�?W�I76V��[��q���Y��Jd�;���G8˼�ӦS��=}aL�LOCʎ"���X�Kj�O?��i����9�^�̙�M%4�����s�R���@�[{����Ǜ�(<�y1�-�>�H�Pr:�6�J��m�y9]q�`�E6� ��D���u�f`�U���n�Q�TBLgF�����^�U����O��g�i�Y���w@�Z�g���ގU�TA�Y�X9��P���~{^�fS�u��՛=���R��qx}5�`�b�~��5�u�X
�E�k�՞eܨ��%1��4�2��z��&W��O��������/�X�/���5�e,��)r�6�x��ͷ�U�s�O�X�,5�-nvj��#flÏu��9O�}���F���c�ʼ��sQ��_��2�3����%�x�O���>��V��b��j��ůy*��'e\�ɣ��͌�[����4�����[<�5��~�Z@���x��-b�3�Lv�ީ0�i���Um���>}�\K�-[��|�?cg(����������a�:�Ifb\�vZʉZ�s�������[��g��ǳK��k݌��fY���yAj�*f7�ܮ�k��zҫpUC�,)5�ǖd�?`}�	�d��Z��>����ԫf��#5�aʟ��p�ecIc��_�ov��ٚ�:��0
V�8+�YaBz����o2�J��z��9�go�=�ql.��/	h��(��E[��v��j��U�Wm3��w}B�׺ӓ�eB�K}�ý1�~���{�1���.{!.Ě�+;���ږ!y�00��,UvƦ7��z���OS�#�*�+c�Ɋّ�C��/���ܺ��M�c�(�O8ݬbM"����W������<p.���ۺ��!�+Q���)J*�����E��-����4�㼝u t���~Տ'�"�j�Pk����E̿/t8�|��k�o�Q�>h��c��Rwa=�آޙՉr�]o�O�r�s!G��g\��ݏ��97_�.K˻�;��i��e$#J�W�t��wD�h'BgL�3H��]�g��Vc̕��Զ�����Wv�/�t�u�߀�q�u{�Q�E�/�e]뵢_!ymD�E����SE�~��s�;�ٕ�a��[L���}T�������1���c���S�~˞��VV�l���Q�3�Bm��;����}�wH��m��+Zp����nA����XY}Cvy��ܡ�cU��0�[�Yے4�����p��ڟS��1Z�;�̩-I��RͽM.O[�m�/�1zt>G�]&����r2��k�ޗSә�)��^&���S�(3���Gs�]�֧6�:�A����f�]�]�ja\�2�j}��N����u뚁{�O]b�Vr!�u�v[�bb��n�7����L+@�i��*:�{r�
������C@�u��q�E���A�%��/Vҥ��+bU3i:�mS�Pf����Y9����o�S��:���
�r�o0�1�М�f�����.b73����B��W���,�&��RIw���W����uj�ѩi�wn/ȁ]��>��(ua{���Ҍ���M8փ�`wLi!tnOg��d�WonT��,;?�9rr�S{=�:�����lj�lIq�zm����t�&wBq�ه��r�j:�^6��ӛ��aI=d'k����e���A�To'k�k3�5�b�*޸u|�:�&V-�U\�n�N>c�&��v�-��[V�X��v�6�e��ۏ�ĦE��x���Gt�pm�c{���UR�y��Ht&��b;}�t�0�tŧ�Y̕(%��T��hf6ʏ{�m�f��_����_��ۃ*��3�K�Ύ�e�V�u8y����1�p�rEL���.&�/gϥ�I���z���O\��Ț����cu�E���}ϛ��n��ZcӞ&MnX喲���r$�<�Rn/}�M綫`��O�ێ
ǒ�gP,;��6�X�[q]"ռ1k��b1�f&���W6խ�{��R�N���J���3M'���h��S��wzx��IU�U���.9xm�*Տ��7���2�n�[B7���@g���cR�N��ҷס��*n2���B�x���~�|�(c�/T����Z�4�$E�v���f���B����,�R�1��r�qOR���
R��Ii���ǂ�.Z������F�5�5nw�"��O2��._Z������_oZ�uU�������(7��T���S��*|;z�)K��T�7r!�@ˬ����1 �R�sZbA��yN'���r�p	W��T�q�Y9�(�q��J8�����~Z�#�9V�ӫ�w�_j�YŸ��nA��P�^K�'K�h���ݔk�v{����>�b��R2��[]�1mx���ޖ��9<WR�hS�6���,ǽ�rO�=�D�5v�k�F�;u=��Z�&T~��2���ȇ�ƫ{��0��0A��}�����c�6+/@�}��V��ˌTvic3,�W�ue�$�e��.V������u��YӴTݍ[��8����׻�3�}G���c�F���z���v.Y�٢��T��$�eK)$Cp��]]�iP�� �����S��7��)����Z�����'���Rus8��-R{WF�1�|�l�UZ��;�"�a�07&�J��|��塮�K�q=`r���;m���|���*���v�G%ҮB֪��p��gg3�Q�j�ޅz���A�
3e�oz���&�y�w���x�����b��b��i�Ljb��m{�w��r�1��ǌ�>�I����[sχ��8Q����:����W�VSW��)l`�Gp���I|6�v�1�'v��R�'S+ak�����]2����1�=�h�Mı����q&���1�A�'�:��v��Ί�F�/F��<mrO�s��0��.%m/g�ܠ�ݪ��fo��z�5򏅌1z���(��V�k�X�a��S��7�{'���u�,Vty��E�xo��OL'�
�zrOIKehd!T���k�?.�t���	�c�݇_dY7%^t~d{ڈ��~�E�����w�7�P�,q�]"��%<���o���
�LV��iηczTe�%���;�b8�;�8��F��qu�R��suo����k�أ!���?���=yp�����=C��^���J�V�Α�<Y�K ���$���c#�͔���Ũ1�?+2�RZ�x���-�7�2b�[J��ܼ�*V��̴��C���#Y@��D�gr����`���Ś��t�L#J���)f��![�a�N���jƍ`^�@2�n y�2�2�4]�ֱ������.A�\�WT�X�V�6F�>T�@��ՠ汚.ͷ�*�>�x3����Hes�l�[s9�p��U�	�۽�y\���r;���I�*�p�e���v�呇I�?<uoMfO	cGx6Hj��Dտn����yfm��󼧕sWAg��N�h����K�<�X6s����N��j�t��El�{���Բmm��m����l�a�¥*��o\��:$:� 7A3�q�����L����]-Ժ�tk��Wjr�Y�pNU�趵��;��h0��KO*�M�f��ѴF����u�I�:��$��:���ӟh�A�w�V=�����#FiΝ����9�z��$�a�������)N�Z,�f�t�~�n&(VO+̳���Lb6>��8����w>`�;�*7��[@G)���x1�s�V|�����I�뒦t�S��t�z�]�M�ʸ&r�ܺ���J</7�Rj�˩����BxR�G�zh���a�{^Df�.��`�wdC���<l����X�0e� �>�2S�I��pn���ԑ�i�m��E��7���f���q�Q�{)3n� 5\���ՖV��H,�l�l� �93hF`)Wc��I�>wu �ݗX�)+�ieJ˼{�u��z'1y�� �J����&���x�֊3;���N�.Z:Z�D��nd�z���tl`7��Ѵ�5��Z�:���"��<��7=e� �{%#VDȬ�نg��=q��h�~�s�\�6`,�ET"ŊR��@����`��E�ڦ0+�IU& L��E�bTQjI*AjPQ@QH,�"�
�
����X�X)&0*(LVT���a�CH���j�@�VHTRE��b$P� ��,�j�+%��V��(�(� Qf$�����@QDU������ZR�[8��ē��<���sD���P5��sV�C�Z��W����W�skV��Vu��o��۟��[��d�R��3�gy羍fYIz��:,��*�Rײz�ם�Wws�@���Z	�m"ܾ�2��Q}�y�9<�Z�ڍ�?S9�&�G��	�i�{�l2����{�=��V�.�!�':���%vc�擞�YY+�׺�W�0�mE��V�]f�E[�ynﵾ��`��X���*�>)9��ǟ6�|T�ԫ�O��w!������7��7���~^��k����>����;�jR_y�M��Y�K<3l�t_,���U�R]/�b�"9��_k��uv�^������.�ER��b�dD�܍p�k�U�#�7X*EW.�	K�gk]@d�B�ho�=��Vm8s-S7�Jٳt���i@,��0�7�%��[.M������z�'��(�U��9D>	u6;�U�Ӯ���.b4_K��Ѱ�݋O�.�|��Z���,��|���׊��Sq�RM�u��c��v��[T�XDcK��e������p���.��!�q��T�ˍ`�Er��{�(���֪��'��\ o0۷���X��*��><+�Ꞑbҽ7�J�Ҟ�y��{���Yۖ\+kY�b>A�bM�/z{�Am9֩��Ʃ�Xs��Q��y���==��z�5)�3��HR��Wݱ@�ݽj��^\7��6��ށ�P�/��q�G/�]��9��kk-F�����L^�I�dc:J�e6���u�.ot:��,ͼ��u󴯹O�T���/�s9��i�?!)N��1и��	�?w;��t%�n���TӔ���+�������So�c�2���2��4y���Q��o��]�)k����}C�*TÛ���P��ON�j��KK�P��\~�:�u䗽;�:病g����:e1V��
89�b/���,���7f���븮sS�[�����_�[� ��s[����������˴��ML��`sx*i��P��1�5\遹[��
?>AI���os�^[/m�>�ƈז!����j֮1�m���8,���{T���i���#�l=U�8Y��yT-R�IWNN�eѹLWI��+�Wك�����HK�e'� -(Ҹ�3��,��$�(�f4���y�B6�m�l�rF�¾��e��syh�E��3�٢�,M��М�֡���)����:ØM���㛗He�f�ŕ5V���-\wK*��N�/`��㏫)�p����p�.t��tS���ڴi7�S���쁮�-L�E��+6�i)���HI�{��Ń3�N����|�C��eH7ݏ����9��ۧsk^{}a�<w����rY��)f�pͭ�04[ג�uaT�ߣ�6�{�3;9o�>�Kq<R	X#��v����o�ߤ�/��V�i�8�¹u�6��5��E[W���6,����ؼe��F�=@���㍬��p��n����f��ݐR�-�Zx_�I9������yg�z�=8�}��8{r�sdG.�S���-�轸&17ӗ9}UUN.U�,��r?�7���n�7���3��ƣ��rNyI�b�>�^�T�P1#������1��k�ݏ������9F���͸�\�ŝ�Jsj�b�sbJC�1��|�x�F�x��V��Snʮ�,uUj�*�R�9Kj��s�Mtt8qe<�����i6��G����5����l��7��nEk��.k�i�Όue��>���<��zQ���U֮��q����ʳ]�Fo���Pv���q�F��[|�Dt��B�)f��82=.���۾M5w*+���m��v��V���_�7z�Ҽ	�f�'84�ˋ]w��jխ���{��s�j�[3d�
����+��Irs۳}����ޯ������׭<�d@���f��'��^:>���m}�M牏nU�.;��N�j+��`Vȶ�-t���7�h�/^�5�;L+}�c�����s���of�/j��7Xw#2#!���s�X�=Ϟ��ݢ��{RO8�I�M�{H�=�r����o��ו����F��`k6�Q
�SM�fqoc.u��Jw�1�[e�5� �����=݌��]�.uBK�G�j�x�]X)�����c�	0��5�KX	d ����ʄ��ZT��Y2�Z���g)И&�q�Sf��y�v��:���=u�q*�;Æ�ra��q�Pi4�bM�EG^�-_��o�]_����0Z��=�o�b��O'�g-�݈�2�R��+�W���(�F���x-'�����D�g�^B��m0�[���MS�ԧt�~M��r�~���(M���b��G�*'��s���9�������9Kz{{u�}��u=S��P��E���7+_�J��n���v�����螔w��w-y�9�i?�sc6s����بE9�+]�z�>��*�w��W�2�zN�o�-k{ԠOt��{�TU
>�!�ͭy�{���o�g�TZz45T�N����/<�*��1e؉�/^�9r���k����@z�u��4���X��6y�G�yk�o|���h�yc��[�/i�v.6gs#�v��UɃp�K��]��ͼx�Ͼ���6���q�~�I�Ң�㋜)5t=���#ŏ������
�9o�4׶L�s&�ϘL�m�ig���-��XO�r��فQ�
k3���Ӯ�K9�&j	����4��^���Z7s&�rGb�(��!�u�xB�<�v���>x�/4,�s	(9��{�&�H�+�usy���=�uq��t�N�4�#�ds���A�b\�n5Fh��f)�r�qs
�o���o��就�P�9}��΂>���mf�/HnW�8�+��+�j����0��
[�ʘ=��E���EQ�T�ާ�R�2��5{}F�n�-,:^jQs����٪e]�%2.}|C�a���z&�X��?G�c�s�Z��s�Nw�w�D��Ꝇ��7�e	]�}��q�Tk�͢��-F��w�_���g��_��u��k���Kt�ɫ�f�� [k���s�gP����p3��O��`�/y���� ۥX�v��&Fi��V9�S�G��g`�a���%.��nh�'�˳o��V��U�&T� � ��.��3Q|~o�O�[e���]�q͙�sٷˉ�%l��yRT�3���[����ڢ����yi�>��0�F�u}]��]��1�u_	:�b7�-��5�oyX��T����uz�X���%	Z�;�c�'���t���Vβ�>h�ENٶ����h���x�=��C�6B!�)�W���$�9F�3}],�@�/u��՝�y�Es�⾯�nks��m��^�bxTkT�u	T��aĉ
�Soj�4����F���q�c��[1�9���F=}�M(���a+��ӸEom�U��UЮ��S=ɾ~��������t�d
ܘ3�ȸ�o�
��wZ���W4�	�
R�B���eV﫝 c�~��ұw�J�u���5�ɓC�r���k�LW�z�V��pמ�yI��Ӌ�C�-^&�F.q�b�u���9������]�Y��ٝ;�작�3�n���E�X{��u_*K<��>���7\�Ů�H���2W�+��پ"��!?���k�;���}x�r����[xqZ�Y�wF���)\Y��8��`s�B��m�nu�j�n��}�K����ݹ�c�clr�PUF�	.��\��Ðq��:<Ѧ�s7.���DvأX\w��raLm�l�ŷ�j�xiI�nK̴ZĔu�޽7L7|7\�g�.���a�9�S�h\�S飭��+Z�B��"����t�)VX��3��k����"����X{mB�Y�-����nR۾�������q�0���n#��Nn�q��Yu�kw;��m�w(E���>�M6�-ɰ<Y{�^hB�<�ݖ��ZϢ��eI����w% uv���R�u��:�>t��E���dj�@����F��x,L���h��� �<�	;K��g*�����w�FL2m�"O(�zhV���?�IF`��;&3�>X��f�)� �4�˝W�z�Z��1P��.��;
ɽ(�Au�)[#-�!;isO�f��<uAcCz\C�T�u	|�o���@!���',_^�sƦ�5��k�
��(�-��n�nU���knkH(^ԉ�V=�����]�u�J��ʮl�l�/�E�R��WCM<yH�|�C)m�\��u��ϗ;�H�vi�{JA: � 쓱��f��V�8�ҥ\�1�o`9ш���U���˲��Ɛ���Շ��z�i�CwjL�r..���M�F���ܬY%�甛�oh��,�mn��߮C3-����د�m�;���P�{v�;S,6҂��Yo^R��̋y7VW�<7�e�*9}/�%-��K�v蜨�g3/��4Nb�Mkm�l����Ůe0�֚[4���hu5�*�%R��_>�1V�MmB�����1���ZN��;���^2���[�.!<�y�@�Pkv.�$"G���kf �������z�n���Y��_)/t#b�G(���VY��o0�G
�:9��r�ۜ��dJՂ�T�p�!�Q"
��+RT*)+%�,�D�NXTY���A��X"��
�����U��L�&�Xc�U!Y%�
��Q �`�
����]2cL��J��H���խERT��
�T X�3bM[f+++@�B��#X���
-eb�q�C
�"��Ⱥʲ���|j�
*�2W]:��G7dw��.���˥㕪9�W��BWO9���_'�[0�ױ�F��V������Z�S�s}|gCsܣ�QIbOr���Wi'v�]*-u@��nȥ�9���J��_�!�;�<�Wc��\mJ4�S�K�jz�IQ]^;-'ܯ{EE��,�9u�\����w]�y�*!�B�Ir�w�Y�Am<Xߣ
Ϟ��;�{�R�ŖX�I�#lh�ST�X���%�WyF:�j�n�A���,�!���{���%�u�9������~��!V�����x�U?S�7���Y�ٳ���o���X��o�L������5�=
�Rfn��� X��-����sK���N�L(T��x��4��I�?]f#}Qh=�)�a9m(�qnb����8�5mj7	.���,��E�s�����N�o�����ż�/��7�ܳ&��IˋԂ��&��4�ek!+#���~���پ��4��`~u/����nx:������}��u�w��{{�#{0oxV�U�2��5;b�e��}��U�D�:�徼WZ��X�Ak��x���U��#9s[�Z���\t�Nm�'�Rt�7OE�}E��5�p
����X���rIDoe�}m���W���b��(�#8�#����Q�-��<�Ò'�k�2��s�;n5���/q�W-��p�Y��Y*
�A��XX�fw]�pd��ca�Dw�A�[mb<:9���6ba�w)L�J����ko2��Wcy����n{�R_����5{�������=
�����ק��'q��B뎣5z���Z�
�2����j�G�I�ݮ�*r�ƹ���;^�/�"��u�5�`�}��b�-�9�{F�ݫ���%���:iwan�TNg��y#���g����h~�b�`���Z���Mp��������Uc҂��r4�a��t�L����Rek<����g-����f�Ʒ��I���۟z��#�^)��-f�������[�r�TywV�����1���,J�b���bk��e�v�����w�3�:��㬷]�F������*�y���!���&���g�H1P��S;�b�j)2��2�e!|;B�ސA�\
}���o/Oe�q�C�܂m]:m�ߙ�ڻ�ݽ�]SԟjJ�Ӎ�T%��N3u�Q��lߥ���y׆o��p��3/r<�-�]U���3��K��f'�\.�`+�A:� ޠ�����f�q�J���� �[����֩�ce��RqH��P�iWS�]^ʅ����J��g+8n&{^20'{%JC7��Z�x�R���+����{nIB������YݑQ{��I`���f�w:<;8�v�����9Uv	S6p��?b?���=�׸Ɨ�]I�`�CG�zT?Le���R�\]�;����%��]�� ~VX��t��k��X�k�����?m-�ڝ��3��c����M�2`���؎�5�ʓm�D�S0=���%ɽ���i����ܵ�,-�uy�/v��s�_[mc��xEv|V����Ay�^l�d%��z-�vYs����B���>/�Cr�v��m\+�y\�Y�]�����9=���2��{V*=��{a�ٛ3�W�r5t�1	y����v���#�s�U�[?a�|�U(���kJ�i��_�~j��ǚ�����m�^��j�޴��n��^C�OT�%�I�{�7�ح�e�2��k���nK��Tsun�+���g!~Sf�tQ��"���un��j��3���S쬗}��3��9	��i���yE���#g�|�eE��N��
Hf�P9��y�
�5��>�je���s�5`��J׷�e�ɹ�c�Z�;Yy$qf�=��3���R<��)�^^W���/��K�o�v덩��ѱh��Q�PKRs'�q����J�f�`��{�T�)EM>�9mD��]��J�X���f�mg�?��!��7���q�)�g�Y|#�.hf�ݫȻ3iAwy�;�H*s�}����O��}G���lU�Ű���K��;s�,�b�I�Z��Z��o�!����s�<mto�~���ܽ�5��L{Lv����#*2�=����n�Т´m^X|�����n�V��G�G����^��k�/�!���$�uf�F�WmO*����Ć�s�\�j��7�n7:�q4��1��뜷1NZ����t�t|��n�q��,�oP�:�r�ěC�8�n����{o��d��<����5;5��ہ�e�Y�r�Y!��'�yօ��i7���Z��W!�r��k�k}�A�#ld�u��,��C�[��\{/\]њ#V&'����|�:u.NM�5=��m
�)�m�����+�q����V�u&�`���T�~��W�.~$mu����q�g��8���3���2AZ��wP6y���^����ѧ���\�u���^���a�YpԲ�WMrMM�Ҝ�pQ{����$�e�9����u."�UmLa����keщ��ο4)�[��m�{�խ�����ͥw���/9vi��eP[{5���S�hH�>������8й��0�U�V�#��Yj��"��C⻓��S�gj]$�Z����_�g3Zly�I�,^�b'�rg��Y�m�!�=f�v��f�1��мx����t��`����A�0��b�js��k���5+o�z��q����Lb�O������
�x�z�ӝ*R��U8�����<�i�L]�a����V,�J�G���ۼ�W5��;��ʀ�5�t�9Q���?�M�sy�������T'co�X��T�r
�)�ϓބ�FY-�K�U��N��8`�d�i�41�q��q�׷����G��<����)��p���t�!Ǿ�����#e+��[]�$<��m朐D5K�-]`�{�R�\*f	˫s9K:�v������]��qU�H ={��u��M���G�W����٪\*�4�PCj���[[�����,	���V� �!�`(e�t9�y�ڥ�q��́�?Ը+tP��ۜo����g9��~�=����G�{��bI�����ų�8�{1xP�K
��諾���e[�ܝ���(G������J����m�s9�xc{d��`�՝P��~�h��c�࠙��m#�Uh~u�YЩ�Y����_����=�S��[��8d3���e�&A��M�]0.���ժ���ָ�0���Z�k�Vw�u�Ǆ��� n�u��y�LSv���OoW���Z���Z%FeD�b��d��s���'��Y��3X��+�f"��%�Jt,0���TL�ܠ���Se<.zM]؍��]�;x���YgrPΰ3�����ޯ4�b�}��F�(+L;��e��;a�R�7�5�g/X6���<)��:�8��+�ҳZԻN���_�jԗ0ƏA����)�N����zpD��H�wmOz�Xdz����>�Tk�Q�����
TOeE}♻(y��f�-/z����l�vg�x�"@߶c ���RAZ���wf��卣��5����>�|\@�B�4_aрI��ș!�-����w���f-��a�f�2}1L�0�c���_7�G0�{�w�~�c�>NlP�B�ҁ������`	e�o��Kkx��K���������)�q����0��:K=��a�PV~^o����N&#�bv��?��1�jeE���3����Vqdx�>K3}�ǀ��ѝ6<�F�Fܑ?q�򛈢�ɘYs9�}�a[��Wz�<�b��΢��7��s�b�
vxh$�ވ�Fz��/S�:?�iM�f��]�3���C���v攴<���lor�J�h�t�+���f�q��N���������`a�E�;Yn�c�T5,�zvG��\���1��jv�nӅl2�Z���.��f��@4M"��XU�q��w���hł�iui�+��+��ԎM*7C��v�j/��}�V
�\ٺ���t^pv#�5�݇|�֐f�{�<�ݱ�%-�EI�'���SXZ{fT�kc���5�S�z�
�X�k��!�{K�\�nWLj	x�]j��v%�w�G���Bٍh7v�Vq�/����@��
R��F~�}����c㩴�^�3Y�;`�*n��R���d�Z���Сj��җ.��kb�n�
\V�Hm���e:Μs3%έū�����#*��&�8�aܦ��}mo^EZ��7��e���+��F7p;�޳0E���G��|z�c��٧�#��a�m�x멎Uɬs�0:�(�gfᣛ���Gr9�.�5��'v����ir�Ct��{��������#����˖��f��v��A�@�͍������K�ܗXri�#cWp =%��:����Cq�'ۜ:[��Ǡ`�H�6���f�q^<Օ/�^��;��� �:�YE��+o{(J�%�F���P��%���Ũs�:��i|�WU������]�U`[l�����="�wB�ɼ��k~8�l�`	�v�5*����B�f�45������]�s�+���)q5.ZՇH���%�m':�=�c��c�	�b�&��Q�k���{WI�fX|g3��y�2���X=���(�-@��֤�I�Q]t��[�evR�Y�ˠh�l<�wz��$��n�����v�r��d=;�P�|�-��u����q'9ϩ�糮|mڀ�P�^�@�X
QR��Y"�/)��i��(J�E���%"�)�.P��`�9E+*VUh���Y#HVf&01�j �R-`*�Reh)���J�՚`kY����QB��J�eT̳b+���P��. �D��m�R�Z���U&Z�)P�[H�MVc&�1�f%V+*,R�����"��,U�R9`T�!X(� [j:��zߴ)���N�,Yȸ��u�ӕ�]�o�X��O��0ݷ�CKnJnv�:9�ީ���5���A/��)�|�ʬ1z@<s��?{8vg����;�U�LT衣�\�z�,vH��8��u��w���6�{��@������'��L�Pљ���s����Qy��I��^��|�~&���)�.�/�YU�����cff.��[��/#^��,*�a�ܑ�P8i w�B1>(Y=�����9�//CE��^,oʡ������c�� I�E����5�׃Ў
O��cӹT�0�T{��,�1�(�<�)޿P��Az:@2x;�T`��	�Ѳ��{���L�	�U�|�g��L`�>�S[$:(��xȎ�a�W�>C������z9����4v&9��W11�,��b~�z�e�����[&^�xP�X10���?7�:]����k$�!�����MD==��]5H�̭YI�����#/E�J�J�]�\�z��F��Z�g�p����&<��}�G�@��dCe��RD��r9��髪�q�ǯj�[�$��FU�{T.X���۫�\!W�~ u"���Z ���.�]�&�^�S������} h�tE#���F/ﺤ���Ǚݮ�ެZ��#�ȑ��=�U㨝�a�>�����R�;��O�W��FT�r꣧�e�ɖ*΅�����P�'�z�ќ��U�Du}�q2�L�:�W�w��=1�b�ԇ���P������}ʸh�%z�z:D�'@�s_�Y��1�����b��]޺�y9��0]וX��qB"�`����9�\��3���ysB��3Va�=86#B�u	9R\ 8Ê�D������Nǉ�u �xX��:����Pcb��M��4���C*X~QM˟�����&�L9�����4.����{8�!��b�]�\�	�+S/�<wP�U��L���06H�ue�֕�:���V�z/jdV�M<�����
F�h����@��9ӎf.dϜ�{���~�ם�3��d <3���g&'�X�*c���*�c(V������]>��x��A��U2���T��������#�\?@�}��:#����k�� �1�\��q��hB~u0��G�8����[��>u�
d��0D�G)��RB��Oc�UV��.=�t��ƞ&��'��P9�S~R����@�F��^��>���8E�w���r�e����3�s7�L�z�m�W�;�z#�M
�`9��jw�Q��1�������:ů]�w"�^���x����Ŋ��ՙ^��z��LT�$F]O��Mn�H�j(?zc���b�T����#�EV���Lh��ߴ�_��B��X�;�i�E�ǗX����Io����ye�0���Gv�m�;�����u�<C1��=�j�J���Nh[��TEa^P�`)۪�����m�#׷y�]8�>f���GC�+#���/=28eM���{����@�9�5f8O�1սQ1y؟��1�H���E�ڗ�<�:TrT�D�g@��1��s؊�΢���k�S���Rf_����1�a�/H��� �W��W�~���2�x[s�@m����{�	��o�?F�G
��#p�9��{҃'D���=8!w{����k�2��t�ku84� G�Pb{&.<Pb��jߐ;��o#{����g3,�(s���ǽ1Ȑ4��#E똫ɹ����]�C�7���k�LLc�*=�x�Tà�	����+UC�S^���GyM�e��(z�U�*����B���ag��Mg	�}�߿(~���к6,T{��8a�~�\xs06�N|�Ï?Y�U��D�Օ�+�x�D�a����@В���a���g]vܙaӴ��w�[���tj�о.]��v9T���	���(�JYه���y�qz����u�>71XcD�4u�7�(�U��g�B�e������PX����;�u�TU��Ry�<Wc{����?���0/ň��)o,���i��l����b�a,^�&�Һ|�xa15n�VN������ )�����sL�Ws�^��[qד�N��`��P��9�ɉ��y��yY��L	��,{fX|6��s0�=,q�����x����v�5���%���:7�`���(�ʏJ��=��������h�1S�5q��:�VJh��$E�G��vc%歪t%vw�z�y9`#�lO�v�v�]�$	����s�aP�ӽ��#���P�`Y���}
���,k�"c�(��m��®�<���~QF�Р���n*����X�J�(˳��z�j�y�o�]ﻱ}_H��0/����kuv���Uox�=Ւoof��l1�c�w�o��L1# �"�<�r�%�<� /���HH�v<m*q��#QBč@�z6]����r`�s��{����k}�=�Ǉ��1x�:�_b�B�M�a�b������t}C�2?l�
�~LW���>5^��#�ʹ�y���1�2� {#�"'��Z��.Lr7�:b��ͻ�_I��>��Eyπ��+�7�*:a	D҆�&�LM�}���3��g�/s�<�����i�F��H�I"Fk��~��X{�^�`���JhM�b��Q�E�c��,!\o�x��{s�Tzh�u�ZC �Ӡ�ۮUV���K�Y"}�Ã��uSg�/��z�b��*.&xԜ�N�w�E�ǫ�60w����������{�.�Z���ۆ�鹝Y�(���=N�]�ʩ�Ƒ���� Q�RՉ\�˒ۨ�e���y�t�He�����$B�W�v�3;�V���e��3:D�4�M|gd	g|]�j/_���H�o���f�W��B��3����"�0!�&D�������jk|�p���;f;T�b�N=.a�N�������g<��Οvo{^�2&	�
+�>���_�	e�厯�kW�J;��.>��p!��T�,SS�d��vyǼ%z������ �s�k:�����Х�XG��2�ϳ|�~��N}*lp>����1����$1C�l��lߞ��B�1̞9� y�c�'H
c'����^�ne���{��q�>�f��8$|1*��Ω��`�l�	P)l���5��wy����"��&:�q� 2"�	ˆU�-�q�슲�A�?�
�w�����qπv߭���YhiX֛�e�׹��EEK���ͧښ9�J�Ǹvm(��缰4�Nu�����x�.��M��ڹb�3��ޖ;T��L�qc�� �O���������a��S�N���s���y( ���5���'^����#B7lL`�:��PQs9�7�婻�ɮ��4���&�h�A�*��� Z���3o�7��������[�}��f���7��`a�LLvJ�.�,��8�:��_����/Ƭ�	Nc�z��#C<��Q��	ʜB��8�o��*�d�L��,
s*��b�M���:�*#oc���n{�}��A�0xL��AQ<)}�PX�ϋ�r�?P
��?�����UJr���?C�jцo�Wҽ,a:(pj� �����{�4#��
;:C�{_7pÁ�V�#��A�옝��#�~�4E���w<�@�gZ�mu��bay�� �����z䳦�䲖CR�h���ӮɎ��:9(�$`�����]Ņ��9���QR�	�\���@���x�����ͳ�(p��4�����2��LO) i��F�{��6�W����$z��=f�	������D�p�@�������,x�ţCr.|=Q
c*f���k�TèS'�0���<�������-��[?���`����6'�6,~��w&���Ǉ3B�\쵧�;U�G�F�r�V�1:W���VLh��MYa��u ��C�}��=�@����bc`ȱ�@����ʋG�ޱ�:��~���8��S��=�8H�#~�8+�"t�yM�^=�U��������1�c&b�-T1��SO�	NpU�WG��k���K�p>���uG��3�:#��a|3�p�r7&$�@�����yw�;�^��|j$��L�$��tp�c��;�SC�}re)��':0��oM0��cm]|�4���Z������5�#�$љ81�V�O�ï,}����L�D��Hǌ[���bB���^�yq�����W�珍m!�	��4�����`���Q�OOvU��<��5������H|n9��B��>%4Lt�tȉ;��^.;4g�Dnyέ���_�S7�}s��	$*:�H��軏2z�w��4<Na�${��ɉ��A��L1��0�H�҂'傫�T�/C�NN�H�'�j<a��R6K&@�z�ן�,�}��:${�4L�+d'�	3W[52c����]Z�7��;��ǻd	�<LK2E���Z��#E��?&*�:s=^�9�$�z<�<+�G��덂�ƞ�D�*ub&*�&3��>���U���g���=�����BŏN����8i��GDu�G��`�^4���>GG��}�� |Fj� {�ի/W䩽�B���טEv$�Pܩw۪��Imi���0��'�q�6�T�<5����G|�6K�.����sp��`�3Y�]�pR�� ��/Z�W@�bZ.i��F��6ɮ�P��C��ש4�+k){N3��n���7;�R�vnչ��H8��q��+��$�j'��%�} C����X�h�RL�8�J�Z��*�&�E�C9Q&�Ж!��|��[��P|6���]�ͬ�p���q��g1�^nr�s�Dȡ�\��t�^W|���j�-��;;NS���5A�4ɪ�fj֍����㶆�p��K���;}��z:���B�ƴ���>��L�'�N�R�]��K��8\Pn�b�kY��.gA�07a�Ά��a�SZz�H��w7���ҾL��$���Ƴ���iݑ�x-��{�x����޻��m�ƭ�b��7b
Φ�[kP���v��$ 6��L��:9�Nmm��9��-�ݤ�t��ݚ�j�j�z�'l�i�3֍K����)>/wá�4Lm������3�pu}}q�-���Tmq�[n*P'G���h���Y���Pl���W5,�P肬wA��:b����4P��YYۛ���'ew|��BDU��}c3��۴�m���Hٌ�.
ȶ�q�GyW��6Mf����Ʒ�|�Sh	De�횀g��&����0gu*N�9�@�����f0���,N.�L�T�O�oM�B�t��'�"mXh}�y�Wt����@�n�-��m[%k�|hwN3--�b��Aj\΄Sq��XY��������� z�VYt�]�,Y�p�u�K��m����W.�c�A�Ӷم����wy��gX��LQD\��KZ���t�<��odr�0���vHArU+<�K�T�`xF8F�r;�.J[wv��
�EU�F��0j�MG,�U�)�*`����R��QaXVAU���E�H�k���b�R�(�Ls,\J�Er����b�Y+�Lcl���YZ�ZՖ؊�8�(�D*B�k�E]$�q�m`�����V,��,B�UIQX�����QT�c�Y��V(�q�J�m�Qb��\I��F`�,"�U�2���b�Hi1WVV��2)YR�(�+����mr[�Ȋ,Q��b�1랷㭸����x�������F���6#-٬�����
tk��{g�Y;�)~�/n=q���p-��1�@�(���fل�gff��:�eV=~��64�2$z�0���E�:�!�o���H���T8v�� E��_���u�7&|*΅Q�"p���������\����tOϱ�_�ة�ZZ0x��j~4����ү�~{�_����o�BӃ�x]C�f���_s���?b��F�ğٷ��˝��F�D%1�bx�W���<5l��B������:�{���]QH��s���t�`���+��r�gF9��xi���X�z=2$�:����8���xK(0�Ѯk����K@8���3�js��2	b�p~1b��ӕ��w������#}�O��N� �Ɏt�190�b�D���D'������~ey�}qŗ��m}�m7fם�<�z���y;Z�?09�a�����_���i+hjPi�(��M�u���R5��z6X*�ٓ7y���RC�=�ƌ ���_u)!��x���^���3�=�
�Bc,������ hY�\x(��3N�=�5�Q?qXL����T�Jd���Lw11���z���߼��cǧ���m��>&��k{� �e3�1���/w��^��Y1?'<*�UFN��B��x����X�����09pյ�����H�{&�_l�"�����5�-g�H*(/7�o�O�ٳ�Y��R�gc�1:U���9%����!}{9�ג���U�R"�}P��H�Q��l����=%4f�k'�_{�z�tY1�tFny�5�<�1�X� 	�-������ע�̋0@��}dxy��Ψ����Cl�m�L*u~����:#BM�U(_>$��W��Ʃ}Y��)We�0@n.��t;�ǚn���kXٰRe�L��},�>��P�}��(٧��R]�t�v��L%�(�1������	\ʾ�PܽIB�����@�lUA�(c�����)
�p@�u?L)zךv�*U����u*�xǙ��Lm���9�z��=�Ǹ�S���U7,�.���U��K�+��G���ca`>��^�K�/ztC92<>�9�5��vR5� xJ��s����g��g_����ǆnM#pK�� u}�TL'$1�>W���9����XA"�I��1XU�T&����P����z.��<����&3Mm��_�r0���P����?O��Y�6>�ջ[��B1�o?|�D=�)�4lX���3YP��z��3	Yƭ���$�H����qb5��#F���p����~,o�{=2�]Ug�����3:c�s�T9�"��X��C�wZD���w��5�����}�dJ��y�	�Z<Í��](08a��~�cwi, o������<�1Ie��r��yy�^3J$o�>nn^rnv�Nu{��d�����w�	�4�
�X��JpWX��ً�7S���d�G����mTm����,!��^:�Ӭ�b����ŋu]ueA����
v��^��:��=�b'��o�2-�<3�h�wې�ע׬��t[���ud�2�u�p{Ƈ(��O�W�<�d�2�����U���=Ƒ�ܙ��$ cꨑ�@�w�vtC�J��m��dB��T����6'��\s��`����IG}Qn{=��\�w�<F���1���^8\�b��BM��� 	��<�y�G�
�B��j�/a���g{
���,2\�x�ڪ��_w��4z�r�N�
 w�{&d�5�H����^�~缔c�,�����%� 8��2���&}���OA��x���?��N���O�q�»|1�p�T�-�]Z��[�%���ǜ�V�E�ƫL�($3\<���g< >�s������Ii��Z�s�?��Q�����ת��=�I�ʵ/�Z�;�����I�1�@�����c��CF���x8���F������$�[*�GC20����rP��:�����܏luC�a߻u��h2���J�I��@s2#�c>�$:�<$��g�}����=K��^�UgGx��� ��/��"2;�
4(n��
���1������p���>څeɰ��O����)x�5b٨�0kZ��s�޽���z=RE8�9�5e�/�r�i�u��nKw"x�C��ǫ|��L��ࡄ��zl��s:�N��Дl�ӟR�t�ez�/*�=�x�lvLZs����5%i53�MN��}gx���ʺ�.k�۹�]��P�/O������7�u� ��Up�W�כ����[�=��$v=�\�-+!LXU���8��~p�Ş��ʮf:1:^V�۟���p�Z�͢J�c������볮�g��<5�e㕝-�������= ����̝�	�ݿ����A��8�?;U�حϧ<�%����uc�w�ݧ�g�ܒ��w��c��:�PЯ%����<Ϻ�/�q��=���b='G�U)0����D���4N�<}��n1���"�)�A��5�K_�<� W�R B�|���g�C[����9�_��bu�3pJ�$1�{� r���㟺��.�ֵ���K)��;���_u	��%�x���� hYᐝ��e�6���h��-TpXL�����K�O�|�f�u0/lF��כ����#��LpP���4md�2ǉ����G�� @2n�1�auZ�����GI�G�����Qr�a����ħ0������j���q�������k�F6�~O_��3�?�1�����L`̋R���i&�A+�`�S�ht�[A�u#�m�W}srM�/�Tn����Mw
�y�ky2ЙG3�w��p�mb�w�j�A�X��"y����mJs��/�;hb8���5��⼧@��S�^�	NpEGX�Ш��P���C�y>T�}���8��G�a��ڑQ�����#����E\D�8�C~S>v'{s���\z�2X������C�8�x1�aYb�kZ���:��N�K��&�f�o�,O��Gx�#�}N���Q�lZ=����:�U�\4;�`���9L�E�����F��ނ��u|��c�|˳[J��:���)!,U �3���cq�y�g��M	�D�0�g)�)���a9f�t�@��W���IC�WUޯw�؏���8 Q@"�mT>�w88�;� x�;t���y��FWLz��=g�X�2�F̱.�:b=ꉄ䀴ߣ�ɾ���oʽ�dh�R�E}ųU��BaV��Q�HĈz��ಇ��y���1u�DC�g.?ja�A^�6wAɭ���
=�Z��ڮf�N�jg������#�b��ڜaA�-Ȱ���z��F�=��x�h@�sbv��-���a�3>��w{�Q�������^���s���3�Z 1�lX�����eC1E\a���9���H���C�_~(-��<-=��U�hL�T׭U�N�M���/μ)�bG�Θj'�P��	´�1�L�oyG���uB/V�T{нΨVz@�{_f�|i����r�JS���w�����.���翫�/����:�����pq*��t�b�V�|�ckڟ��9ygzG���>�*���޸w��L\Σzd[(dx�;Q�]���O�}p�5���;@-.�����2�������Dz|9l�m�v���x�&�6�i�~�m�H�b~J��� S=��~}/����b^Y�/�tD��p_.�V�;��*�TJh�Q3"/��O^��(3.�O/�n(D]��=6�����������8ƽt��L���\�JV��_����v$����+���H�������x� ���{,�Ǳ�.9c5����榿G���/.����^8�uӨI�P�p��≍=G����|"����%	��^s
�*&<�v��r�Ͻ��4�&+n<���( ��� S�X> �|!�̢�&H�*3�o}�Jc��$-U�]�?� Q�B���,k|u>��ީ;[���wT�QG�4�yMĔ&=��&4,;���u
jX"Q�W����x�y�&=�z���|*��9�68`�IՈ}������I�۷�q����p���.�xZ�>5��"9�7\���^q�y�w�����]U����.. -�8o�z�qU����I��=U�� ���&�1d��_�P��D�q�-lh�驺��ג�֤zlǽRE
�aT·P�����caƙ�`O��8�"�m!�5�-O��v���J#��r魙�l�t��j!]v���"�˽���>Y�_�QZ��JQ �x~�`t�]�;n�Xx:��+��o�$%�]���mܼ�n�tءD��vf:�#��L����bS��J0h~�O�����G:�.	G$�&�g������NY��Ow|�֏��?\*�ņ��:t���q�	�:��{�����X�&�7H>�1�V9��/�U1�b����}����rGu�;��~��|0T�9�qXUs��v����aE����t�ޜ6���.w}��2}`��j	aҙO����e����>�C!{:��m~~h�!��G�������-�0az���:D�<�G�FOw����W����,��,zo�Q�r ��/d:�����O�{�w�y��b���b�GI���<� �	�=8$���Q�]{5z���5D!�r0�N��x�sސ��1%��qT>����}O��.�bh�����ϱ�?+��QwshZJ>nżG�l�t����F���j�8N�L�u��* �v��v������WYJZy�HMR|Z�+F�u�������m`�z���p. �c��-����a��{C�o���� ���*�����{[4N(4�B��,������碙Vk:�a�V��^�Yװ���RU�����}��^ʏr�����|�%z�NnZd�w�eB4v���=g2��52�c���g:��]��ލ��MBB�ؒ��p��89����{�T�3��4m�F�����p��}J�o�r��v-�tu�X��2
���l3y��/j�;zB�r����Ǳ�9+��p>w�t;q7�v�E�m�y[�ZJ�p���#��f<Kk�����74�ml����z�^��՞8k�z��;��%gN5�"��,�MF�9�})[յk��ܮOh�`;ܛ�@�k�|��}��'x�V1�J<���:�����֞vۡ�tC3��Q6�[����W�5�<�`(�Vn�bٿ*��W�ˠUtRRT\\5�舭�j>�+ii���V%w0��.M3���m�vGM���E���+��˴pl�3�WI�����V�[Օ�K�����EY�Y#4����;ó���%N�ף�#PA�&��#����L��ZJ�����oy�
z�5���eq\����+36�Xb&#㹊���|˫�sb�x���ш-�*v&�!�����71�Їe��}3$r����BJ�%�f���x991Ԋ�.t�q�W��mo0�4L�N���u��@_e�ъ�[���wbkb�T�	/�aN��X/jfA]|b��}.p좞�m9�V�˛5s��t7}���[4�]��l�L��(�	����}:��A�-�'��E�"�꽫�5q���a��r�2����#nqo<=u�^\����B�Pb"]f(�A�+Mf��e���2�E*Q�m�&0@R���-QPb�C.e��33E`�3(UEY�TLs
e((k)1m��GIEPQQTf%�YR�V�L[��V[dE[UQ�m�+W%Llb�\jc,J�Z���R���E�"0F*1h�Kj%im������J��2Ֆ�UV+&`��Z�Q�DGHڨe�FZ��[���`�##����UF*�ppE�*��PK�`��(eTY�R���@�:���@�2����N�]gc͔���%���ܢ�v��f�rR�d	?+�ڋ�Ga3�uƾ�K	Lώ��gT�N�ߡD��U����FzƉ�s�
&���<N�uz��X,�������θTiD���*����r�aa秸��E�����_��P��A���?�կ�_���b���'EW��1Qjw��s&������zs�e�����èSc�|6#��LN�d��*�3N�;S>�����,���ƪ��u��b=��Z�S�Z0\3���=�=��e��O��I���%mC�KLo�F���HW��H�c�¯B��x�c2��m�L���P�*��l�'ʃ3K~��<�kC�m�����w?G=�J�Y�����@ލ�\�ƿJ��:���O���]���_(��G�UE�G>uꎸN�!f
F����d��W��nk�{�4��5S�x��~JZQ�S��1ӟ��m�ٍ7a��_������mڱV���GA�V%�Ǎ��^���˒ܭ�%������"��	���P����p�j����C��ƒ���77Pu��C���w�:��ܷ�O7}ݜ�v���wMY�UpD��(�`�0���p�80J��ƿUe�ז����zcG�����X�ܚF�c��� �zafPu_�'1�w�|@�Ll�#F^�ĊE3���5
��k��H�,��E�2��g�{��H"o��2���s�S���UCU�{���s쵾g�vc��
��z��&?#�p�D=�lLQ�b����������k��g��<3���,��P�@�GƠ�»ڎ|�W���8k��k+ݧ���_ST�1]r���*X!qc�60�9^�Ws��s˖�0�Ǯ�^sa�y����SXb�6,E�X��t�Ǿ����r�|�2�ɐ�\�:&��C��f.��N�e#�W����0�s$EPH�@���Ԋ��bVsH|tᖱ0^󙕶��~�V`��Wd��5l��ݲ��E=f�w7f�}L��V������;�����Q�=���#e�1��T5��Y:�F��K��d�'ї3����1�nW�q�uh��қ��ō5���;|���w��+�P�hg��<#�#r�΂@�zf� �}��5���G��HEq�0k��0�O��p�3��(s�_O�U�f��݈�G�*�auD]B��+�P�f��Q�u:}�w��$�^2&
� v��1��<�U>ۆ0�T1���N�S}���v(�G�(��>�%b��x�ܙG_�UFI��=�����"G��Ncd�酦��5/�8�i�d�K��4��כ�Q��Q�Ԃ�x��x�bx�4jc��B��`��]����׷�/_�9���cx9�����0�B����&9F���#�j���RW}j�j�_92���Th�o�����g��V	;ƼCZ�y���}{�B̓	�,�I�:Z��Įݣ$�W[C�u��À���amR�ݎM[�8?;���ʞs��]B�K
d���uB*bc\���ε��K���=��c�s4X��>�zm]0@Qj��!���qG�y�
��4QɊ��X\����N�6#���Y0P�N=�mo�my0fTOT�B���t6g���Pzd]�:�뙗ݱ���x!i��U��OFX�̮(��ɟ��ݟ�"5:����"�v�옷p��%��<`��Y���^W_-�Ho�L{�<�}��~4�X�*�	{�1�N�9��&���?5�s}���ŉ��Gx؍��9�QʢbԱh�x���|�o���p�c��kq�zt�C�"~=���1�j�tƪ�^+L\{ra�UKM�{yݶ=����NK��A,6H���������ܰ����ǀ�ۑ��6� &v��"y�3Wϡi�t���v2���Q�;.��9��\&���m���[�FD�Ӹ�+�.��9���Ob�\���h�>���a��&8>,���Pb%Ά �7[{:��z}�������Iz�2��H�:��2 V�&��==�!�����W���~�B��vT���s�_9�,L{� O!04�[�.f}���{�W�%?)RG�d�� �{�>+��3@�*`�d��/,`/d��F=��	���L�K
d��0��q���u���^bc�H|cFA�����#~,x���ǱP�rig���5{�l�>K����tt�����(V��r��e�5��}�c�����A�_��*+����&,m�'Ex��t�QT���^H� c�uFi@�Ο;��pD��QZU���f=;d{��w;պ�y�}�:*�s��n�E;�9��Z:�r��X}�� 0�-�d
?�5�~� D�8V��+w.�%���W�]�m�Ps��Hq�%--�{��E������Ֆ��9�T	�.%�h��R`v�-7�4����*b�}�I��A�@Mk�w����k:#w=�bƣH�aZ���&Ono�Z�{g?�Ί�����f�e���*���_p�!u��4�>�G����gP��\��_��U����/��=]���~����A���I�^��H@@�,��R@�;���k�]{����_�ُLT��L������ꡊn��X	�;ݝ�9����?��g���^5g��zp@���,aT>s8&�ѹ�V�k��� <���&/������Q�%�wX��'�2}棧�Fz=$�>��1������3�eH0����'�my��d|�<�b�D��:4WƦ2���(��MaA��,?;��H�T������s���؄Z/�|?qa�������ª�ʓ��Ƒ�vV�lV� ܃*Tte��u�[��љ�9Z�q�}|�r���M�0LP+9��m����Ŋ.���%Y���喷���]�>�"o��^��^��3,Ș�,F�c����V��N�)N���m��\f�3�ԀF|c��7����%t��$vq�ױ�p�&�2�㩚�����������������b����sY�{nH��������ם����y�J��յ##��W�佼�������9�V@s������=7޸w��L\Σzd\X�t#�;�\�z��z8�b��k�c�^E�Č튮�x�Y����A���]3��۳袧G�_��"���u�H�_D�@�L�^l�Uf>��a�=����|#x�,_}����3 wM�{%�^w{]�虑}�>�auE�!1��h�O*\�H�@\�ǫ���\l�@��#"O�
'��Y�F��
�*'�9�_�=��?e:�g���
�?�a�gc{�3��a_>��f&���|0�U�b[�B�>��]�ͦo3qK��s�2��aҐu}���-d8��+�(D)`�QښN�Ǩ-Y�k���T���;�Rj��Fz\�eN�
'��d�l�J�����*iAS�$\G:}ꉄY"\��PJJ@���������F���ś�/�b��0���'�}��&/J�$�n:�}���,����z���`���$������Кs �%�;��3N��nOSh���5�m����C�,�D���凙^c��~�G��8=�<!m]U��u����ك�7|y(�~��^�Ȱ���c@��T.�uB�=:�@�>V}�r�r�<}��)�8�D�I,P쉝	��A�1�/"��΂u�婭�My�j`+�x_�Lu)�1G	�Λ�ae�����o����b7�31�q�i�2ǫfFa�Җ'�bӟ�>��F��'����A�עv�y�n�K��w�G���x�U;fI��<]�gS��إp��=mvL|�B���v Pc��x�lͭ���8i�H�r��A坎���K�|�i���l�ծ����(Tx�v�C��|��K���~m�^@@;��!1^�&(�5c||�.SŊjb����j󼠨Y�^�����(�B���9ڭ��nNx?U��V5J���c�M���F�r� 4w�PT�@�M�/_&��gX�IS2�҇#RP�7T�����t1{/fc�]Sy~��	���6pI6�1eO��E���\y� �+H����q�vU�����M)�-��b��=4����{� �B`}���+��v� ��Q����tD�x�5�
���ϼ@^�3<~���j�r���@��!F�Q1V5u	�Ic������^�mU�y9�	,�^bqI��nxz̓k�|��<�`��MS�tfl�=ȉ��bt]�qp��OC-��W'�, f>?_�v_QQ��#�ef��9`�@����ϙ�*��-n��8��}[����;Ц<?��?P��S��TmSx�GV�<*���c۔��o��˔����>08���K���B�YD���E_7�ܷνHǣT�o} o��2vP~�å6;��!9�@��n���D��}�؉S1�}�,T\�3xcz�jD^7Q��P��pXjj-Z{����9�3�Q'Í�k�VbQ����!_x�%�H/\Y9�^�Zđ����R�-u�̪���Pfiʳ#���:r�\��׳w�(q�8��fx��e�@�5���uPbT�*ǃ��҅x���w�x����|�6,��K��Ψ!F
F����FO�������.�����68�|0p��7(;��bS�n;��c�w��3���9���BC�?�OJ_T)�Uf?��?�����������?Z@�@r���HBH���P	!$�~�.���L�B�Yy��C&��=�?=M�xH��I ��d� x�����Sn��h�P�'(HBQ�� �HBQ@<����t'�����`�/t?��dFc �@������w������=6�?���2x;�g�DO�e��p{�&��P�D�D�{��C�s%���y���y�����?�؞~Sp��*#�=�"pm�@�@����~��5�����A��>D�����x	$��#&9��]}��P��H��> ~�Bq?�'����0C��G�nI�)���d	!$O�����0Q��a�``�� o>�Y��z4�=�P�@~�6���Z���A�������������`}{�nS������dHI�ۻu�=�?��@�C�8B �  :eR[����0.}�C��p������?����$��<�xM�I}�s�}�{I�����y�$���� m�1��=��p�?����m�����k��?�?/����t'? �����YHIo�P�c�=��P=7����>8z��)��z���P�8�??��>�����'�.����'���=9��y��!�����?�8=��$$��'�2 ���>���?�؜�&
q(w�hϦ��I l�@�@���H��C����l[!��5��d�������hP�������H���1'`d���'�9�x$�$�=�� ̓r���C�{�xl�gg�I܉�V�����	������)�AIi:8�5ɐ���	!$�`}~��}��������>!?�$�O����$���O�<��@��=���=@���=��������>�G��>^l?�`��|������$��=��z�o�=_X_�B�>_w��?a@��dd��
)AV@$$�I�nO����$�:���<�̟?�Ȟ�;��&�w�v��D7$����C���4��>Gۇ>�� �}���_��~Ӝ��D�`�P����rBHI����m�k�u� p��3���	��OC�����{
!�N>�﷓`4HP�I�!���$I	!$�"@��O�P9@�{���>��{gN������y�'�n<���}V���,F�gې�367�C���a��(�Y�����)��O�