BZh91AY&SYzX���_�`p���#ߠ����   b;=�  �Q=���CF�ѥ((� �m�)�	(e�T�3b�*� *���I� d"т*U�٪��*��m�J� �%'�ׯMmD�Qg�N�m5��V�Km��hV�V��T֪�f�iU�0�ڶf��F�m�&-�����V�5F�h��UU�kS�TeA� �ݲ���l��e��*�Tm�R�M-��k-)�f��[E�ji��ڲf6ٳk,J�lص�6dY�f���5����V�F�Z��4��צ�kkA�Ӽ :��kRS]�Mt�V9�.��=+�
��w��OF���u/{��]oCj�ѩZ�N���[ڥ��R��A�N=d�hv�t��kT��+[�b�Ģ�� 7ԅ��A�|.{e=�л�r��-e=��`����Ԫ��������/l��m��>���"V��(U�N�=�=RD�ޣ��{�����0hUL��˺�Sa��β>  u�>�m){�N��c�}*�*�}�}���MJ�����Y-i"}�j���J��5��}��J�.����
}-�����ުT������_}�JUR>���|���7}�N��5VژgYխ�U5��  ��J��>�]�MvεU_yO^�ҚQ�x�R�Ї�N��R�s��t�m4�<��턩D7�l����Q�&�����eQ��2kmj[V��5���3V��  :���Rz�x��)6e�9�T�U�ӽҺ�*T;=m{Oz$��M��׽�J����{B��/k��T�+��c�x�T
����R���]�/KEm�ڑ+A!�j��|  ���Z��R\�s���![�7Wm*P���uݛ�J���t���Yoz�^ҕ��.��T�]�Q���+�N��q��/g��כƕ����;�Cmmk)��R��e�eZke��  >�`%+mV�Ki�U+�.x�C�^��Z[��=�!IO[�W��%�֖�����T�JW���t��e7Ta릁�����������u����f�jb�[��j��)�|  =���:t������5ЯAn˕�T�.�K�I�^��N��<ۂ���z�w� �^��Y��w� ���kQ[j	XV؈�Q� ���:�y��C��y��^=ֆ�]{���UQ�=J*��`ٸ1@�=��@�v����=]���R��	QKU�-��l�π��>�Z��΀=���z;�V�{������{�w���ޯ[ށ����\�P=�m��y����Hi��{g�٠�|        �*J� �     ��0�(���  C   )�1	J��"4�`�#&M4�LL"��M	*��      ��&Ъ�Q�L���� F��&�A5!#B�i!�������4����#�*����p�W��(�Rg�j���V�޾�^���Mֻ��u^����}{�TQ^x�;O�E�AO�
*+���" ������oH?7��o�����}��~~�^QTQY?�UU^��
��T��H
���f �A"��T�%P~БE�B�	Q�
?�%Q �E�!*��B���>(�� #�J� S���!|TG��Q�$���� @0!�!|	T_��U�$A|	UE��E���
A(�J���(/� �x���(#�H�/a*��J(�"�	��|	D��� �'�"*"x���"x�z	O@@�%D�J�#�J>x�/�@>��H>�x�!�/�#�(���H�)�B���C�$OQ<	SA����Ӥ�C �o����0ϴTC}-n^bk*�^�h�y�E-�W�YX"��,�ZXQf2��T��T/n��Jit]#r�^S��[�v��{�,��CmSX^i�g4M���9-0��9t�Xt���F!���rD�X�إ#6��>n�A�4v�@��bS�����(���b3*�"Z�j��m�	n��F�ke��8�����J&(�s`�$6u�x��$�4n�%3][Y�a5�R�L5�ݢ���<��լ:d�X��#M��dB�lm�,��f��7jT��Uf�B���`�5�N�x��9��k����,f_a4��Wv�[�أ�uĥ��6��d#�,����X��;e�5�,��$�.� j����li��(A�]���fe� �ȷVP��Չ������G(Y��f-@�\yW�{�d�Yӌm�U+kl1x��ЁM0��W���&���J�dM�ǖ�ǀk2c�ůt��rʡ��P.��l�YY����$��"AN��n�Bɫ�ڔ�c�1��m���n�:��0��PošWW7`6�6~ioĄ�tY���vq��+ʎ<Z*���J��M���%��s	@�DMJ҅��1�CM�+J84�$S�N�|�i�f�H�<w�WYu��\�)ˎ"چVk�N��K�'g#���ܛ���U+&C�V����N�\h��6�6��c0��t
#p��G6m�f4���n��#����ٸ�j�M��n��	��͘���c�S����ۥV��"���G%a�����le�T�3p:N�h4�׏Bx~CU�j��yO �i��z��#*����Ȇ�����dV��]tS��PWC���Į����{ H�2غxrP9��Bwm�^���\z�kN��F:�Rњl{z��I!V�$���0TF��<9Vdor-~�Ѻ�-��Y�	�l���wLzF��u����Pɓ�Ke=�,���*��J`�Q��,�:���*ab5ᖓ4�
�� ]�R�I��/�bl�@
��̶aNv�;v�9V�Or���(l9A汶7w�����!��3T�z��q4N��Y݉�����
�y)7�&�դU�y���i���x.�ۑ��j�7�9�6�9a�������Yp��e����&�*�3��OC���`�^ňJ
�n
1n��p�Q�=�)��%{�`��hdM���sP;���L��@:)��l�U��x�R1,bg�e ,����"T�ո�	��'�u�S�7E3��W�f���9����v�j�[%�v�Y�xum5��6詂#qn+��A��#��Y��.�Pٕ��l�ę�5��6�H�������E��U7@k�w�!�˳;4T���g[�{����͂��۳�U��P�f�	%jƙTŗQej	�w�+i�6^����Q
�_��Q�v��wqBC2I��-��"�Ew@�)E*Vn\�wB.��>'�FǉK�m۔,ܬj�xSܫU����iô�8j�o*�]т*a�ʅi^Lo)cP�j�?vR�a�B(*�5�)�>dj��fF�v�z��
ЉWsospV�� yZ, 2�`�u�f�J�0V���INl:K9�&�Ĳ�I���ᴵ;�������P�,�F�JdSWt���j�\(̕-�������N>+@��.�6��Ǆ�Qy�X]��Fۡ�-�8��6R;JT�n������cj��7[�qZ6���;�F�"p����r��֨��� *����"3�eX���@���/-f3Ln^�,�a*fb2��a�VFD�[��ٗ�J�gw��&f5[���3oEZ;4	�����Y� �mP�y�Jh����4]�?��Yǃ3T�U�4�dJux��ĞJ�)cUk>�e�8���M��:v;*6�2Ѥ��M`�N��_��ݜ��RA��.�"���\;WZ v�Vh�E�W�Cs(�oP����'x�+�JEVl)hL���4+/��嬃X��V����ٵ���M�Ob��)�i�ܦ�괺)�=X?n�A��G��{�9��m�5b�٢��R�m�É�t�����O����\�jv�+L�9�1�MHE����f�u�4唰!ZUH̛+S4�沁KT%�n�K�Zш7K7!���E^Z:�9h#hǢ��%n%����Ji��p�����$��ں)���Z�{�U�ݻ�]�c�4v�r�$���P�Ҥ5��CU���ax�86�pTT�(��A�b�{-d��Ԏ�H�.�$�`���.)P�ы1�����Y��^=,љG
e��
��X����T�;��4/4��N�2@&]����-�3q<M�k�H-<2SD�FP��ĔR�N������T��X��^=ԁ�1�w)�B�ݱP^�RAi�/M �2�>h�.E��zm%5\pȑ��c�a�P$237EܬY!�ӊ�tK�cX�Ie�p8��h7�o�1���G��K4e3�]��w�E]��C	F�+�V��CvLr�K�So���eKY )�����������&7eL[i��h�`¥�S��XM�cu+-�Y������ۥ�N�ڸ��`�u����n���:�z�Qŗ���o('�C0�a<Х�2�v���l� �2���Uf���=a��űG��3S�"YcJ�F`�7+m'0c�I����Uw#��Z��"�M̱M�Ϥ��f�٣��w)ś���j��2<��+pV�{������*hX%�V�3���A
Qnێ��ᥔSU{����dG�	Ԉv��	�-U��R֑a�z2R���a	cTF�t^�r��t�(L]^=%G��+��*�UrK��ω�
�u���in��e7�휻0�rfm���MQ�.�W�F�1� B��Q�4���b�/U��Df��Z{kl�� %�E�aV��x�۟Z�`f��X�6�J� ��J�Ѵ���"��W�]9��
m�w
�+�xP�H��uYj�x1�L��`n�f3i}��L����>�(q�2=WZD<ɼ[���|q;x�&Usf`y[IQ�)��{�JL��'Y W��4��Z�F��)��ܳ3rJ3�GQL��hH*�Y������x/ ��XB��3�X���N6�/ִC�����-f�T��D�G�3r�m`oݖ�+z����=���I�'Tz�^ړ2�@�x-ՠ�ҚjkYe��8�̋!%(M�-��7m�z��+�Lat��D'7F뵪�#T��&e��^х�+&���T��:8��C,V*�[��I(�XR�[`h�e��OB��F������SCr='�GO�[�teK�t>̭��w��ܿ��ʎ��vX��se�՘��{�zY
�ZY4�~��R}��!���m�Kk�e�h��"�f�v!l+�"�����`+VI�+^n�4����i�)I�)4�Դ�m�^3�V�5
U�,�J')&-�VѬ���tM�@3U=����fL�vP;Uv(ɵycn+t:��&\Ӯ�pJt��G(Xz�eX��@)��q�6�ɱ��܉�RP�6��[�r�X�z�I�tRWA���-����4N2�u�n9pIf�܍T�X��lc3�Eu�@;ͬ����'���B�ɑd�VmI���ё�Ұ�nQ��%�.LaӸ�ȩ����a�*5P�yG*JY�FŌ�%nV��P3�Y�Q Awim��fяcgfa������mRy ���LcJ���b����an:��dVk�Mr泆�	���M��%���V�؀�7E�5�(�xct�Eڢ�f[ڸ�,���Ȉe��+SQ��̬���ʵ��|���.�%��傛�֥�V��g��1�7hCU��m˴���+�J$&�.�\"Pv]J���"��U����e��3N�K"����̦����Al��Ux��Q��/2S� ��'䖅dH�����5y�Ò������6�	܅̦
 ̳[gA�ˍ5OP�dPblَ���f�Z� ���f��B5�uT8�l���k-b2����C���`���+%�24�[)5��wf�`r�&�	{b����ĝ
Ô���#��j�tSy��v:t`R��g�2�����c�<oh�9�!eU�I�9R�z�����(-[2U貶��I��r���67���q�iX��eS��D����1n<�ە05$�ޘm@�8(	Gr�Cv��e=CM��Mn*�|=�u ���`��n�����<��pS�cK$#KʏF<Z�,tpgh��g��������v~�&\x�q�NCY��{�����v6Ũ ���ì�ێ���Y05GUբn��e�F�Z)᫼�.?���c�	��)�[�S52\�66ؗ���@�W�q�&K�=�0���JԞ�����m�i���cy�1^�Q��+/uiBj1E;���u�޿�v;���o���mL-݈��5��/�c%bjU�AkT�6&��p��&4(w"4�T��^�I�GiJ�$��I�ǃ+*�ƀ���
��(�wtB��T!&���(R51�e���Է�Q�QZ+uӚ[�5ةs�w�^��pl �h�$�+[�#��I�L"�˛+Uں��
��2v�z�L�`�T�.�+�踨
f�0sq�hn�KV�U+0�!ۤ�cŕqd��aةUm�n��iLձ�j�����mYNrT�Vi�L�T!Z�]���]��V�V��ck��MZ�;�񯀕d�.μ�[�s0�yv���;D��j��1-#g�R����n�r�,t��	B��3eeJǁ�Y$IM�ւ",�����M���ੴ��q�.�#�Mj��(5PeJ�Y�U`��da6���jadQC�ZLӷ�@g��Z�����j�+/m`�s��	[HF@;����{��=����&�9x�:��LX=q�s\k+a��8误&Q��a�ܵR�;�>ku9���H��`��M���q�մ������ɕ�.H�(u<N�xLpo��^lwZv
{��.$�&��Vۣ4L1;��Wdk �&������[�*f��C�I��Cw�p�q�m3�?�B"%%ti�mV&���v�I�7��i�ׄf��[Cm��u)Z��������M�̦��'Α{�2�HX��W"����ż^�;��zV�W�l�#7�H���غ�L�:v���KS�V
�
X_p���egR]���J��
���R�4��n&��͚Ǘ)%6F#)]�P�
��P`�&8`��͉P�;��A&"�
�u��o4�IeID�k-bCn=��U��E���i�eL�X�SM̻�݃�p]�X+h�6ޕ��Te5�F���0bkf��|n��)��7��j��-���6�h�u�����"�t˸�"��Q=ˠ�j�u�N杢Nx��jx����Z�XUK`w�@?��(�Z���0�^Yg69y"��M��ѷ��z�,KJi�4+���۹yD�!);�[�ւF�!&Em`sS�2��2��)Aɀ5�e�LH��7,�kKv���ݥHwj�ե���w�0���gq]^cf����C
�:j��i���Q[����	��K)�Ǫj;i�*<Vj�E�q=�6��Z�ݑ�Cod.��]0Dٻb�����y�]%D4�bJ�jc�C:Y �`�Zst�ݺcp�tې0�JM�!=�Ӛ����
#5Զ(��P��3i:˙��50н�q�YJ�r�f1�Cn��F�l�+E���o*���NP��n�����LT�ˣ� �6=j�K4S�A�x��W�mS���(%����,���Cq�ܕz���4�H�����Y�l�CCMß5"���*&�w1�Ű!%�]en�c&;�(dsM��B���)+
�T���W�М���f�Q�Z��D�El
PZ�&LU�B1m-HZ2нA��@�m�xjJ��P\�i�ڕ��i�������Z�[��+P�L����+��|h2QȠIP���KW"B�ٵjC0�ۦ�ŋVix�K`+Q&�X)l@LԴ!�Q���Sr���yn�L�4�Iza��v�� ԫƱ��{BLF������U�a��eD�h��*��;��#��[օM�`Im�O�Qn�����<�@�)�=�\4�^�?-�f$�Ia�[�lSoɶ�L�j�n��F�l*��t4�,3F�0lZ:rf�,�:��4��ĭ�ύ��J�"n��"�U�0�(P�Z����˔��{@�a��:C^�[\����R ���*\\�%V5E����^���r'���9�ӊ���fB�__�f��+�ѹ��ٗl6)�ô�Ͱ��-�V���]���m��J�-�bz�K
���G�yx��Ci�P(��a�NJѻ��.�͌ ���e��IH&�K*R�6�:4&.*1wp!^�>��Ԙ��8uʕ��=� ���J5�3�W��(<��J�l,8E�O[o�hD*0e���5b�Z�%f���⚅Q�ZɺQ3�b�u� P�fRV4<�#Y٫W�&���n��CX�3�
�L0�ڹ�%�Pe���T�H��J�*;t�Q�
w	�j����'	�X�nFv!i�h�m�{�wVl����6kl��g`��]喑��C�)���JO �Mևur��vV$n�䒖M=���A��nd"��V&푺h�S�!����tͳq�A�9�f����nc1M�n���6Ƽt2�U�P��Hԓ։ܡ��^k-1H�Mf��(��Ɯ��t�Lm*z4iv=�B( �"�"Ĝ��  �B�  ��X�6�z�l�u�;�0g	,`�2��m�Dh�3�@��{��� h뀀��)��P�'4y�m��X���6X���]�-C�J J���0����sC���	��v_Y~Y�H���f�Ā9_�����������f.��U�����rh4�E�r��/疺��U�i��6�eh�-���� ?P�&�����R�L�nTU�����5T�7�@
��tG��X�;��]O�DL�r��:�;7OLs���C}\R/E[(�=[*v��ҡ��������%P��.��̰�W`�b����(���]W�0�/^u3Q}ٻWݨo��Վ���(��1-i�$,܋�]��ѣ��W:���`�L�Ei�4���� ��7�|�s4bʻrK(_#k���H��8l��u.�-;�{S��⾵�se�1�ʹ���"�� |^ N�}N�9m����[k]�J�	VF7�j2Aü�SN4i֪�����Wqui���y�����L��a�jb���*VKgo^�ou��C;R]eh���	�"=�\�|�ܔ!Θ���}��[�ݠr>���7X}��5��'F��=Ƨ���ˠ�Vwz`�l�:��;O.���+��Ň��UnkۺO5N�Ss��0��]���[�!����g 5�R����4'�`�E��g`�:�_	}NJTE���#3�j�ݑh!�r�%
�ttKS�+/C)�č��/+���P��wS�}�dRY���:����;���X�c6�^�=B����:��s+r�J��v��]�M
��:u_[Քtn,i�l4&nF4_^�e�1���W��?2L�ԪRX�[�*���B��Y�:p�ۭj��M�tu�qe�e�Ę�C&�c���&�>҅O9�m:�x��̘��w{���֯$���ܖ1�=۴�)$i(˼	fD�0��]k|�M�T�ۃ�P�U7�!��?9�E���X�H����M�֨���)��7"b�`�3�y�vge�U�՟v��txǹZҦ\���d/hs�	��۫�p�Jֶ�l�GLGJ
�^�9
]�6�n"{4k�V&��O�����E��w���!x!D�gV�*벓�R��j�TG�O(<���5o�]���m9.�v����M9r��RX�xV�{��T�
X�ZY����q��c���y����Taq��S;�P�2�3ܳh�ʓǷ>%YCaٗ;�s;`)qC�v��Ñؙo�:��L֙im���m�t�FK{"޽4��p鱮�ݷnvP��}�Ѭ�zۉ�O����#l��ZFdk`�J����.�TX�N�����������c������MY�+X�>�z��'�g���x�p&�����UL�bX� m'WY}W�*S�h��\�Q���1Z}v=@���sݮa�e�䄾x���`��(�Vj}��b=�nS�R��HU�Ȼ�2��HN�+��S<���2vTܸ�e��6%�Ƌˮ�Z.�mE����E��\�np�(�M����(1�Ԡ*i u�vҕ��G|N5iFs�:������W��4�V�vL�f�[+{^��Xx�Y=v��&���q�d�{���՘�ҍ*�7���)�o��,5���o�|������\<�� \�p��X���֧`U�e�.]��*G�޹x���j)%kX��L?r9���ޤ�ܾ��b��fۭ�f��ä� X������c5!�sp=��ҡW�����Z���I\q�����@O;85@��u�oM��4�*�gv�i'��3�x�%@E{>�"��ۧ��u�)�qR*�M���-=�6T�V�zռ��F�b�n�icq�MoM��e"���9�6�F���.�w�CijBχs#�+Z�Ŷ�א�9g�ڦaׇ�X/��vS��!ڣ2�n�Yl�՚ְ�+�O��KD���&�y
�"b���/�*`��hbPiJF��e{���{��^�jN8��Ie=���nY�Wn�81�691��]��:�p�����80负��崎dFWl�
ESUh���5�+���Ӳ��ޚ2Z��DRVe��9Vm��:���k�0~���\7��J%趜�w=�J�� ��[�YGv�t:��,�E�����OV�e{���c�J���K��0^�4��R<�E�S�k��v����[Ӭ����)1�;+�uHz��k��b��(���s�r�:�j��&���fsV�G�ȇ��.�[1���}�����Y1��+͗�Kއ5򪊄�I�bt�'t2���2�풏'�qQ,H� ̋F�I�o
=�)04\��	ְ{3@/,50�v��M|8�]8Sݝ��h@*�X����yϖe�\7���U���fNR��^�������fR;N�ɴ���}�'}ƶ�$� �'t�U�O),�@�CQ���G�+�-�E�E�˒T��Z�������}u�vmجm�����E_u��1@sW&	xk��]K.�gE}���TP�.ZP)[�oR�ŋ�3�Z�(��n��ݚ����{�/54�Y��q�X�%]�`��Jl�*�N���1��l)�Y�ËV���nq�qY]�����ܜ��.>(Ӯ�*�E<ܶ�n�R���Ŕ��{�����6�j�K7��4�b��1�`�Τ6d��S��ö���H_Z]��P��2�[����>��Y���,m&�ͭ9�u�������L��6�Q$N��oi�ζ�����B�U���2�D�7%f�N̈c�r���ga�F�g�+J�P̰&k�h"R��Ѭ�_NqD�u�@��ֽ����<|��I����J��poEmv�vl[�+�{��H,�`�dxnf�����櫔�!���V�Jz��:�r�&��4A�4f)\�3J����Z ��{G�;_u��*Ոv�2	g�(I�����gPǉ� ���@T�὆�P�OSƺ�����ԃ{�I��Oi"��rh�ېѦ2���m�#V��o�KhL�}�bXop�,2m[���֧
w��^Ef��kz�������{����*�3dWS:���������u���Ѩss��o��}�te�k�6�xy+���}o�.ڎsZ��(��n
Ռnn�Yb]n�)�Rk$8:|�|�\j�5%���f�k��]9���u��9>[�v��a�k-�Z�޾ɵu��P��NQ�)1�:�ͨ�o@�]X�E��+")љ��wK�2Ԙ�J䓳��j�2�������nX��}����Y�İ��W4 ��u�����!�w���$�|y.*��Y�vŢW��!b�鱾U ����{Ho��� ��Դ�V4��X:R�ϴ�B�i���-:�[��S|�׻�U�m�~1�4�fo��If|�9XH�7;U�{��-�ǅ��]X ��.��ټ�'D��LU�A��ԕѠ��Ҙ/��t嘨�֖��j�u�A�[ٙC�@)%��4YU�\N�t|ˬk	�P�Z�s�R��A3�j�/N��u���_k�u�.���s���ٵ�b����=.�9�ؕ�1sܶ]+��S�*cj�Ժ�z&֤�hc�6���]�3b���>��7�V�Ō�5�B\���x�7�nL��\!���˽����ꭡtb$�xB���%�{ʶ�bT�MW�<��U�sp�و�jZ�+7����MЏ-�a�R�'<(�k���j��N�s$n��LuL�ہ�jv;�y.}]%�Ojq��V�|���m���X"ۘ�SѫK�*���޺{.�S�S(F�[�0Y�dt�΅y�MCG]W��i"^u� ��l��|v��v�kV6���O���^}���L-\��L[��5�qvQ��۾*�WN�����s8��]������t�p�;���/�����eGW�K]��ڗ,}���B��Ө4�l�;k2����0��.�V�P$������g�C:˴�,��Z!��R����´7s
Y��D ھjƹ����Z�LN�a�+�}��9�<x�uNq@m�ݵN]����I
�,<"E�2V	��w�����6��J#
_g�`�o:f��yn�}�����v�C)��;��WT�!:��3}���WGxP���ڜ��L���`�B�ۛ*5�#.�TJ�����%�ڭ�[j�Y2�:��C{�Q���i��I�Z�GU�T�v n����k��2���e@�-�_ue�\����w(k����v3ScE��Ɛ���X��W�㢋��e��D����*�5l�(Pu��	����"ܥS���J�Z�S�.;���z����S��V,�f�_Ϩ��X��rMf���W��ݫ7��A�N�x���vΊoV:�"��g;�7*���$<��Dq�u5��������i��f�G�a�r��_����o��Ysq(�	]D����ڷ;\x�Be9��i�Yg���2��)'�cb�>�B�dANܻ���{.����P>u�kR/�����o)u0�^A�	[7i�۲��
 ��f���Y�kk]���0tg�(��@���)pu�}B��;7���O���\�j���*�$���ޔ�%�%��Ƃ�*�Ҁ_�ܫ�m�)�X�xY��-P�A�]nL����oGj>��̭���Zm��̜Y-Ζ�\HN�Έ�vPli�#�ou2F	`���i3�K��« �ɖ;�y&�sD�nқ�`Q����Z䌗�^�3/yZ�[P ��R��t/n'��4�7ƛ`Ŋv*^@9�2�:�s�(�� ]�%L�lt��Z�6x���Yq��@Y����)᳽&[YL�b�]�3,R�"P4�N� fs@V�����4��ΫkNv����n���v<�!�����{qw(sp+��.��r�q�T�ԱK�ql��Y��/���.q�"V&���u�a�Q67\m���4@7�Aݻ�،�qY�o��`����tp;hv��Y�M�
�`��ڥ]�1k�μ��$5�f���Q����i� X�y��8��F��5K�L�#�)�omXȺø(Ы��U�:h��H�Q���|���v�Vu�hGf�^iΉ�i}v$��b��Z'M:s{%��@��}���k6��6��&$�V��TyΐYF½���Ւ⼼J�0��9#ћR��-c=�O�j��=*`a��k���zX�'�(u�ބ�Y�j,�p-��v
-����atڽԘk�fmێP�k�����$���e�lc�y�F�X�	�Zƌ�,�ۑ���2��Eu��L�m�J=�]#ݎom0�M��N�I��͠�@��G
yA�*���5V:���a�xH` Y��&�ׂ��-\+���4η�
@>�K2�	��D'r���N��F�Qi6:벂�yV],�#����Z�����s��&�+
)m�7�ڧ]5�&NN�}�����9`,�'3.�-�Ht��-K��`�Y�Vu=Iݮ|e�{��WT���V*�Џ��3|6�,镧��H@���'�`Qx�ʺ�t�&��}�B݌Sfmj ����`!z��z�p�@YX�{-b��[�c�0�!����.�g>�4J�����X'�=8�J���͉9��ل<ɵ���\�bF*��b	A�.���5wWY̹#{��3v���7��m=wz�X���*���k�뵋�%gb%��{ݮ��wrī}z�����`WM�l���]�%�R��̀1���A���3@,���RC���Bխ)RtI_X��L�s������ž��+�d
���%e���ۿ�!J31Ae�a	��3q���1c_Yr�me��Y ��m�u�E��nJz:e��o[�-4�R�0a81W¬)c��g�S�^�ħ7��M��0���_ikV��%�$�>�u)�KS��V\1l.�kPm��j�5F�fx�ԳkUNܩ���WY�O�;�:�AB�,kV�
��z��3��m�Ԋ��onpٺq�5�o�ogM�9شt�k�R5��i��9k��te�2C8�эu��NK˵n^�7�ܹ��-vR��kI�����T�-o���
�iN����/)�F�	D`-uȦ�ޤ�n��(&����K��ɹж�o³&�`��-FE���#5X�)��Υ��6��`q���t�&x,��:X�v�5�]AR�a�� �ɧ!���*�;M�J�K*NᝃV<�0�<��jq�x�+�w�D������S��;�0K��Jadz���M�+&f\��?��\�(ȄM��;Q��l�E�.�9�<�[3Gw��tݮ�ޡOC��m0(V">�]44��IQou�d�ږ��tm\m�c=ur�M�2F�oz�ً%j�7:n��,�/�rl�ڃ�Ů���r�obe�v�K;n�9���h��ȓ)�)���r�+\Ȑ�����(�+S٤���;��"�X���J���6%tz�XU +�<չb�)��p*�ݒ���!�R�E���rY���޳��O�L!�=���ml��ȡ��˝@���ٳqoR%.��Y%cW�[QV�L�-d�h���U��0���
�թ��� v�j�/`s�:�:�wv^��+7~�Ō��"��齗�;�\���Ҡ�=���)^�U���{[�Ojfk�!�&�bnr�[˩�Wd��yk��/�����9�א�`uh��}�Z���s/�e��Y��Q��a��X-^��nN�d�¨".����2/i[��(�6R�a֎��j��8�i�]�(\�-�x!�]���� ����������#�c��IX:t1˾��IW����f�n+���a�$r�I$�	$�Zt��r��r�I$�#�$�$�H$�$r����.�������zG$��j�J^f릜Pu(~]Z�l�9�I�d���%I$�I$�I$�I$�I$�I$�H�RI!CQ#���Hۦ�nI$�I$�I$�I$�I$�I$�I$�I$�I$�I3330��ǋ�X a	$bHX�<$�RT�" �%�$pk+��5QZ080��4`*��*�U(Ю��_n!j�ha"���>$�
2'�"��"D N��!o��q����*����㈨���p�����S����(�� >�����������#�3�/�~��?W��צ��p��:v�^F�CVX繸ۊSޫ��72%m푔V�F!��s����{9l��,0�:�z����k�5^'w$0*�z�S�)��c��������S\�#�l� 7լ	��C��9(�����5P��:1�N\쥘eE�F���PF>:�N���,	�t�y��U�r�k��^��7�����W�:�,�wj��Y�c{�yXWX��2eC�[�X���K�⮜
s�T��9Cep�ku<&q�S��Ɣ��jU��讔m�ogB�Y�d��9�j��.��u�֓�ݫ���Gm
6a��j�|+I�{���땊a������ހ�yA���j̧*Uh��䢖nѷ�����f��;#v�+����f�����cKILy�8�c��M'F?]�/w^D���c��ܚ�j,�����/��&���Ҝ�j�f:�ԕ"mc��,A�,� EY�O
J��:�ފ�I	����y]�Wu^��@�!��W0�P=�n�~C�r�2�^��37�˪8��h����ӷ�A���U��X�I��)S��ٺt�)�-��&s��d\3�⺾ȴR��X�r��}�C-�V��Q�mʾ:��5��b���X���-]D��}g��N� ����CE<�r���N����?bF��h��4R1����丫���L�ZQз�̗��Z�TL�t�����A�=�(���(��Vk$覭�*<�p���IfyK���N����\��94�m�Kw2���5,G(͉��:�3��\��Z�Ǳ�/���ᕑ5(��)���]aB7�r���S�ɮR���PXκ�nڃ�+c���-�̕��o��-��1%Pۙ]a,��5qv�. "�*�P�)Dz��Y[�/��7DE�V��%&����4p����x`܂C�.�grgP��lPu���}tM���u�$C�O���̻O+t�n�]dC���<8�b����!2��m�J�@��,Nnq��F:YX�Up�3��6�L�&���M�)�H��g�v�d�%h�����7�+�et�%������wb�w8�mv3\�ɰ�mH�%K�j�kYʞ��Y��;��,�d�n2�l�ϵ򍝾�<����[1e-c�wS��VoZ����*P1b�g-З��g
%ޒɘ視�I�[ac����h����6�*M9AÎ�-�7Jtw�&�݇�����(��l�tёd�1RɂL���ڧ�T*�tҪǦ"�^�COR{/���l\	���hp�Δ�Z��3�*�M|�|��e���]7j%@"=��:aY&e�k�0�u\:�\��Θ�$wfb��(�TP;Y:`p�V�wG���:S���x��tv��1�N���8�Rʎg�����N뻴�:�㮯�ȑ)ήYGu�/;jmY&�ְ4i)�n��:�j"�+ �ꑤ�b7��k��"����tH�fC�Frue*ƅt<���sWA��-��oce�{���]��@)��Yw���ǜ��Uݮ8	�nna]v���GC�.�q�s2Q.�����9,Z�9ep��G'l��9y������\�*�H���;��;.y��ﶙШ�'�)����9����{��ڶ\�X�;�UID���s���\9:X����CY VT7bk�q��FJ%Er�j�Rx�̫ۏ"���/(���[AZZ�ʛ̓��	���r��#(U�gI�b����E�53�nh�7m-T�̓>oP�T(%��7cMer�&�S����r��ƶ�]��h6���S0+���l�,���vj�C3r��#.�V`iH;�iU��.�%�MOȋ
�:שS�[��],gr ����N:�Vu��OfL��Se^�����ki_춓;��:X�]�掦���p�Qحi�B���㹉Ҙ,1�m��l⧯��T)�#Ρ��*�8���d�Ss��}Te�樂�k\�&s��4'1,���_g�s�������ZԺ�ȞB�VT5���%����xwr�J�z4�+��Vuꖕ����C�C[�o�u,{o���,	K5�4�ۇ�=+���r���{U&��L÷]���t�],[0Z�svn�<�^��U���ʋ4d�wS�R�^�wh�R.+[�/)OQ�\D��[�tܤ_
t#�NД��u��l�ְwq��J��6��)p|w0vM0����l¬�+17V�ZN��ʺgQ��N��[w�lK�RNJt��0��`���q����l���K/���]���-�C:�d�]�4+�x-�uWb�Y�t�EΫ�����B�e��δƺ�f(;I��2j�8��Q�����ݺ�t�Z�'����r�h�H���VW1��8���9�\-�dέ��¢��.J0vl}�pu����Ҡ(飐f�@���׸��:��&�I�Ni"�A6X�[�J��I})�*;���Gam���W,IlW��i��I_.o*p�y�����+��AZW:a���뙥^!�& ���R	f��9mK��J�sg�����5�Kk����-8�|�m�c��kt)�qJ�XM�7A���3+n�:�shŻ'U�#
�.f�vRń�]t��y�M-�&�9���Z�]�K�o{qdpMD�B��� 'G&'���U�k���/��u+sLoiӍf�xu����"����ú����=˴�n�k�-[��έ�D-i���zV���v8�yA=��wjR�6�F�#GS��ي�-�V��>YI����� ��N��5=����*賷���3��l���)���OErlT6���vi�dH��.��B�:�����3AW�m䃻�������*�˻I��Ҹ8��ZQc7��6��­�2q�[65vuғ�gʦ���>���>[��,�,�C������N��6����e��e�(0�)���g)�޳N婶��o+ݾnۭ=�!��/�4F�}��E��K�^YQ����u;X�j&y����7/�uӖ�yu-�6�O���[�����v�1YY��K[-�(M\q�SMy
{\Z�������pͧ�0�ʝ[����c�ZCQ��r�{+"��2��d[
�6-��3�)�m 3--��YA&�m(3uK�ա��`��u����5����vs*��/�횗���-G��q���y�o�(ֽȺ��,A[ꭸ�a˲�g�3s�<*$]^;ک�\�t͉nke��+4qFk鶺e"::�vi��F���XOgWkΥZ{6��T�ˮ�k�㕏�H謙�U��f\DN�k��S�En��{��	�g%��f��.Vs3��|��:4�]V�(qr�����`}e�"#�c��WW|�9���ّ���e�EV�@5LCpwU��Μiˊ��rh��RL"8�վ�[Y%�6.�pF
�Xh�)������M^��qE�o�):��#��i+YWφ��nk9Mu�E�Y\�b��u�.g��;�ۋT���6�)�E8	��"��v�4�y�Bǝ��Z�qLjy�Z�r�7{11���̫��(�ݾM�ZS��W��՘R��6��ʂ`�%[��]�Y�gD�e���X��*���B�M��v��[�oE�w����Xy|��<��|{D��G҅�B�����U�EXԾ�r
�k]N�:w�U
�mgjN�ۙ���K��M��3�����%C�KAR'T����k����>�me�RuZ�S9�u�,�{-�T�u�G3\�g��k��d��]�iL�|޺�rn�.>��z��!۱9@ҋt������^;!5|j@8��W�457r����f��51���V��+"mi�K^,W�ek�;viOy�Av(�:�۱n�p��X�,>�����2��ݲ�R"`��w�k�F�䫥�fܚ!t� Sb�6�(�ch[��aHN��p�����.�teֈ-
r��(�-��
d����M�N�V](�m�1Mgϲ<:SJ��V�b����n����Πw�LY��2��Hݡ+�Ӻ`g]b�v�cR<��Ό���r9��Fe	Sz ��Y�<��7\M�"T�UxRVv�}��2�m2M��B�w�r�mf��s��jq���f+�m���J+�E��i�����Ñ(V�k�v�}`.&'���e���9k���i�ו|�5A^(�&����5�c��R���6��)�!d��r���E�W@��z ����T�z�q�T��*�];K���Ίخ�}{��B�BTK>�{�k�-�}N��Ί;��U�%��K�e���8)bY�w��Z�2�*��V�����ׇz�I<ں.�ΔZ�^m���ke��8�j�.�Jr���U�=jӮ����\�1�1�x,��?0�e���HBJ�WJ�H�c���d�ܩ`�c���k6��5�-\;��R{�9��X�}�/i��>o�Fk�^$U���i:ͽO�lE�U�Ki�C�5�r���r�p��s�R-���0�Ql:R��s/k�
��WK������z���h9]����՛��P�|!ŕ���T)���V��D3B1���+�]�]�*��̜X�g*��]<���(�N��9��h`Tێ�1�tlS8�� ��9,.z���C{U�l4��
�@'�t0�ѡ�<0-ð�*Kxۨh�ԙt��Rzu�W��\ױ��Un[W<��u'�e�Nl��v�<)�t�o]���6%�re���n
*ފ t"���'>or��n���TGe:�CK㗗M��%�m�j�V���u�"1�s�,9�{ߛ�f�bb���ŵ��a�l�"�bkܮx�_�2�0l����T+J}4wF�B�q�8�X���Z^n���	$���X�����mv�� B.�5���C���`	F��<�j�@��^���ʌ�ܕ8�ͺ�otL<KNk�@�e�Se92v���e�YS��-V�ɻ�-�;8��Vŝ�m0B���̜�#`�Z}6!S������\����St4t�i�Lu+8h�]�2���K����F,[��3U��� �Y�Q����y��D�n���Q*á�g:h��"�)1f�v)x:��WedW�����ub��V�yu����y,�f�,X�:㚠S:U؂�ƞ�u�sRJ�j���`
�u�"�����i�-�z�3\XQ��\�����Q�\��T���u�,�Y7_W:O�KX�Rn7��� ��Qۡ`�u��	�9U�7z���5� r��Q��&�E�u��]-ּ��I�۠��r�ͭ&���f������ש���m5�d/z���Fc�ť\Ot0D�S���u�d��T�`[fW5��C�j��$���-�r����r�it{��[2��/���:�B;��[�h�\cU��� �ɱWI�-�\��m"Kߚ�����$�0j*����>�����\�t����A�s�8�g8�Q��m3-�rr%P�ڝg2��ai	s��+Z�V��g|�h�×X*�_c���h��Z��do7
��e��quC
�;�}3����0�[������.���ق�l��DЧM�(hйY�"�uݒ�ި��eC)L�t���㔆��{��bQ�W7��\x�ޣl���kU:��1��`�qt9K�p��_V�(X4��Z�Xo�wچu��s�.s��X�ߵ���"ݳR�<^��kM������������	�p]��V��C�5��%)��s6N8�w`�x�h�}t��ĳFfR'���h�ޤ���᧍�R��YϾ�+a��J���-�­�r���)�7RE��AU��xc�:�2�S8
�\ֈ4t�-���5QC1�R��B*��Mnf�50�wϨV���_��<nV\�̒��(�0�_p�'��j���֮U�!hn5'^,�AR��T�� T���o�+��)�U�2�;����_h��8�XJ̠h�Z6�C��@;9T�|���VZ��zs�ؽ/��"��X�w�oof��9��2eY:�j����mf;�a���P���r�[KS�n�����r�E��4�V)��N�fGm����F��T�rK0jQTV:�1kh�V+��M$l	��܊PK������Ņ��;㹂.��n���6�Z
���;�$�@7�q��]�p�h]���u���f�[c*��i��FXl��u^NԔ��X��\�A]�g0��n�Tg6ۀb����K�˺��!��m��u4(�_-�)�wEңHf�zi�H�b�ԝ6�ޠT�7%��wmBj���$Oi#_-�Ziԝ�z�pА�]��sN0'C�Ӡu0�Rf-��P� ���n9�u��8O�,P+	cPGN��m�ʭ�{1+²Gsq`(���Y 0�F�.�Ƥù)���g0ɼ�֩J�}Clj��ׯB�S��y}�A�k�!#�;`�;��v�8D�%�[[a9L�� b�R��1�;�P��{|j'7a��_V�9���h!����)ow�а�)oQ�c4s�k` �wY]��=�x��F�kh���Дմw���IB�B���V�*a���V*,�W���R�(Qy���!u���aީ�W�f���KJQ`�ch�%��w
�"F���*���{�>�,��U5ҵn�w)���Ѕ
H�P���swn���n[��9��nkK�1�F�3[Ce�����tý��p)�oz�F�{�!�n)1�.�y;bI��u�s�Cz6�aq�.D�;ArZ7�:쮶�[��(���u ��<��I8�������&�,�;;���o��Oct�9tú,+�#F+�У��ԙW��R�9n��E'(�N#+���V�ɛ1��#��P�.\��H��WW*X��k�ʣ�U�ê�@�3�2�:��6��9��]u����ᯒ*�+��__�~޿ԇ���}!��|���;��%�8=��|0�	��A����T>���C��6���47i��wu��L�Z  խ���1;���S�F���ӢS�Ǫ�8h�h�%΁�mf���/��e�ܙ�K��pŜ� :�mgW�u�鶯X��n&Q�����Q�,����"�}ق���R����F�^+�����k\oK�: ��[0LҶ�=,�{ݙ
��e��nܹ�Pu�j���[w��)���:�aQs�x�4�ͭo,Y��Goq_u;)i���=`U��If-�o��:3�{�Ь����T|_]��.��BE8���m�X�s�*�ͪ/ht1�pR��p�x�LӃ�XC>���lQ5}8I��J��e$95�m�V�F��d��,�����h���S�֥�0��y�&�p�d�2�`�cJB�5�A�vhUo(ax�Y�oD����;v!��r�r��`�\;U�I�U�Gu"�2l�^P����4���o	�VfZX�:
9�*#���Z�h����rM�+����n<�ޖ�\BUP�庶��"�-=s#}/�E�I��ڪh�Em��zn����a�!T��;Ya�#��Gk�n�Xz�v�"�K�&��g�I���wy �A\����XJ�h\�%�]�_ٖu����r�S�)8INHZ�$��!��T*��تBE�XP �)���E��%�2 )J�%% U��%��3xE��P� WS�8�7��nss�r9�%BPReYD�I��EnJ�hL��h2L.##��s�.M-	Z�(D�!u�UI��G2�#Z��J��7<N�B �d49R49)�r]Mn@��ܑ	��"���6��
�-J<C����(��'Pj ��C�CI�`eT@���,��G' 
L���7�44U	KՐ!�Q��CW0���C3�
���5֍��y��k��*��
��$��Npd��3�Og��Z"�)�.c��1������O�ߪ������$����v��[�*	Ί��1 �1���e�ii� T�S����^�_������)T�&�7<����rK~��]<{C=]�I4�4�x�����c��ʞ��k�"_�4����֦�@{�q��L���Ůo��.�v�X�w/���"��L+��u{�"���_ē�I��;NHfbO���S���Ў��m*r���=~:�V�0��U�.o^���鮯���]P.����������s�һ|�Z�T\��mK����������^o��7Y�/-뫜������+[|'�I�j�|�r�j��Ԟ~���>���1���M�a���H*<ul�<�ݯE�|s��%{�|P���7�~�)��}ouf�:s���~ƍ6������Y�����g�f#!�6�ۤ����A��ٍ�N�c.Ks��H]�F�t��Z0F��6fvz������sϵ8��S���;-��v�Sl��Z*�u�b��S_w�
a��}�Hv�$�f7t��i���Ky��s�0��/�v#��N&Ė�!�j�p�h�-�K�1=p��p�����F��oUI�I3;<�u��9��/>�鵔�Ԫ��������2��6�ޛjːp8o����w*N��O�0R_�f�x�����ʴѤZ>��r��Rj/A8{�+(���P��&�5qKӸ��P�7�����G�}�V��S��M���s|;��p�u�~��2�w�_��(���> a~�(�a�}D�o�?Xک��}SJ���ޝ~��?{�h).W���kHx�s댈���5�cLD�b��2<MOh���Z�	0(���t�:�7\��2X�j����w�H�O�o�=]�n�\f8�;��'n箉78z�ϲ��qF�^�k�OK~� ����U�! %<&���{'�W���i���<V~�v��o�=i����L^o�W�����͔�
��~FOt~"���q�ݽ�.�YF�T�<��;��q�Ӊ��M[�lW2Vuo�ʋE���MP{�5�8
���|��"�b%h��5����l�
���7�2����Iǒ���
մ.�r�.Ic�%9C���*�?[����58v�kZ㚵��u��ma�;"1�MvT��6a�����R�����Ow��/Ēj���Ѓo{1�.E�DNY��1���>�=��[V�I���}�˘�����ݴ<���������;�9ۉK��զ�ħ>m�<�����?C&mC�����mX�;L�%x���3��>�Ygiߨ-�
�ǃ��c��f�s�;~�{�������%�U�>ؽ=�;\׵��n��1�r�A�]<����a��_��L{��zt����g�����e[���lXeA8��؞ʊ��r�/I�zdWދ��V���jU�q��ӽ�٫��\n���ޫ6��ʞ��DX���N����{���>^e��=�֗�b��X���]	��3m���4�����[��PS���g]g,�}�.dn���]w����)�U���y}j5O=��wș�8!�[g�S{p0x�'�%5��g���˲���(��+�j�<��t/��,��W�'�#�3ͦht��D���
~��حW�p�~;k��mV�}�Ձch"�mi��o���wk{h
mK�z9�S)��w�����rؓTw\����w�7����V%A�9�w�Ɨ��I�~�b�\��'��u�NTY�w�����x=�o����9^�E�&=�K���q?W�R��>�X���dޡ� ��Ӿ]����c �UX�#}oOȂ<!�~��^`{������Ǔ�;�|FW~�:s+���[����w������w�I�\�y�y�}�~�%\��A/pڐM���BW��q{�x5�H��׫��Q��t�����2wb�O<���]Ըl�s:O�S�Oc��f��ľ]���M�[�0�|K��X��}�ׯ;�5��nz���U�y�{�V�E��+�`y�8�8�`��Mgz�JԜ�\�Ά9�;@��l?ldSf�5�����i������H����E����^�3ދ������z����>qU��==��'�u�W�W���+ْے�������p~Ju{��!V�ݖZΡ��?9��JS,Z��F��*��+�ȏ�ʿs����E��9d��p����L�b���M[��_Rd���uIF�k9���i����I1�st��=/V6�iO:��uź�a�ƼZ����MѠ�J��.@�w��5k��{[��ҍPK����C�/�3�L�(R罾�����ч/$BW2�xݹι�M�E�gE]�iў��2����v_=G׎\iDw�}�ew��k�	�Vn�QF��vL��/lM��՘�KS��+�����{s�I�G7[O>��kM��������n��=)ڷ/DjT��M'�2N���z��~F7(��䬟ILL�.0�7p���B�3��ǹ�{ܧ���yn������nz�����#i=���"�RkA��u����(i�6�2�F��z��ڳy�Õ��&-�*�n�4i�9{�\�y������9](v��:|;��hNC���y��l7���j�fï��Rc���};�T�9�o}�τ�;U���2��t�zg�u���=���U�C�C���3{�={Q�q#�C
���k�9���~>�7^�G:7#�b*�G�>���6h� >�k���[N�4��2]t}�;@�������um��[A��͸��bz�_ei�]JUw'�q�%��؜'�:k�yZjU����.,���)���r���j��7j�rh��*�ŭq�-���v�x{�7I�lg����.�rҺ�޽�זC��aw�H>Ξ�DX�"��ih��w�㦼_���ܑ�_v��.��G����{�Օ��T!�@c�3~��E�1 �?I;�,�p�/4(yM �Ճ����!w�=�}�+��<I��r����׊�K4��ӳc~f���.>;/=IjN���|�-�ʵ鵔��;짍s9yL�ʍ���s6H��y�ٻ�u\(�!~��Fo�^1&{�(�/;M�sc6,���i�z�����ǰH�.F@5������;�yR�k�����b]ܡ�"��^��:�@������rN����$�iI�pB�}��:*�����>���{�)$��W�K*�.eg���Y��?!��3ޗ��2������i���a3 Wa��ȳ���:����G^���w�O��[}�3K�2�Ӷ���գފϞJy�}�3��4���#*h&S�RRMq��'Z�PY۷�ިƜ�泼Uv��s:9.��f3����Υ���܊��a8a��jg]�\-B�HN���~��1�����ʌ����1/�U#�_K|����{lVz�I�;��d�Y�k����x���z�<Ƴ(GS\�9o�G]��Lw$�&�3�	����/o�jߧ�*�������T}����춧�y<#�W��a�Gs=���/k�u�+jBsj-'/�^�(Zi*;վէo�x����Y�f_�<8G�5�i=MǍ1�̲{���L��6��!��|��@�z����X~���%L���^UqN���~S�W�V\
��/^�ߵ��h�~[SN��Q�m��9���?s�U�́&E���	[^�1	�h����h�-�M���v<�O�0�F�/�r^���<x<\Ȼ�;�x���P���^�}y��<��j秭\@*2���x�u��ӟ:z�j/-�z�G���3�u_����E�^�l`.5���F@f(�Ic�-��j*���KE��#��;V�p��؈=�W�Cl�|!f�d�y*���o�77�+�,��t.��w��u���MY�%m�A��e5�J�Z8d�c��P���Īc�����w[����a�d=���mn�I�R��<�2��鮲D/�Y�r��K4��?^��m\{�>c!�t����l��w��}<�L0�^�Ѐ���]�ʕ:n��)��i�5u�M_z�m�zs���0u�_OP�E�v"}�%q��?���[	��9k/ۜ|�t��J��~���(,�r�}^�W��w1�[Y�q�\��֢_<�W��7|(N?+O��x�un_��ᾒ��a�2/*�:��0�:�Z&��FX%�n:8^�)�b鎚�=yU;��S��>�X��)�M��$5�b>��k^�@��S͖��3����M�q���y{OG���o��"#<���%r��O��E�X�F���X����6P�W�`H�g�5�zN��J�N�GK�l��\��k��}�_1�}�US�Z��$�2Y��^zT�2�7�Jc���Нgqܓ���s��<��+�F*l��X��궢��t}�_U�n��맼 cs��̘��=�1o\G<{�q\S��5����k�-��J��sR�j�;éڢ�'dQаA�M@���6N�o#=��t����Q��?FO-�O���8D��줍����i�sɃ�Ŝ��2���s�9����������h����$���{�c�_�yʠ׽8�'��[������S[]wsʋ�K�S�u�T�����}�I<j��T�>>.����>;n�
"kLnJ�N2]i>�1���˝�'������}<_��ϜҪ͟]��<��j/��6a�k�\��þa̪�I������{u�	�D�o=o���j�����+!oז��)s��T��jW}"�.߬rݲ�{%�ZM���z>ٛ�6�n�c�1��+�k[�%�vk�E���,$i���QI�����ƽ��~b�UA
�0g�����^���]�1��-��WO��}�Gw���y�GS��)��S�ї��|{�M��62�E�R`�=��?P�|-�u�<�/l31N�}������l�m%�	�b�W�k�Y�Z����~������N���葘KU:�w���+x��wv]˒�v��8�x<�Kl�)�G�x�V%#�6*�
7�h�L��ļ�͚� �4�l���M�w%���:e�D��q��2�n	�k+�V���JIE�9��cx�Ŏ��+�"�	R8�f�حo��hK�	�C�j��Z=7�/6M��"�� 䚽�*���Ï�m�n6�AU	�|�ݩ%��?]���5��8}\Ve�{|#�q�/+���v3d֎5QTgfC�1��R1�r�Z���7E1�]���j�y����Or߻о����ܫ�zіI���{�Ș�����˥=�����s�^yι�w��{�w��b�;�=&�����/!�Nw�Hg�ɵ��"~��fL���޶���/u�h{s3�$-n?Qo�공�eM����ۋ+��V\n����w��v,������VP��"�a3�r���_W/����e��{k1`I�7��� ��ڂ[��ISё�3A�׹^z�ҍͩ��/>�鵔�ӾW,���N�!z[���\��zE��;[�r�ڹ��0+�^�*�_h�_� �X   ><5����1ge�{t�V�_f�⢅�ų��r;}J�-�(6�B�h����&m��x��Jus��X��/�'�Q٥6��ܟpזލtw���W��عq8%����V�U����W�k#��L��{Q!�u����i��9�U�r����sol��+�	V�&!��K
Y9�m��o$-[�2���Rˡ�J���D	�2À��E��y�t�i
�l��ժ�qMӣ���C@L�$Q��;]&2vMH'����}�̋O�ڵr�9H�m'{#�Z,�1�e��¼����<�[!.xN�0m�"�YMr,�v��������
1dv"���(T�`>��GOV-�����+ɛ�lis:̫��S�S��,s,r���0|Qj���YN`C�n3R�������m�T쒤|ZU�vTɓ���;v�����V始:�Jg��ފp��lQ^��[:��3;N�i�E�,N�1;�i�zNf����};��/��MP�R۴���CEi�dX��Z�q|��}y�˛ҳ��� i]��'z��#� m9n�⧽C�8��"mh��7ۗ)�m\G��qI��VS�޻�h]�G{w��֔�b	�'#g��O�f��t�<(�¹�};gCfԵʷ2��Sޝk�.�4t��6��3`��&ʁf-�� `�;%N�U��x!sqݬ*�]s�(*��y>ğ.x^�0�c�^�c!�Q�{��V�R��gVY	գ��;E�:�B;�z$XյXأ+�B'X�!P
Og�_�0ʾ��Hm	��ݷ]�=5�n��ޥ�rH%}@Qu��n� tq�2����r7C��Ll�SJ���#��m
�)�e���~�'<�$�2��wW?fK���}�{0�A;�m#lY-H^o8�-�8bqY-u;�1�����e�)BqΦJ1C��t:��F�+��]�B����vY�R�PCAB�f��G67[e5�K;76�6�X8(i�&+G�KH�I4�VHم��j�f|���m���7PTB뚣i[ڻ8X8���;c��
��`����;&ne>��s�r����t,��p$[���
�a��*E$ӱ�"�����}'�|F�;,Ė�нV����3Uƭ�]\�X#��f(�dA����^v��bN�T{�j�
ĵ����:!]9q/sJv.I��ق�G��`=��g��h׆�b�VF��:��:��oAL\��y��[Ϻ�\��N[.��ac�W�ή���D�_p4780/2��ތ�2��v�N�����T��l�{�f��累����I��\��Ī"���Q�sH��%�0=�5ŨT9�.QC"X�_�a:��IW��f�)�"�q�a)�����^�2 ��S��;ȹ�A�&���ǎa����Sf]j{��y*q..�И�ͮs{ww�ې���,�1��D\��Nu�r#��)���s�ۦ�G�?��$|<B D"�$2ɐ{J%)��.��/sư")
 �9��p�	̉�8��K@j�J2�����5 d��%5	�nD�% q�- �'r#AZ����Ւ<@�Wpd�Q�Za8�;���r�(�N�a�HX`S��7!�A�uFI�P��2	x�ʨ�r8�%
hN-��;���b�B���2##S��X��vAN��&IB�C��$�Dk0���0����
�բ��9��^&����sX�g���߫���o��˾�>�4��	)�!����4�u�����SG9l|���B�Iͮ	�וW0��� |8����9��_��.'W��`k|\��1;�(B�MA�P(��7�����c�*K�ޱu���z����������Nd�T��b��fŝ�!���i۬��D����'��t���G[�UN����.��s�
�9����;~?a�=wU&�y��oGlv�"�pOFm�=�Ϋc�z����x'��ة'ԠKS�W�r�7��\{"q�bQ>�|���D�^MR�08\���5{]��_�3�YP�]�Ч^�
^�������˝�`�`j}ut	�v#8������ϝ�O*��*d�דGK�s%��֟y��Pg��dJ^>���c�K�U���=��T��7�h�g��s�������E'�P%�AS�d���u����/�������A�-�L�y���ߙOl�u�</��

Qqr ҳΓ�~�5P��Z�a�^''%Ȅ$C#�+wO����O��O�B�O�/'����L�>�䮚�p������^+]ј�����s�+�#f�x�"�ǠV��*;J�p������y�E�*��eH8޹����P��6"=����k�M�=ydV1��b>
���mAQ��F!�3���^���0h�
yL�S%ۅ�5���ͮ�G�ׄ��h�Q�R�s��,WIgk���C6�*�];P!���x_N�a���]���z�$��L-�)�<z�Z���������?y��'�g�� κB`bJ
�0�\�m}*3J�Y����:E���E�P+U�u���;���ܜ:��lV���B��q�P[��⿥KZ}������ך߷��ė@F�P�$�a�����?zk6+����k0DY0\aB�\-���'ى?uw0!Y5}�uO��]�]`�E8�FE����b�*�ނQaߎ��}ǟ��.u��ŷ���5�N�em��������[�um]z�۽<�j�q�hB�&9>�S��}Ux��碐�+�)I��(�Y�X��pM�`^:�^Ť��Q���8w����Qk��L���?Q�`�u��KL9�I���I�;�2���18���8�5ϙ�tR�g��f�R�͛ޤWlR]y�?B��_H�8�Y*���[s�8���͊�cu�;��=_A�=�A�G)ƗNC���xi��sb#���YӒ��I��e�힖S���6�E����e�c�Ǟ�f(��r'ψ��_d�&�B�-7��wg���v��`|Ӯ
�x��7s��c۷���g�Vv�7����J�㏀���<�a��dv8m䓧�R�V���-u��v�}z�D�!=��S0ػ�}�R��m�xeC1V�C�jǰ`��gfT�����N2P��W�(V�b?  ��l\ґ[u�������
Y�����'�ʝn��SE���e�V����yu�ڐ�1��A֝.�Y��(�{[��8Џu?C��BWqBG����Ũp֦�,����O�"��0�k��|N��D�k�,�ÙAZ��:���l��T><ː˲�ɐ�>�R��4�q�B�c��,�S�^�s�����*�l̍�&o�9���#a�.z�7r��O)��M�+ٮ@��u����*\��,(jS�T�GD�u�c��|�WJŮ2h`�����?^�~�c2Q�o������|`Q�㖫�ZFKwX[8D�}�3CEG�']�u]7�^�Ɖ�����t��-i�O��G�|l]��K�[�	���q�
�.)s\�?l��EV)�%����°��Uҡ���y���^Y_���z�+lny)1qi��*��N��͛��vɊ��d�\x��j �G6q4��G�����_3��� Η!�oW�Yy�ڢ�6:3�5#��M|��Q� ��a�l����y2/�x�����q&D*�&�y�u�v��Q�.�M�㪓�1nQ�uj�i��r
e�����w\R����L�k;U��I���l�}�r���7��ӈ��Q0�<.��yRq�F��ʧ���c}1�ޝ�Ț�x��܋+c+�F��O��_}U���a���;5�&Rͬ��`.g�/�V��twUq90R�蒚�8��ȉ���ₒ�Q���_j�G!��ì/t�!�]�B��#y,Z�lv�7��=�`�u��/�C K��������BzF��7�iC�z=��^�_�cYP�ꦖ��La�(A��	u�Ր����;��ȉ�g�FE*�Ž�I�y<K�:�|uOr㚪"[�ѩ]��r�)@,��]
ǈ�A��!Pa���u�� �áj{��D���>�ٮ`�_���<��m�Sm��,��s��$I��+��W���q�U�B�Zʈy���C�xcHw�X�%�v̀C`���
��]7L_��A۪�Ȏ���쓌�۸<�S"����Y��(���y���i�vʘ	�:���	\����2���Q�D��1)�T��ª�mA����&r�\[L�E���qKM�:�����k���M���܍2/jB�<�u eAN]E�j�n��c�Bpa�iiw�֤���ќ^P�@3ǌ�"1��ҡ���D��R��%�EUr{Q�9�R;_�d2���i�*�������6]8�mҴ�CYfY1iY��a���[��}F�U�fGOh�kn�V�����v��9&����Fd�ɘ0Ԣ�2�C8�z���)'��Oe�%�:-@v�k��m�K��̾������Y��$e,�ۿ������7�[��K(g������'�ڕo�B�9`T�sv��m�R��@�0О�'bl�w��v�c��E���Y�E��j̐��f��8�ԩ,Ȇ�q�t�o�E��ˉ����*����і��c��cW��9[;" 3f�S�qڠ�W��ʮ�χae�m�z�K���cv��{���r6*v+��v����"֤K����q����L��k��U��u`)8�{*PʄH&F5�.�1]����A��J�T
">�F2g4R��G]L_�����E�2'��B���u���͹G+T7[�E�ޟr
��>V�f}p9D����k�گ{n�r��JL�Pn~+��C�t����c�2}��̻��7��u(6�����c�FGz����	7=Ѽ�w�V�n�躕���b���]Y(Z0#ќ�W�T�|F0���V������nb��0�yV�Qöp��{�x��e�a+b�"G=;�z�>cϜ�Q�)�_�H�U���}U�:^G[��e]p�j;]��&��,[/���m�
�ֻ�a��w �D�^*i�d8�S���]b浪s�q��C+t���ς�x��-��v*d{f�fwD��Z�Sy��u���Ym��z�_�7���~�_dW�.ʖ�Vz�oV�]�4xI�8w�QWbi�#���ZSM]��)�Ԑ��t��Qe����Þ�[��5ǹC�*)B!J
k���m;�O�@M7�#�:$����}Jy=��E�ޛ��oM�*�¥ύ��1��N�`p����8�����JL��{(��|c�s�\���J-99�T/�ܮ����?-��¿)|�����\*�k������Hő�J�I�n�	���E��TY��TEݾ���E����9QY�{�����,�������9P��q}D�^�W�P�
[8�M����6^�n�,����ģnS?��WLY�����	��()�̮r6���.Y^D��-M�.�����l����(K l�z.SI{H�e�O�Љw��-&|�0�њ��yBy舎���*!�u]�^��Q*SYН�>��O��Q��u�F�t�Y����y��ؿ�j�󝢸�L�҃���Z�'6�x��N741��F��	U\���:x�;������wt�P��@j��H��)�Ky�Ý����.cvGW���z�%���=�վJ���9Ss��ٽ����P���$�� �u	���BB�pM�`^:�Ff�Kc\��'1FyK�!�oJ��-W��S4G|�%�(�l9���ӷ����Ri��ݭ��A��%�y����KQ��0���ʔq�0{f�h>߮1*�s)e��*c� ���SKs��/���Qt�X"��(��7-΂&����*S���}U�UW����=�C=ږ�#�ܯ]�a��|;=:k�Er�R��	��{"$	�dH1m��G��L� ����׃3��q-Oi�&w�H���|�s���S臝y�ّu9%<jVb�`Z�Sb�v���3�� �^*m�r�-��r�#6�>��5����.f*fK�C���z�j�B#M��������[	��Z�΃(zO%ւ��j3l%�TD?
쎔��<��W�ώԝ�1����VD�UѼ�꺖s!G3c�/x����b��<[y�B��jꚔ��Ǝ������#��P1���3f��L�E�f��V�Z��d�R[���3�zǺ���Ң�z�ׇ�]��o��1w���PMȘޕj����W�#A�f�&�3V̚��ڋ�4֛���>L��(�\�T{cÕ���&o&+_�-��1�2�!��Q)���-r*��ƪޫ���ĞC�b6�_��b���%�1F�;��
����	�5ADY�\��*?p.;2γ}���z�Z�K��Eg�ɇ��Z��6h�Z�� Z��|j�fAE|*��ç��#����DM8��e���Rܬ��j,dzy�>�n��d���n'�e�|���e�B�K�����N�U��^bm��ǩD�E63O@��֝Y��,}���o:dd0A��®TTÊck�L�λ�����Lĳ0�7v����Ư|=�{�"c�l3}���U�1��39��t
��0*e,ڂ�r;���A���-g]���`�A3��"��H�$#�
�	�њ�f1��E2{��ʡ�GEƦj�cti�3�5>|�ū��«��TY��<W*܄
�����>�D�;��͉>��7��$%o�W���hvd3��8b�U:NЄv�@%�E��+�sz��(����c�h�E��an�:-�����Z�@�4�ZS6�?wUq;0R��L��Ǚ�30�T�gE�S�Z�Cf��^h� ]��,ż����ݦE����ϊ�Y0��21�·ɞ�W!��Z͌����Хdp�� T�{�7cZ���R��/����������lVC����iƂ���Qӑ�m	�*�#y�q0W_3��z����!�#��HM�g���k_*���}���S��H?�?1����Y�f�Ol��:�=�M���{zUc2�Z��uU+��Z:/���>��q��M[�5��
̱~΢��iv*�v�z!j�;�\����~������n�~^TF�;N$;���v[�ҤԢ����.Q�_���������\6L�4X����j�;�Ab 
bӈVu���,��`�;�9�6�����ކ�%�X���j�MwI��J倹��S8���g}j������"-��������i�$�f��戴ރXP&e1��*��s��cu�Ͱ�T^uH���"��n]���B�=�����!۱�܆Y�!�GE�?D�L,�LN���Pm�D��d��ƻ-w��/�w�"��<h}c�|�&�(G7P�	�݅�<�x�.,4��iQE�����(6��j�),ؾ\w����+�W@t����-e�=#���C	�@�\�%�hk������d����ؾ���z׊k��q�b~+q��x�	���2���%���R�k��=��P�sp�#���q�AL��R��K�P�̐�њ�	S���Y��<�E��Y�]S�Ԥ��xn��Ny�m�,�;Q3:ċ�bA��g� kC��aQs�p�="���A��8��]P��z:�	�}3���3��zɐ�lO��%-4Zو%��ќF��x׎{���W�G^݁��ţkg;���d];�w^�F���4�z����Dt������{\\Q�G��	p�0g�˞5(^�W։����2�I��K��0�T�T�zuC�O��&=rf�js���]� g��r>4l��`�����M��b�	�Ҁ ��}l=����o�tr"�������g7͜źϾ|N�\�{d�MK=ՓY��]BKV.S:sJ�2K��0����1t��^ڪ�x��ۻ���O�ﾪ����=��9�yS�,���Z��*^������aR���'x=��?�*�J­��n���UX�EF�f͍}��n�>�DY��v�r��RO��Z�p(�x������S�^��G^5�B��'��I�Ƈ�&�M��yB�d��6>��i���m�O�P���3���,��P�>���9�L�v��W�C�W}��:�>�֬�ZB���Ed�f���w�r�2��{�3Ő&��
|���
��	�t5��v��	�n��9��'I�Fm9�6�ϊ�绂�e��?gzb�k��3;�<���]�ؤ�hNt����{s��Uq|	E�'�ۑ�z�W��T��~+~n|�x_E~?v��,�$A->�0���9�<*���گ�����	0��q[q�¶7⎽��y�=����^�--��<�Ĵ�ސ�0��ȗ�����<[�)D�{	�:ާ1�v������q�J����v+f1����n�JJ )���lJ��R��oV�<��9}$[�D����x+Z-�46/�S٨M��t�9������/e�ݶ\W�G� ���< ��0
V���}%Z��j�_���zfՌ�1 �J*�T�v�̠���x��[�����vY��?�\�jý�nWm�=t�5W�(t0��
j.L���Qi�gy���b��.�R�T8ݦ0�Å+F��x��«��=��]�� h�٣��(J:�w6��NwI0�4!rs�}�s �[x#z��W�u&aajv���5�t̻�
����M����Ktc�[ס�s7F;b�ͣ[[w0�j�R�A���jQx��ݷ`KT����Z�:�6r�Į]YfD�u���]ۜ����ͤ��Z9�O3�K��X(�s	p[cv��u���P�os�c����׽��B͑\ϖ_tM�%2��dns`\��K*]O���.����n'g�zk����cN�I�ŌE����lL�n'���[�����4�㨧9��)ޭ@m�vx�u�	҃bd�6����}��Hp(.�6�M�kY��P�N����[O�֓Kt���ҧ�\S��S)���� <\�]�G#��:޷�据�ݮ���T`�4a�xF-vZ����Ӭ����ݬF��ti'�q^��tFjZ�yK�f��ˀ/��˱���͈l������u��|��%A�h-wC�l]N����Wl��U�Q��5֍�1������z�l��%�Q��)��ꎖ�����Gs<P#�/�D�qM�ݵ�S�Z�X����!��c�/S2���7�򬺝��iKCU n�m�J1�U��^~�!��gr��8��zb�I[  ���4�p PD��"�O �bT��D却=G= �x�Oq][�*ݷ�
"K�Ś�� +kf�[Ý��4i�<l�R�md$�%���;h�)ne�Sl�:^�n��j��Т�ZD���o"�n�܅JV��	�t)
��zs-
T	k��Y3w����� �u��_K<���.���x�I���K%�!Aaՠ�����+�YUχ�GB���Nu��EF��0	̥��Qۅ�Nq\ŗsaf�� 5������:������U۴y�|��y�;P�J�)Ӎ#c.es�9q_	
GB|A.�9W\��M2P}�G`����\��R,�[�9�H�>��2�偭#�R��h:�]id�����}"Y�r'\)f�.c5{��>���:Th|j�;��B�i_fv�YqԛW7��,Է�'�{{#ݡ�T�me'R���'�7���+��P��k�]2���IJ���zQ%'y	Ycc,:�M'E\u,{s.^����-k:3Ա(�/�X+"�(��>��T�,����F�J7.��k���[9J\G`�H���eR��;j�鱓M���y6�ےo9J��]M��@�dkt�!؎�����.N�-���%�w0m×o
�Y�����5�WN�����Eׯ�s��c�t����g*�%���ïB�Ȭ&V��Vf�y�ڊ:n�Ψb�k�T���V����:�[�f}|�tL;��!|Z���:I�"��Dml��>����.�XDh��a�"��kAkK���#��p2�eM��C�QK�$[�	�|��"7�qh�8�rn671�7F�#	5�s��NC�Ć���A�F%&�7-N�ɨ�v�5��A�
("���r4A�6��7:�@�j!��ɠ0��5!�Z �3��W-��ĆXY!fsR4rA�a��RV�.sWR8�&%�	�`FF�
��)��F��d�T��dSQUH�a�
UE�1f4�թM��\�bDF�2�%�M.�M�'Y�]J�o;����2����C�NMQT�1\������*�����d���h: r�*���(N�p��0rL�(��r�fd����9SQ9�*
@��G0@PE(�J�WR���o�
36'oǗ|C`ZU��P����E���ֲ���8���
p�;�M�`�ju�\�1�}��؇$�̡�����諭���D`����u��J|�h]�U&al�Au����@;l����_���.N����j}}�F�'����W5����3ϑ�hu�3���F�1�d>�Uϖ��q�>�v��O|�{�Ox����@�!8L���vН6���q��{~��\���ϔ<�)��{?
���f�ߥ��X���Y��S��$��m0�1=���LU�lc>�����$��,ۅ)����Lz�f?.�������$�3�w���Er�	=`(ԋ��"A�t2$�x�tb��c�!��j�qC���^+�2j����7�i��L���Ev�%ב�}!KS������t����5��/R�R�r,�Ƽ;!VꚆ�tC�\���yR��.��	A��K�`��h�uxa�Rk��+���QS'�]L�{O>u6°�\�]P��(���'k��
���O.�<���?uч���l�����տ�9�w���i��Þ[P&{������sr��Oc��kv�nЮyuO�ܠx���,ؕ�P�,�Z�X���&�xQm�N9F��Y��%�*�7mWn+�;utk�(�8�~�N5���Ԕhn�I*����#���t���=5U�ލ壸J�)N�����)m���de�u�����0�p�����X|�G�u�EXU�H�7O��\9��61��B)�0�Qث�{޵�^��]q�Q��G����֡�km��*|��V/^��fP�����B���ҭT��������.ɣ:����B��7�Ǆ��BN�yeϼ���f�mɛɎnk�ǈƘ~=�X��y\C��n�F�sWZ�8�;S�yÔ�Q5)�|uRYbKq�n&:��\V+�l:��]�Y6ٱw[���j^��eB`kq|h���+���㖫�ZFK%�g�N(kgֹ�n~�cW���wWu-�[�W$<L }v�#���;����b�UW���_T'�,��ƻ�c�����0�eWd��-�����D��@� � �[	�|���FN�H:IX8���N���g��9�%bs�^�=TY�;c�j�Dҁh��X�	���_U�2N����yU2V��p�t�FO���f����N��!�2/T�-B�%��cH�=1.�F�,r��A�>�░�?sy�>Hk+(j��Uf��g��4Ԕ��D���Gω���*I]nr�5>�l��5+\T�Os�닷V��;��r�A���$��!�t�<�8˴�LS�^�Ȕ7�I��
݌^�8f��\�n㭢�w�a�%����`�W5���M!���|��j݅_�^��YZ��jq}��x�n�n�an�"q-�&����8Q��o�u�"멆���SP��>Ս1WH��]i�n���γ��� ������H�r)��������!�5��|����DxklcwwL�5^t�0���6�!"K����p�ז���9�K�ÇF��7��M�]�Ƣ�|�P�T���X��-�:l���t����y:.�M/zڎ��xv��;'~��T`o�	��]FP0�{��qT�C���KRZz:��s/#���[��}I��̱v-���|K�PJ�O�Q�U+y+�w�B)mutD�І7�]� �t�Bn�J�����u�udP[��
��b�Ḻ�w1^ޯ�c�zٵ
vs�ޘ�Vx��Pz�T��xNX0[ux�x�c ��&l�|���P����ߕ�BtY��=��R���@M�����H��9�E>�Z��ч�Ps*OS��G�oW�㪖�.
��*x!t�&gk'�'{�{,��"�U��A�^C�*�������s�p5�{+�IYp��]�m	�"&#�Ɉ.ǟV��g��B�.n�a9LgE����8��Xs�4��<�J.�/'�� ��f�1������w��v��4[wB~~5��s���(އZ�xD_[�\n�j��]5u�橻5���Yv>KuQ���C
�G(;t���ڤ z��|;���UhTz[�Ѷ�6�5)�z�wEh�h����o&��C0�es�a޵ף�7�^�POt
	B �(��&:6����E����mc�*��]%��u��v!��(�lp��af�W&mfFM�}��7��=�z���^k��\�'�hu���2�|��}�:���{����u���d�>���Of���y��``��/X펕�:C#*#�FF	�4�f��cL��l=۝�JzDv�#yAA7 �q�3�:jP��B��`��e`^m�/
n�6�TgC/T�*�9��d(/ټp�t����1�8�K���i�d�_p����,����Ak�x��з�0�B�3����fC�
~��.T1RO�Z��4����9s��qOp�=�V_f�G6�a�B�W���ĕ%�=%�M��jO���"F*KڨB�Gz���ܴF��fBZ �Lo��\f��s\p<k�%�e����
����<4�pܢ�BݡS̠n�b[�kA��*����Jh��&�ls�Ǯ1I�>j�O�1H�Ң��a�[�R蘃�ּ���nU�G+�1�y��N���`<�w�ZF����K����5BSĉ�m���v��Y�9�'���93�"�Ǽ�f{��{��;އͭ9��k)X����[���*��q���V�\���zT@Q����8��b���X��#��s��>�2�\T��g�9R�q�8A�`�M}B�[����e��&�.������{����+J R"/��on���������d6�;X�5x#����g�a"
i H������	w�E��;�G�L����/"9W#����q#@��Kht+�_� {V�ܨ�T%h8|Q�wq���=�a�˜��a�Ry�{Pk羞��W��4d�7]�~�$��fW9��w=�b��,ҫ�1���ep���N>f�ۆ=x��i/a#%��g�-���ZH��>�;gwV������R���;��U&�9����{�3ٲߞc狟�s�F�P�q��u�	`|"�X���t�vy`]ƇX=�8�FE1�]AFڋhM���P6v�e�s���������p� �%N$M�i�{�r����}bnۡ���a8�_g���@��4�^K!Ў��B�Ѕ�E�RQ�j@E5�^�`e�.�|�/-�w�(�7�6��2�r�~�q��Q�}�$�3���Kb��X�'�	jB��=,�������cVF&�Pݎp?�2�*���Y���L���bɞ�R*{g�v8�.��%�/]�u�e�n3�,�'\�E���.����;y{<N��hi�j�S��wEE�#;���Q���vc,+5���6�V��ݮ�7�mf�ĆfJ)��NY�,�,��TXL��i$��=��[���c�W����R�iA�Qߛ��ָ�;��íq��xioaM�8v��ܪ���aP�� ��X웄�b��L��u���u��j�����w�P/G[Ȼ���-{.�uj)>�YB�7MJ���{��v9�<i�D.��#�p�u����J�糼��ǁ����L&EԞ1��Ƀ�qu7}�ٵ�tN=�%�V!ʷ\]�ʆ/!ԣ����ك��-&)�3��̃�I���^�gn����LN��ٔ��%>���i��wA�g]9T-4�V.D�V��=�܂5�.�u}鴢��it�m�۽A�3���QL�����v���.(b�t�Vb_hδ$%,�ͣ~����ױ��v���S�5)�|�K#��y��R��zsC��|��ٱ�}5R��.`z��̉U�h�G:\G7S��^m�o�H��hÊ-W0�.���v0�v�v�{}n1O++E@HY0\3���5���w-�?e��ޜ%R�aoT'�{PL�܃D�<��҅�3|d��w�^�� ~W6~P���	�C�Bf-��yfN��k��W$5�zlFpՑ���^���J�R��k��d6J#�&�9�n��ѝ������r7Ƹ��#BQw��[k�=�﷖
ۨ�.U=���ޭ�ܼ���.������|��fjh���7���-H4�O�\Zg���;'��Q���r�=S]9&��}_�����JB�A׷]�/=y{u�{��d�EQ��@I�mb^���v�^j͐�!ϳZ'|�=���71�03�O�����l�ݍ4����l�i���Q�@���-@�DT�'����{�������dw�����5�YYY�P=�f��lwUq��%.��,��io����aE�Z��/Ry"&zoP�&�{��~�׍�J��w��%���F�ޟl���md�e5�3]Nuݟ�,�&�&5�_
h��*�j{�n�y�FM{#N��\˯X{�4�]'ڽ�j�ŕ���=����"27��Lc�}��/Cu����1��~��2�V�O`��ծ�����ƀF�V=��Щ���쯸�p/��{�����]v�ѹ�
��uTC�D�k-2kZ��T�̨�[���^+2�߱:�^6�b'�O����[Q����վ`�w���޾�]��A���W������g���\�}�m��ec
*/&^4Rui�}(��� �Ϥڙ&�����7�j�w>1���~R��xO���Mݞ*�_�7��o��w��4�Ө���S�G�DVb�䫶�����+(���X��AI�
�`����ȱLɩ�����yX�9Fן�z{����)Ř�Eٓ�ǩ-*�f>�z��jJ�$3c"���W���@�\�*�lV�齸�K��2�y���Nhq���@�
�R)J�Jģ���f�++1�Cdׄ|�k�4F4�{(�8#NZsڠ*��ԇ���yI~i�ن꺩�&/����f�)�t}���HY��*>ԗ&|' ��ē";�z�� ���T�#yR�1Sp��S����[��7�⚡�	%�b>+��������T�v�8m�F����P����-�5��a�����Lsrؿ�cL��Ԣ�d^O�d�9f�I�!�i>(����;.bYK�&��^6t���Q��>W^v������v5��ࣲ}�:����D�F��@3J:����c'$3C#&�]���eP������U�4	����-���]��-D�,?M.
��[}���z��Z���:�bgX"���ܣ#���9������4mH(��{�Q������&G\i�({z*�7�z� �f�G�^�f���Ή�v��y�o��Ƥ3ZF	\��W�����t F?��l%���w���'�ζu�u���"xvgC+�N��#H�gN����DY��f����S�����))����_c9鍪�݅XT8'�UqTKHe,d�}�_���AXzJ��ImJl�9i���$������#��Ŝ�^�A�.רv�4d�tz��Y��1�c���q��1G�K��@�%A���aU0�K�I�U-�>�h�˚�}���/1s������ �0`�(�F�����߮<<;�91��){i��Z��Tתʖ�	Jfפ��ɿm�O�ڡI��d��s4���wR�<�C������2E�T��7�y�k�����Ȗ-�d�f���v5M4�vmzb�-��fփ�Ѿ��yO���!@-K�1'^��):/���������L�.C���TM[oV�嫡�{�s��p�z�|�ؤ�k�ޔ]f��Q�'�
Qqa�U.s3Y�xg�9I��&4�dVr�|���V��=���\}VJ�=�o�c`�u��c�)z��6uZ�,�����Wy��[�z��/ܠsIe�9BSt�h�phK��ZZ�i?3�)���U�e六��^k˴���oT觏v��}�ԎW�lL�Ad3As��6���Gg�~��/+D,�^�QP�4�"SȾR)�v2�,��]�z�-��ʔ��Ť��ȟe�*�\!0�(�7W0����ϑ�&o=z^K��,��{�2*�iV�v�nOB�ϗ�f�a/Ԣ7mMj����環c�ʊ�����H��`�Ҥ���{3�#3hg�ճ|��ݴ,��,7v�ɜ���P~���k���/�E��[4Y��=)�R�#7O��v�M=����*ncܡg�\V&ʈA2�mn1]��ܬ��tY���-���ާG	A���A��ZF����+�J��1qӍ-[V�Pn֌a�-����4ɯ�s߸t%(D�HB��>�s׶v�{�k*�*�K�e�V����&�}�v����zC�s���A�XuR;��0a��^n�1{���S�6�l֡KhJ�X�'���tb{H\w�����:#ϖ���f<�xŞ'Nw�׷��7qx�w�L�`i�W)��b����)=(C^W� ]^ȕ��z�<��mss�GIw���w_��,'L��<�Af�Uӳ�3n��6��/�7��R��f����]?��x�^m�tm���y��A�=����Ke.��ty�q��ʡE;���]ᐪ������Uf�e���yr=l'ωRױ���R;�Z�8�"�m:uB�scْ���?�^��{�՝�#̑���c|���D�T:7��ߩ���G9X�]C'�7tF=��7sLj�D��s�rEm���՗(c�.�4[z=��q�K��&ܳr�**�"e9��O����)&M�A���g��(��8�^�,̡��Y[/Xt����:t��8c�*wn'ٯg�>]yٸ��m!�w��7a�\��\���:��O��u#v6��ڋ��{}��� $	����Z��V���eS�n�֡Ϻ�ʣO������J�&q��]V"�@働��떨L�Wؚ�-��o��",)v�S����,z�v7af���t)7���.����|���t������n���!��+.���6EK0� �l�ꎳ,��v�h	��n��%��o3�|�3���d$�*Z�qț�ѵ~�n�^�;/W;�pOhz����Vo�,�(1G�K/�Q�������ˬy�KR�b��)���c�(tô�B�P�N�^RF�/s��7+��4S�Zv��J�f�+�\���b���9�陗5:<�"gU�WJgU�l-ٔi�9j�
gq���g&�^R�^�����}ԷenVKH�5�M^�f&���)�XK9 ��ON[ڧ�F�lC������C*]��ܧ��s1��8��H����]GcT�����k��9b�@�C��!Rz2��؆��g.ԉHȔbo�-Gf+��'c��r�(�F������Uæ<ʸ^96�v�{(�w�$����҅@��A^�O"y���IRf�݇��%���f�t�1ԘƱ�(uN-� �<����72���u�+��i.��঍���̆�����v2�r�<�Jk_&@�u�ј�#�Ǯ���]&*R�F��ڷY���|΀t��(i(����i&�c�W�y��nt��g�;��uL�����[X�˾���gM�t�:4���x�- �+
tO��2�F�d��c'~zV�;c�_�u��
����^Q�Y��ǽ�3�@�@���2$-�6�2�)	��)�Ĕ:Aq�Ut��6Q��Q%�<��b�6"d�i��Z�U�ޞ��T���\�aΡ�Z}ʱ7���.�Z�z��N���D�-�����q��v�$N�P�`�t^���e
O.~I�W.����9]���'�w�]B=S3��Ƌ.+�䳕���{58�+�k�;vA�1p[���W	��csG/�J��`�C����{���e;�\l��V�=�w]��I]Kl�*��L�$�١��$�ZTn�V��=\3�nS��̩�{�4�t�K�묭q�����,3˰
����}�F���6�!�¥׎՚�	.�m��S���Q�٢⩘���aW�|4��A(���Ő�-���9�U�����ϛ����|�W?���oF���;�->	�׵%�t�w�Ū���&�C���+�GW��u8���͙x�Σf�� 	qD����8���Ԯ���'��6��խ �7e�du��c7�	2��@���{�Ң�N.�ɒ�wrH`�WҲ;Yb�_A�c�r�WX���n�8xpʵ�phhJ���G��P�ˑ�_,�"�eH�y�u��Y�q��n`E�<�6ܝHYr�I�͓���v��E�}��}���F���`9�/����dP1!@PQJ�3�:����\X;�����(�eQ3E1'C������h��oX�HUR������.E5BW$D���s�9�URRPEYdQABy&F��q	"Rf`��� �k1��VIY��C�j(;�&����2)h(�i��J
*��J)"B���Y�F�'��YJP�s.QPP�EP![�-N�LC��@�4�PPTA܆E�;є�CT&���$��Z�iR�M�UP�r((��(������Lr)(
+��}K�͑J�LB�;�����7�	TS���F� �ʊ�g���B��)��EĤ���� I�� ����2��%7u'l��N����nm�OX7�l��_Ow�,4�sK6���O�-h��&��f�s��v�R����y�x�S��!��_�Uw�IC2MS�>�.�^�g����>����w=c�y��<�����b�ê�e�:'���X�mҌ�g7o61��v{�vK���Rg�J�9B`q�X�ψav�U�}���iO0��y�KN}u�;)M�1qY�Q�̩���>+���AY�!�%�>��徨��^o�߉T���jy��;2��D*���Ũ���_���B��>3�I5��a��x�L�徨��q{`؜���[W]�54j��+���	�z��t$�6�x�x�U��A͐�AJ��1F�7���Nٲ�#�g�a;G!sMͦL�sh渰	�krg�1��>sb]�{�3iy�Dv��c�D�G5y���8�Qi�#�x뾖Z���P=�Wٰ,���AmIK�]�!��������S�U��*�����62DO��O�n�yy�Ё����wBN�Ӻ��H�~U���x����Nێ��s�t$ֱ%ɸ�$B����޸�՜�n�ɡ�v[�:`x*�>č�%�N�Z�ֽ�"n�ڸAOo������M��o/�.�M	C�:���'�؈�g�Ÿ������j���#��eFw���Ooۭ��q�8�̵nv�7���W���;����ip��˼Ź�#:B�6��6�B�����y[�I�¹���r�m�+�sz�F�B����<��{5��R^��3(��!�M��	uhѝ��_ڿ���<0�a�l���^Y���\%4ՕA��H�V/�O�S�D)j��!/\�ڡ�����t@yU���ROj��-�� y�ο�1m��b�x��u�c{J���~}�4��:�Hf)�B����y�:�!��T�k׆�w��h�;@�tIaD̦;���EΨ��Y��
z��O���=}�د'sJ9;�K�J7q�Z3`��0􇑓��=��tU)���l֌��W�Jy��~�{��<�?W��ɳr���Rb<dF��`\q�p8��/!�x�.ʒ�&�[����غ\�kfq^�� ��o�^� �<���wϼ ���#���F���� �#�s �Llf�޴#s'y�Q�9�;_yQX��EBp�Wba��b6;`��沠f��M.�r���Z�׉*�_u�q�]ч/��Di���J/%�P44 ��M�C9~�t�h���u��	S��M�5&�!�#����Z_�u�ɪA5Z�<H�v%�71�˝���Уy��c�U��z/UJ:�U}j�:ʐ�z:m>�&}��g�>l��{�!Ц���p?�[C�M��ʠ:���g��U���7n��� !"�j��r�K�<�X�S/o��B��X��r�j��-���b�z��yߩP��+μ�J��۽yp �g9yVKU�a}���ԶX�r�����S���򆜸r��u<���J�pDfKK69���P�|��F�/3�f�;�>�˪������_����7n%�/����B6�D�n��a�
��ױ����`��Y* �yݘj!U��>2E\o6z��
�,�ȠQ�����_����D����F�2��{��4�UF��Wn��N�����x��LE'������t:%�8�)���k�G[B�̜��k��su�u����3m@��1���#M��2���*�$����Km�>�&�FcQ�{��:2�MG���z�X,�r��P��\��k�	d���_w<-\7
��5���
�r�����u4�eԄ^F]]`f��/�]M*�[�/��6�ek\�s���/z�k������h��47�`��0Dwk�2���k:����g��sω��b���է��u3�zK���C�Ϧ�x�F�g�8��N~Z�/w������O0��(���ټ5M��z�\�oB"�K��ˢ�ӓ�P�#'kI7&Uk���TY�o�@�����a=�[a�)�=�/B�^'��Ql𝝯���0Qn���璠Kд��B��@��5�pd0u�~`���jE�˃��U��߮�q����75���a��l�7Yq�j���{f�M
;�0v4�'λ�=zB�Je������QU�bu�WҖ����(��6���S�<d��~�4Ϭ)���#�����Zwp�+���*��m����fŻ���^�P�8ܢ�ǹt0�kK����� �C:��_)W��9O-�,�p�)�B^u��H�y�H���&^����^�����[?G�f)+r}p���!�qC�;z��=�I��-"��ڤ�.�&Z��4.�,�0�u�QiOcO��<�]�֝<Q�-O�u�ty��_NZ��7w�e��Չ�/�Q�H��2��&�A�{]B�%s�zu�ʅ��f��W�OU5_��KMr �$��F��ӟJ�s��J]�xlN���������C��ÿ�br���C�5�R��i����@F!Ǳ%:1�W��zU}�k2[Qr�㏘�/�{H����J�d{R݂h�8�ʱJOi@��+��)!s7�v��BԖm����>܎L�(,���Z1�J�vyFm�5W5C+UY�����/C�<���.�''���^�ƿb��n��{�:��ro�H���z1`/���n)ً��~h����������%�*y��S�VK]�-�+��xaP�9�D'q/m�Q۷UY!4��P�J���"m_R�o�`�=��Mݬ�IP�N�N��Ԉe��c(U��#U�]g�
�Od������s��]�DH4��\��']�4]�=��񈭑�c-c�`����+�y7�q�w��Q�����������U_j�s����/�����T���L:�F�u[h�������Ef����)������c�M�s4Ř5Gv�T*ne䠲�a�OخEbS�⏵eC	��e��oi��l�)�TN5\u�������J�%c1^9\��d��3+���O�7�V/^���c��cF�6��6܋�r������Q5�^���J�qзC�����ή����o(�زʟl�Hݍ�3�0���8�{Y}q�#Ѵn�(�(��W���*�<�/T�7Ɠ
Ԧ)���Ids�xy���f+g���8�f)Vfl/��C�\Y��-�j����*4�L9��b�w�h{׳���\��U]h����jz�;�1ܱ�ן���/���hbh�	& =�	�k�����G�;8عU����9�Opӻ7}4����2�z��,��Taq˛ұWڈų�&WC�C�|��p1hA;]���S�
�Z�oW�y.����Q�qRj[Z�&-��f�P��B�w�$+7�=�R����z*�6��,�Ĳnޭ6�^&3\Q1�o@��V�N�|%�y ���V�x�u���;+u0r�f'��	�X�	�e\@��5l����A�V�l�1U�#�Ĩ�ۢxl������F�θ3k��ڕ��P/C�[�̙�܏jWM�Y	Д�le%*D�����W�̘��V�i������ن�����Ӵ������ؾ��a�5ٶ�#�g��+��`c4��Rd�`�j��1��k�;���g�L��0t���Pϝ&���)�nVe({�)ܽyD نjLa;F�wFcu^�hX�PY�lF)�~{���X*�xRF{���ӵ=�n����0�����x�<����WBe��7����.͌��D��� ��Ԉ��F���6���*�0Ѝ��9~�z0Q-�f�v�v73���Ʃ����k֤&گ��W�V����Ѥr�(J "U}�lԱ�ږ �Uc���!��j�qˉ�l��5�J�O��~���/��oj!x�O�1}�5�Kn.�ō�{u����2O���A�m~��,(���p��9�m�eͰ��6j;�oP����K�蹁�з�Zf��0��C��nC@�M��b��UJn��?R�]�v�x���Ķ{\��|j��Ɉ�ޔY��y/ڠ-y�چ�y�;��̫�W�����o�rجX|�0��=k��lq	�|T}�
&k�E��<~�:@u5����>#���
=�+�k�+qg~N�#�	���x�MX�3��z��KG�a]xoCz �!:��Eʹ34(�J����]�"R������9*G�H��- �]Y�BZ�}�ӕ1��\":�B��]��(Г7�#j�5uf�9r�@vR�+��n����(^5~2����z]9)Ȏ��0��7�����&q��7�{��	U����]�]41�ʊť���$��5n|;7��n������s���lC���)T5 �(�届`���R�?
�	y*��FÀ�}��δm����+��J�����o&�ft�Y}��.�믑��L��7(��7Ӟ�/�}<A�}(�8
���U�����c�y��9�?Bǻ�&|m��@��\#x���L���^����,C����	pv4�]�:/U}h��P��ȾG8��&�9�?kR��Y���c��GMj��(CI��Ѧ��4%ދi[�˧���G����~��np�2�zݴ0Md��M�^�t�P�)2J6�A�[�&<�B��{/�Mው�1�_�\�������Ѡ�v�"̇�2���\��O�P%��C���#�����ur�Cz29=N\���N0O�M{yC'���'ЖM6j�v�o�n�>eB壩�n�Թ�{�@C�<�R-����H)�.���xZ��d��,[}�60U�6�_.q_}����?J�v#N<�Zcц���mu,o&Jn�w�u��-Wf�HMt�8Ǘ�y@��lj��g���Ɍ��$��kYxJ��NV��ܺ�n���M�:�ړ���͢��:H/q�h\���1f ��>���%sΥy�+_�SV�"�L�����QN�u��h�����ׯq�N��v}�O����n�>���Gג�M���պ���s���*YQ=T����I.�0 ��.��~�﷨���3�2��dK�D�A�z�>�ӓ�EoZ�a�@�����e�<c	��} A�O�Z���V.�\C�;Jd��c2j���ך���!�Q}��T	{K$wJʆ�t���,Q欞<�B���;�^��A�1����x�4�\�{�r��!��BG,tl����.��4Ū�b��$qߕ܇R����_�ԉ�{�"�0�F�4s߆�Ξv�~�t2%��b�����J�)�.���II�Ada�lf�1��0�Eb��f�]�����C+�X0���b���9��ߞ��^y�oMkP;l���`���5�q���->��U��"36�v5�3��{0�UJ;�Ш��41�-��	�U�r��p�H��F�������^�{R�"����A���V5=�;�:��S�q��\ė�4%���IF�D���������U�!��<��6��ͥE<��cI����ް�l��{m�75S�����G��� H9
܉�nj��7�۰���#[x�wv�\8^:��9��W��X�{E���)m�д2h�S��SP���P՝�+����xs���[�s��鴏����C�oVK62��H�3�f�X��M�#��ƾ[W,0��2�p�|{��<�-_f��<"������1�ڽ����ڔ[Y�Ѥ�_v��iV[������A���*��4�d��G�xb���w�`0.r5<6c�e��@�r���Y�Ô�6]ݻ̖�nP�|}�^e�S��=���E%�P�u�\y��N�j��>���
��+���W
p�p�W��)ʹn2���5�Eb~�9Ч�VE�DB�H��nMF���zNS��.��ܦ��s�C��+�bKcY0��QI����.�M��`�!�{����O��Zɴ����~
� �[��t3�[�E��&�%��Jm^Hחu�B���:�Μ��TF�R����c�C��.��"�V*V��W#A�f�f��(���E�'�\�B�lJ7c���g���-���W�^3�}^<2)`uN�%h9��r���AP��"F�O�c0�֭an�T;�\qWV��ׇ�ն+��B�d,D��8��(�9BT��!�<w
�?Nw����ߥ������rleL���1^@uBr
7&i�:�!׊X��2���ޞ���c�E����ǝ�Κ�9̢J���Μ&e�kl�7�b��u�M�<�8�24�Κ�f6��XFP��H�Y�2�C{7S�or+[2.ݸ�DK"����cx۽C���⌖K�0�P�ϭ\���E�'���1a�[�]9�2�a�<LSm��gkC_)mK��������/z^�_vJ�Z�9��1a�]{I���j��`N(���0��hQ/j��&4�oP$ⱸ��ȴ��[�5M�@�^��n2�^���4u1�Tr�h֗�A��l&�Y��bƽ�j�1{�	�>U�maMV�N��o������H��ޞ}��>������� N��GS"|X拏 ^��`{J����Q�� �ű�՘���OY��):�Ĕ�%��7�":3���9�N�h0.��9��|wC̙��"�s���>�g��2���|A���\�k�D�-�|JME��ݍk�B ���j�ʾW3J�C
����(~.Cf�&�j�H)��Ԉ����Q&���hE��V�0�˪�E��m�[]{2����F�L!<���;��Mxg3"��1
��IY�w��ΪӲ2*�=2�
�-�/O2�
��@�y�^-�
q�ĩb���Gb��Uu
"1m�:����H�|�Op?�5 �Zޟ#�"�M�LG+�s��e�Q�C�:�^�)Yr�+�t�b��vi��ʏ�=0��ѶH̘+0V�
��-WZ��K��@�n�)f���O��b�4]c&F8^rR�)�	)��JC�9�:Z�VuR�5 �7y����
���`����[4;;����ukd����ʃ)5g�%J����h��|uo
wK&�k��)���t���|�����WzZ�JK2�os�\��&��^������mO�>ğQ:F�K���U�ӝp��j�i9��P�� P��ˑ�Ix��6����8
�ؠf�p���B���X�7�a���������؍�2��*�e����VSN%�R.5�ѴHw�m�p�k�r4kz�Ǫ���Gr�@H�˘ìХ�W:�2�cbc4�()vj��Aы��-&�.N,�ٙ��o$ie�]T�[��GY@f���W��Ǹ��(��G�y[vͷ�����]�\��T\�C{NLTq'��Xu<�י������W/J�	!%v�]�������S�X=��b5�Qg,s���j�٣��:\GY���K�:�j������`����vS+������v�3&C�PؾGڝf��s#�D��N�Ye��Y���B�)_rC�� ��fU�%���L��Zٗc���Æ�MH�)�ߜǛ��5Q.\�l��+rl6.�f���dրV���)㏘%�+�|7jv�;�����]R��ee5D/��5����Y0�Y�ҽ��eKwi���`-Y�sB+�؅]n�6��e�'�c�U�-�6@;��ܫ7A�3|S���կi��n�V�Z�q�"(�y�f��#�����Z�%���T;G]�RYO��Y�v{n��׍�i�v�7/\��S�`��[KJN��e����	j�'�;��pJp�����*�5�fS�Y'Vp�lo;Ծ� �k���
��#�>�;��}+a۫�72sXF���ˍ�4��M��V]��֝�O��oj�V��{f���c�E�����v�{WD�u����Wv���t�h�,T@��+d3ܘ��LB	}��A���${�3�J�[A�t����$��ۉ����|�����e��U�rȧ���j�t`cw���z�i�I69g`���5 �,mF�2f��j� 9����ծ,8�uʙ���I�k!�F���.��MmA[sQ��l�Vf��ӓ��Q,a����J̏����C ����k��]J�=沅^s�-��1�d�/�I:�p�� ^gaB����X��h�d�b��)r{�S��-<h�laχd��tu�<�V)c���j�g�9"I�co(ҠwE��ˉ��Y��T5��y҃�2,	�D�w��u>a 4k|$�O[ÛٔIRM6��%��cE�������Yy.������8Q���H�'���\�$�I>�5u�v*�VP���ֵ�`f����E%5�L`�Rd�D�ՋED�M&� �� ��*�y����i
�¢bh��QTYbMAQ&�&�F5R�]�!�c6b�I'�O6IUM=Yu9SRDs�2ɘ��\��754E�2b(��
Z5&�c5Q�̜��"�������UTAQ�:**gU9�a���9�������[����x�$��ZJ*����J`��"�l�������H��k�����������2"�*�9���Zh�"$"a�h�&U�D�ADPUTTPQQFHd1UAUIK@UQE5M%Ds�0QPM�����$�hf�7dE�U4�F��l��&��
	��*"��h7d�MSR4s���$MD�")f	���`��(���YDRt�G~k�]��~N�>��wY�oC8�֦�^7H�܀_4Xs���+��9�j �������u�V���\����k+5f}u��U��z\�E����z���>V@!����<LxK&$��\�F��٣R��@Z�8̮Ί�	�����
ܮ��3��Kr�_�}C�h�9a�F*E�;�~a�<�x�j%%5�b<�ޙ��G�յ�&���~�<k[i"����F�`\s>�`eꐽ�7{�����aj��#������X�z���ְ�}=`� VP*>و�LМ��xߣ�acii|�Eϼ���lX�Cz@��ň*99QϨ����ɭ{"��C HC��5��ޕS/�����YGX!�n�YM���0�P�l�%ܶ9kBa�@h�}�"�'�(=�Ȼ
���D�p`��HC�����>RYM�ѼΗ�/�t����͍ڭ{�D�x��>ܱ0}��=�r �#b �ڸ����x�z��r��rC�&����6�l/L��b�<�Y���(��ƾ|#��~��)2�6��	q��,&p��!F�ls��T8T�B�K���3�*���tRՎ�Fz(B��AlP(�!�r1�}z�L�({z><}G2]^SD����N�l�OE��Y!���{ɥ��.�EZ��J����ԥ��`���͇m���n�����R|y���p�\v�f�I�u�n�����Z��	�V��낃)�6��a��^�cwi�q��Xޱ'(z>f=���!��4��T.�L��>�F�.U�Rd�n��(h�]B!���R�(��k��u5ݗ��љ�PջƝ��Q����0ƝV�Q�\�$�׎�����B��I�e��T��4�63^��x�^�cs�W�ʖ/R��έ�5e;��VGC�V�4iz�G
T���
�H[�=Qr(��❻��u�=����<XA�
Noyy���N�}�~��/D��A�Cܙ2�3ވ�wk�4]-�ltĝ|�.!nD�!�=8�j�&���Ku�*)?X�"���՛�/ZG�/�6)/��E����x�]��R��_P���:��m!Сk���NNj�}jm������ǰ��W[�{���]���OS����~�ڨz��k)i<<��E�t�:�f�.���J�O|5mj�[�'$ws���W�i�z
�\%h8g�(<e��)Pv�S�C��.�?�l���H��v�3Sv{��繽���]�)�f@Y�yA_���K�~6H�y�E5�&^�f�0����t�@�kzE��F)y;�!�W8�S��z��+{*؝ł����q�a��9Y�y�=���+�����_V�}W�$,rf�.�RJ�[
mwepW��RM�&��2K�rsj��#Mˣy*,�f7{�/2)����܈�5@�`��kyh����IF���\��a�ïah>��������,���o.��0����CT���1��K�?��
ؾw�s	V�r͍/�4����p!P����>����WgMa����FZĬ���§ⷖ��2�,�-�l\F#E���l�UhcV�s���q#C߱#�qX��Wڈ8`�� ��X���m�m��6�W���Ay} \y)��-`9͡���z�<�hA�.ȇ*�)I�(�:�����T���sp����TU�ʺ�l�c��l���"�ߌS`iJ�5y�S:wA=h��=��*�͊9Is(E�
܈�=,��&<sW�я�E�O�|���C×���cI���L(�KϵSߋk�5��s䮶>:b}:�̋�NIOR��-��[`�r���\5�.��җ����r���;�
�R�%���C�1N��;.b��إP��u2��+���ߴ��e������b���z���e�V��핔+lr�ac>�#�h���,�C��<�6�k����[ER����v��2X�uM���=Z�/�nEf�[�-�]CǶS�8~�o��)W�%|�:���FjD_������@n�+6�0��V7���F�k9��)�P~��<��,��\!VumkA^�]��-k���ǅp�ܔɼ�Ycpev(��P��>W1Y�wN�Wۉ�{�6:�S:���D���=W�V�ob8������.��m<n�����ċt�Mk�%��fQ~ħț*P#�M�˽��X�*W<�����
]�d���>>K����C_�ܥj���j�*OZx���'A��I����~���>���L71��J�Y���s���>���<�ɤ����9����d���{��ݵ�K[q���n6:0�E�I%gң�BsS�8��R*�s����1P�Ӑ\���&��1����=ֶp����}���H2c�F0�qi�w��m@���z�K�����bݱv�җaoT'��;��C��Mh�A͕�+%x��f{ ż�͵J�y��p�2^�����*)��IomP�Lt\ ���}&����g�`�Y�𙋧�v������ ���JCϋ�c	��澸�I��i0f���C����u^�~o�}��OM;ƾ�g����$r3àx���gH��\ު�&D�Y�9W���6�l�iQ�~�����g�{=L�v���hϭ��G�쟁��zoP���w��-v�EW�Z�A�Z�+�BGw�E���9%RS��`2�T�q�Y�݉P���*�7�VLou�J�$��R�+�u�cpa�,�Fi�c���h�J}�E�Ⱶ����0ю,��:g0���l�W}J�Mm�ێ��[��ݧ15Zp�]9x�v�����MJ5v?��ι�E�w�N;�����@ri$�� vϊ�C&]@DIr��'�
��\�Y�Ȋ�әHV]�#�{��z0��K_��t��Z9	z����F��H�c#b[%���qʰ��d��l-u|� u='+��0�9�.�uQ��|&G*����o_���nE_zb⤬�V/�H\�툔�ܛ\��Uų��� ��ڿ��:�	R����]`b�oiWt(��7{�y{���G{^�Z�#c���&B��y��לcz���@ׂ�H%�l��y!�`BV~�ƪ�y��io����3��^�=�,Uu1Z��KC�Oё�S2硛4�=!��ԭT�C�k�(,�5�[��psZ��x�O6�)��g���͛�_j5&#�czQf���9hq��<鼋�DKц�W{-)\[u���[][��L�}sz;�}=`� S���b!>��u�^T�غ��5ن�N�HȖS���X�P�%W'�PK��$wߔ��r��ڋ�.�_�Ʃ���N��[Bw�Q�\^ة���t�b������lw/ˍ1�E�E�&:~#>8������D�G�={_U��FC����J��]	�Tυ�Ĕj��\Tsi�r*�+�o#��}�,�P��ǩ���mT��&�΋�i�uԣ|�u�(��LB�4�+{i�o7��'SwL��r�e�����(��F����g�x {�C��"�*qq���|0�v��w�s��_T-�}�=�c2xN͉�<��4c#o�!C�Ȉ�͐���W����U�YBwF'�lj{�N����c�ST�&�zl�m�W�zk�ݩ)i����=D�	����t^�&�uZ�Elu�zO�6;�u�u�29�9w��H��P������ 8�o((&��0c�4˵^�������*�M�N���ޑynĚ�Q��i�����r
�j�*�T(2�+���gB�>�M����^^�P�D�9�?q�wuPh6�u#3�<��DY��f�څɮ��{>��=��NGy,k�q,�\�5�٬a�5)�P����)�^��M6^��bO�.|�9YC+�|E}�Iߔ%|n'��0�@�<�����sX�2h��jt�=�0+�qaӗZ�kY6�-�r�ƽ�DPچ���#c��]$��.��_��Ά���eΛz�zs����5Mp�����S��SiQv�TP���?�G�E�ө%㼑��)
�/�`���p{�#�y)p�;�G�I,
��C�t̡�K'������y�.�1:��v�2^Tk�|^��(�>9�3��  ��]�T��WR�y@��]�5Zo��hgӽ1��=k�)�����iSǠ�:h���R�s�g5Vzd���O�w���|7����'XO�:Iqa̪�|E�'=���U��?{�{o�o�oN^��{�z���sx�EĶ�|�}�Pm]
�&�ʰ�U�0P��f���im�H��u��T�B�z���7�ӑ<.x�Ch1��R��_�J3��{��>ޗ�����oN�O"2l�W��!�>��JT.��IAZF�ؕ��O,��ϣ	i�2e��E��П�$Rn�q�{�c�uYo��c>5�g_e	W��-&|�0����1v�J�H��B�gw"e8�j̃����,�96���h/AfϢ��f���=��x;k���oK&NF�&����P��jp�G1�׾����:��g�(X��ȌF�EJ��C�<
�_j ᄉ��ң5#��}~���=K������3:,��:���)��69��m���۽q�a�h��4%j��JO}�x���+Ș��w���.U��r�p�;t���8��6m,eV���l	\�齾��Ŗ��c+��US��g�,��*��G<�:~z)�j��,/�.�j7�
�z;���R��V~7���V
��7�Ij�KN-0��`��n���
���t^Wt*�t�����#{��e�M������������N��yXF��/in�u���S+P�p��K!�AI��l�{�3`Y`mV]�����x���0�Ŧ<��.��X����K9=��u�f��Wy�n_�7�w����_$[�mYZQ�U,^�^��k�ث�7�hǫ��{|�7.�L�M�[6z��]���˧!�Q�w��:����@�{ځ���k\NT�!5]�m^w9a������<��e^�_l�+lwU�F����R2��1f���#�&�̓ad�_y�C�c�u�ͺv7�	��t�_����b��Un��յ&��f����nS�O8���a�͘ò��Y�ժ��_L�-nfQ~ħț�^�Y�6�^X�,ޫe���hu����Q�w"~�ҭT���F�ٲ	����V�.���s�n����-����3f��u���,���>D��uP�x�i�,��J�sS�"�$,��.|�9g�`����<%ܖ���u̎��n����$�D�7��)`�e_����_���s�ݍ��1ذ�z;b�"�
GdÉ7j��;{{峄M�>f�4T$,�=�	KO�c�f���`)}�����%E?K���%�0��.2��]<��n����
�ұS� �� ���[؞�;���j�c�e��x�.�����)�&�XF�ck�:J�����Y+�(L�����ˑ�7c���q+���2�&?��� �2����5dl����b�X/[���r5��Ѿ١�f y��aʔ��;�
��t�H�ҽys�A��7�� +��*yjda��Ey���O��5���}�[�'��%&2(Z�g����֢b�ˣ�����:sewp7v�e�����͐��	���W����Ն���L��fS����4e�=�3���f�7-�\nO�Qھ�J�-JQ�Ѱ&C��"Q�dx�t�Ő5����(���X&���:��x�eu��gIق�fD��Ј���"&T�qSY%=�vצ�\e̛�5J`\�Acn1���.�v;����0,a*��P1l���0�꣦��� �� K�"�S�1��$l(ۄv5�{�Z[}}	�=y(A����Uc�y�7Náݰ�%���thbg8.i��W��Y���k%��lx`ZlV�[+USs_��)��٩]
ǰ5kK�5V,�����4�Õ��ngB�Kǒ�̄�ύ2�� �˚ �2�X����M2��X��yq�]�v��-�$W�G
�z�!HV�b��ԥGmP�������s��i�3ǜ���J�(��g���W��v��E���7�z`W��H��{�F�=��kA����j��c�/����i���Pk2�	�;U�U���^�n��C[y9��] ip����n.H�$+Ѭmm�5�c�{c��N���;��:"1�E�_apږ���nV��qv�o��G s�O#�8WQ��eA�f��J�ӧ��	��\D��r��wD���\_�Ȕ酕�E�Ч<-��I��8�/@���m0T�kW��&&m�nŰ����P�\4�{<��+�՜����>Xr���a�AhO�)����\�*�O\�_��¸��__	�lu���T7��y�����7Wm����1�Cw�ǩQ�뜾%۫�/��f!�*	./'�-�����+��q����n[�^��ϵ�f�od��=|୴'���o�@`�Y��~��PcW��Dcڶ��gS��Z2x���QN�L�qwc[��#<-�3@f�z���@f Y��\v��q^��\��@����榪j�Wû��y��,g�k�>�55���L-5��DAj��&��R:/VG{��h�}>�����t�|=�A��zY��"�*��Tt�*[
!���y�!��ڹ��=����]���z�Tx8,%������ag���P�2y�qU�-�KH"|��y�S��}i��v�`�rp��ѱ��V���N��MM��|.~�R.�Q��i���_l"<l>񐗀 ` P ��hܰ��|��ش���sQ}N��u�KE���@�%�Y��5|pރ@���%35zy�;�i��a���CR�PVT��Z`�j����P�k����QBz����,��T匣yZ�eqރ�<wUά��[�H8���Y6�k�,�c�E֝ag��|p�WK��Ў��:�nRL�`;��<}mF�y �h��I���-V�9P�����i0�����I���r���o��t�3&���WQ�PuM�'�WDS[��R����e.(�N�8e�Gs�	���v�B��tCr�M&�^�J�W6�<����ݝj:9T���t�t=�V����w��4ۤ�z���0�*S��T�07���@t�H(�i^����<�x+۸�G �rN|�p�\�MJ�Sd����w�z��2�yޙ�\T�<�#(mTS�7����r�c-�R�m5B��u��_Tb��koj�Ym
���Do6.��֍��]�\U����i{���d��,��+Z�5[��N��R�E�ݳ�2�S����	gKd`c�L��qg��۱7w�\���C��1�W+�i;{�)8���ഗgu
�2R�f�{�����d�N�@�[�՗y�	K��4�����u�:��d8\ub9 u��[Y*�E u����G<w�h;������N��c7Y�sj�ni5|����s@��z�)�U��vt�2pY�-�7�6����^Ҭ�6 -%Zv�0�F�W]����ֳN
̡��ִf1�^��{�s]�oh-\�y>U�%��� �c\x�����>I��ݮ��+��Z��m@uf���p�<�V�#+�U����1JFDJ�Z���.`�D��@�F����/���Xl�F}��)\�e#�^V�)S����$ˬ�%P�n�D����-p`Sfn����}9������{,&!�i�U3������kY�uԝ�Rk�����H<+73X�З׉�C�"�A;��=����ЌY�����:�� u�;�B��:��X#fS��u�%�����z�(���@���{���?p_&���1y(��k��]����h�����^�nPr�:�ˮ�!�j�T0g Jgu�X��*�P2������,�xCG�Q����G�*l}� �e8�*<>W�k�����<�f�t׻9Y3��,��{:ږ���3�/�5h��۹*rط�H��v�+���"v۶k��wt��PM�y�Y|��vj��TQ��»%���kN�b�:�O_O��4�3�l̳��k2gh��k�P�}��jq36>y0�J���f�
�r�{���N���҇�fbw�ѭ��G�51@���υ��t��L���b��>�G*f/�I��)̓=w�^���ׯ^��9u�ۮ.��&x�������("b�����
-fM�EUID5��cQUUV�Ȫ&9�(�)�i)���)����q���&"��.'
������eU�d�D�U��h�l(���b�����H���h"�QQ3UTEDTPTs���S�[��`EU���UE�%5ő4EUD��rb*������� ��Y�9�s��QMU$C�(��������

�-X�DUUEHQ4F�jkWF���*k������2���� ���Y�U5TD�`d���Z̪�""�&)�
��*h(cvA�2��������Ƶ�s�DE�As�Ls��KS@Q�8TP\`eMFLN�Ŋ�Xg�	��)��H��C�EyZmj������8�T���b05���a2��f�\�|sk{�'��f?,��
���I^PP%�
�Q�����ש��[P��a�#R���T7<HJK2x�����|ԛZ~|�=þ��dS�P�<��i�1�9R.�d�e�R
y�y`�أ��)i�w̮���]1K�4[���z]����}F~��"��O�XIC�VTFRG܇^��pL��mQ��Ƌ�挬 �x:��):O������"�l���E�
}p�z�|�b��z�]��(�[ޘ���1X�ڐ5�t�s��I辬R+hͰ�^�u����W}Q�t�mfã/�dw�Xg娴�\s4ާgi�䬶y�"��zO���^�-�۸�c�;P�a9�c:��@f zUU�,5�W���}C��
��v�W��ˢ�3�3�KYgV1ƛ]y��_�qG3�/q�m	ɏ�B70�D}F�2�	z��~7�:���a��uJ�+i��fw%��x��n��.{gO;�-��ʔ��8��s�<��њ�^y�{��aS�Ahi6��͝hټ]��϶�!˨�ձ���z)3\�v������� 1TlZ~���`_k1m�pU���U��l����&�Nk�ւ���œ�Gy#a�r��))P��e�4�
��:"�&�����P}]d���B�5eN|�|�4�-�E�1�A�!4{�8���>hsg��|����Q�r���5^����ǽq{���Q/���x\��Li����-�����\�'�#C�#A��MsP��i �$�{٢>�%��3��]C���4�;�a��C�:���R;U�j0slu��vp�Q��@�Z�G�Se����\�vV�/a@��@F1{��Zw� 0y}����y����&W���7�T��{8]����Q�<�(�Za'��Z�}"$	�dLLx�+�~���M�iB��:����U�U��>\E�?vz�[�Iv/��`�-H�#���(3hI�7�K(�M����4��!�F�D:*82��"��6J�w�f�ጻ�U��"�#�����:���tH�o	7����X�:�fn��j)>�+(V�gU�F����S��P1f�ޅ��t��v�5}���U�����5u,�ɉ�ƿ	�{���P����8��vQFm%oI����:E\0��E���m���3����j5�o����_L$�a)�'
�7U��ce�c����;�㞈+��NUZi
2��LnʵA�b�h1���f��(���E�pk���樦Y,���5�U���m ���������&}弞�B��y&J�oe���i	�J��=쏡�3f�P�T�z�.m�U�e�bkp\3,e\֎BF�� 6��`�30;ע���*ʽCl�s�|�#��`���z��3|�����>��U�߆xLh��L��֤�>��1A�s�{4���O�ƲЫǣ��
�/T�������#�ad����Arf�♲�@�;��x�I��^�¹���
O:�r'N�Z}}�xG�����U�--�;����/�����|��c���n���T����`�;����)������ƅV�K���<��Gs�*0���m<k�D�|3B�\�C��|d�w尵�L�'2������'�čF=Y�<b�;TpЊIJxK4:z�VQ1�U.�A�P-Rސ���&g���q�V�3\P�k|1a ����u˧�f�݅R�Sf�xJ;_d_)�jl���ģɑ?zLg�ү�K=f�� b3�Fb/�ꊛ�o33D��ǜ�Ҹ�&�uWjJ]]S[Q8�DH���"n
|�ʆ?��RX��&S�-�y���d,z��I�>y����'�M�db��^L&��$���i��Gc�>B��W�p�O���Q�q�垼ɓg-i�T;��u#9|hTS괂��R"G����+�Kث�|�-@Cy�?�rVv��-���C�1[�P��sX7�SFg`iٴ�F��[�&� 7��/��-؜���+Eү�uCRwe�������̴������i��±i\2U����e)�[k.P���t"�Ґl�ٙdA	ʇ��z�}ϫ��(y�?�o}M_y���S�B\��mU�9��tŬj��@-�⮅c�խ"��5ev�Ŗ'�����Խ���|)R^3�V���fڡ¦{�`�Cr�Z{M+���>�&=�k԰w(O]�x���i�RK��_��W�Q�kg0s	��@WYǆ)��� �����D��L!Kh�Q�"*mkY^J��s��cu���R��]LG���}��|>�u��68�����
��[ipR�(z;[��by�T�����[m�]G�����ƴX��hv֊��mr���ۛ۞%��Y��>�\s�TS�y/��Tsux��X|'�l!d�H�5�FVU��U�M]��νJ")�T�6�W�%�b�oW� ���ۨ%��H�}OL�쒈�ۈ�c	��痴��G�xq�-��K�꩖���[XC,q�c��n�p��E���D�e�1WA��d^ʀ���$!�5\��ƾ�%���}�gK�ٻ��QQ�^nh�CM嶑Km>f��Vk�����H3Af�S�b;U|g�Uɐs��2#;�a$��U�������.���Ma��/���3x٢E���J�5�ƮW}��<9ve�A����̬�H(�r1ċW	��e��Kn*,�6��'Z��Zv�!9M�ك����w��egJm���!DpN2P�+U�u�i�����F�|�f����u��-�F���=���rs�5􇾓hE��K��F����Pux��iu��S_�<�Ït�Q���9�L��&F2���ހ(��P��P[
!�������qr�sk��t���<�C���z����<�R��dv�4��E��r
���\�ԋ�	��W��jk�o����&IF��j�Fr�&��߮~��uPl=�&$oN���(�����k�v����#<�`��x.�/ԭP�I=(C^
�Q^Y�����O������YR��4s��{a���ΠsjU3S�����dS�j�� �&x�#�Y�Υz2i���H)�7/,����.��C�vk`{=�T�
Hdŝ�f��Ll/��I�~x�rd�+�Ve%�H�lc�]k�~�F&�:�yC+&'m{Rr_5E'��Sm9�vT�>���]�_�����&��H���a}����Q�$gJ�N/�J索ӓ�EoP��x��ۛ�[(���\wǤ�wW�}w���#��ˑ��фǞR(�gui�9���='ݰ�]� �^9��'��1/���EG��V(�~G=BX�a�}�{D�`��w$VvAC��jz��a�A���Q����Y����[n��5M�u��8�=��`W�5J��ǯ3��FW�pU��#����iNȬjفL�n��8�'�_�����Q��߽*�Ch��v ��Լ.z�!�
~d�6󢝫9N5{��.���lL"w�۫CH��!�o�8<=g�ٺ�7�`bJ
d3!s��*3��D�ȾR)�Y*����	{�~��e��]�������K��I"!�фLtf�T��SόQ�y��.~:�4�.�7h]��6�v�6+6}s���TW�0"�%d�q�C�A��p�=4�7�^<%{-W/FfЧ�7�?r5�cu�F��J��I�;�:�?����ت�E^�ك�haD�F�ztА���>^ډ����a�9�wO�&����z���:��uk��09J�	y�����R��$�����,�������vUtN����_".13P=�?g)IX��Ȥ�iȤ�^��ӌۓ��G�2j[pZL���dc�:8�
]���l�ݑ���W����PT�ϒ�� B���znw��(�yWi4b��#.R���Н�8zf^��c����׋�!�B3n�ݕi��i�'���f�R<��i*466�8s���OqCG/�����}�����ճ^��^�wO�^v}d��|�V2�S�ݝ��Rv��Z����h5X���L���(^+L��TOj�H4w�(֤��pV��d�|{��]_U�:�4c0���iT���5U�u��L����ځ_Tu����a^�2�7�,a�B��i�z�SΟ%�\�)�*]ᖢ*�C�sizKw�=���Z�@Q�Mj��YS�����0���)?b��Un��םh4DX{/"�Z���
,P�r��?Ma1fN�B)i=>�æ�gkI؅ϼT�v9���)����H&�z]�o��v�s������5V�BL��ҭCˮ޾2��J/}͵ҺH��:����M.��g��q�EO�i���̘ÇԭDY��*:b�����C]�����u��Ѹk�i�]C�a@���> ꤲ)̖���$B�hw���C1\���ҏV���K��d����+y�CȪƌ8�r�s�J�K^9����0pp� t���~��&��δ$���&�g���s��n��>��uQ�R�moT'X��/��.)s\�?f^�\N���r������ �G����LƗ2��#;�����ZS�q|��E��z-)��7����h��ǊkI5����!Iq�O�>��<v�WV�ٶ���R�Z�8�K�I����Z�׺�+J�O��*c_S���5t�N��8�[��IN��&�3�YfA�Gx
�+O��Ov�o�`m�h�'^���)T�
���dԾ
�X�w� 1&p���u4��7{zl����D��\���R7�1v���UG���.x_�_��2��:�t��	Gh�K�0�P2"};8^���h�Gw&�w[�H�A�vCcp���9�w��?@����3���K�dIMm}�odDt^�_zJ5q7�M��2Dd��u�v. {3$�׻��r���my��ASl@Fm�={�]TD���{�]I��;�\��Q�z��O`W�^�n,5g�E��>�Î;
y�e�����X�Q�vL��&��k�������mPzX0���#\Ԙ�Ԫ��{
�)@-�+�X��� �{�X��R������#�� ,�c�k��ӂ�7*�Z�ЧZ��b�Po`<�L�'Wn7���q�%8��j�Vbڈy�*�����@J�F�\�}�F�ܗ��:�p�^�Mջ�#�͐���K-*e���m�eͰ)��x^C����4ܻeL˞�q�6����U���°܅�Ь��4��t¼UIn��Um���yyD`�V�% Ÿiv�����{�
0�M�vƊm�d�;0��2��iW'�76_�<����X��)Hxg�pb�v5�\�
��
�����a���d�(g�#�6���k�DWH��黜�j�6����ǝ�/�jN�<^�]uz���V"��PH3�YNyJ������]J���kOB��;r�	�Tt6�ۦ5�Wi^Y�Nx�4v���f����M���:��2>��1�#�Ck�{"XϺq\��q/"$�Kۘ%��(���msJOmR�9����3ι��믄\$5<V���*0���/=S%�>�>,lwT������_q��J�1���e�z��Ay��ƙ��B�A+%� ��
��U��k�J�́�x�seg��Z[gl.��sF˕��Z2���Ԏڦk�ܣ��8u!e��d).;U}(�S�֋3}\#x`2��+/����Ӓ5����	�u�՞�����f�L-4�����$�p�"�;�S�N)��Y��Ŝ�^�c��;c��#�01�:���@�CESI�9��$lB7���ܥH\J��$e�S�6xi5��f��0E�C�M���036��/�kĴ�	)�p�����r9v����NG�<X|~��x�{ꕏ�7~���l�Ѡ߆7(odd'EZ
�ʸMccVc�G��d)��,T1ROA��]0�_~/��jx+����'$o��QQ���o/�M4�Ҏ{8KU�m�}r��T�3�T��P�v�w�$��
�������������#�n��h��9,�sk9��. 3�z���дT7�ZV�s��n`���)2�ͥqh��E��-a
u��8%y-	��y:��ju�lU�i��C���5=��I��:��Q��nG��*>��fV�u`9E���N�˘L�o3��#a����k���t��R�}�$�߰�����-�8��n�+Z�j�E�L�%}d��Wt��XXj����	��}���bz��<��Ej�p$��W��P6\*�R���`���s��p����rK���l6:��ÙTy����oH��Ul1�;=��=ʷ1O�9��M�\�����*,���c��~XO��GwN��l͂ҟ3�dFGv�8f�C1���AA��5��=�b-��	Z���L�7��7�L�r�Q��^b��߾6C(۔�=ˣ�	?�9�#�
��6��Ak��Vb�*yfˑ8��vZO�vN^��n���疒!�D�*{P�Sߗl��-��ʔ��-$\�"'�Qњ�F{�Gx�Z.l�z�ν��WD*ԽOZXJ��l-�h/AfϢ�q��j0κ���,#�b?ׯ>�&s��r�Jҩ�4%���Z�\�o���ŧ��E�#��BUW=%��hQ�fʩ���q�1��- �$��
��%M���a�T;������)ހ&K��H ��X�rZ^�{=��T��#�t:����К9�Y��>��wa����q��zs��&����#���<z��*sVb)-�z�����u�����,Y}�1Ziܦ��(f-����$̧�}��������~'S_
�� �������_I�VY�D���+K�3+1�F:^���W԰F���Q��ڀ;��Q�a���v)�Y��$nx�[E/!��j�w Q���g�v�O�x�,Z�_��L��2���������0P����l��b���|z=.�nT��a�Jm9m�Jo"�j�t�%���F!m,�-�i2�y)��b�y���T�2�����v[��
Q�Q��1T;�gi�Ll^Z�@d�n(f����J����Ẁgf�<�<�@��1T�M)��v�J8�`���/#�2��.���T�-�A��B��e�twH"�2֓��ё��Tz6��,7#DsOX·>�"��3G4^CL^EjѴ�^fJ��[}J����u����Z�j;G@a��-6	e;�ā�Y�'G��8+*ڡ�-�(!L��R��a��3nt9�zX,ͥ٣7�6m�1[��j!�d[�B���y�=��"��L�±hc�b}Wf���d�jĆ )���u��}�rl:vnjV�H�6�e]�'-���49�';����L �#0�A��h�1��͸��$ҷ���9�lKv�m������(����Uĕx4�CWj��M?ۺmi7apT��u*5d�ZC)ýGS�<��4�u�͉V/V���$)SC�B�P�P��J	��|{&��7��Ґ�B/-6<��)��
�b�Ʈ���1Q���ՖX	�q�N_N��e��VT��u���R�a�
b���+v��e=W4>X]�ۣJ�V��Qy����:���Vp�%�˛36cy�Woq�n��
��c�z�s�N�̇�������Ӆ)-��`�ŋkFu�KTf�t�Vp�ҵ��slݣ�uv�l�@P	���#�����uM�5G0�u9�u�D���ݔ��*N=�(�h�g2������|������	[QV*׶M��:�ǉtL�S�أɽ���B���lO�V���ދ33EY��j��)vZ��s>��wv�Hl���W�L��mU�O[���YN�^η���o��&��@>�`���x1�a�z�l����FY�:��q\�J�<2i8v��n��Qi���k�ܻ�]�Hsw�����gV6�E&�h���:H��q,x�ȭя*K��m��}��X>�KH���uP@�ԣ���4��uo�
�dذ.�8Ŵ���5%,:���ܦ�!���y�oݼ���_K\u���U�q���ݻf�E��{
XA��8��V�M�W�[�$� oTe����X�[���^P�Qv���puNgm����:Z���*�WC8���
J-YP�T�����^�w1o�e�ئ������zRfﲑ�g�dӏ��"JK�d��!%8ۏm�̰���`  A�`�$(��7�i�s2̻̈�F�b�k,(K"�b������2�5ѐY�eDfe�fF93e�dfedb{�Xᙙ[�ֲ-�OPd�)�Ȃ)((�0�*��#�Q�d�E��V�ʢh��
ݔk0��s(�i��X�LEf&u�%����2H-��%S��9�AQ:���+�0��U�c�S4�beD�TRLSTQL0PDPQLEN�TTETUAa�LR4�To1�	�����0�b*��
(�j�j�����1H���'	�a	�8�T�\`bD�SKT�PDF��bB��5a$T5̚H��(��")�(�e��D�n\�J
�("u��z�!݀U!�aQK$QUU�R�L&�����b&�������(�][T�~>W�*�*TjЋ@�-k{;�ӣ�Ɓڀ��a�쬘^"���\8 �;i�.��	2#�(Ջ�k�$I��虺���ˏ��K��yw��^]�{	��[�Y�n~��L	_����gV�C��⟨/c�[v�����:��Xa+�
�*�DL��/7'�`OB����M��E<Dm����62�&q\��c��c2U0�hͻ���j��<뵘brJyե+�륅Og����$Z�qM��C�G����ˠ��A��-����<�ۼ4���G��'O���{u�ō��wU��4��4�(_=�0��=�A�?Y���d��CHdQ�{Φ�~��/+J����'_�v�B��W�ǋ����"R���SW~�y��[�{/%�b���Q`�&muy+�XÝ>A��"G��_|~�{�6hJ�(O�ZLS�y����kĮ�:�����)��Y��x�RA���^*��컠�2y��E�Aw#zU�:c�mz����3��#�؆�ͫ�`/$�V��מ!'W��Lu���"��s�w1C�,�Ǳ\�1>�KUƃ�2�9��ٱGǮ��^�vz���q�G�2�a�Õ��
�Cѝ1���\�,�4�M��nST�:�[��(yF��,�y�n�����1�뫺j�X�;їAN���A��t���Mo���QѺŭ��k��`�>���DAi�}7��@����;���1�z �5VV�WD�7I��p��,w��˨�ea~�[4���ZP5h:\�l�b-8�����&��=_�g���K_�4'�v'�W�L8㖩�7�XH�d���W�:8BW�����������=�]f��LF>�L�Nn�����%J�BިN���_:\XG)�25�6oh�����<�w�D�NA2	��>��>�5QL�Gm�qX�	I�����*�+�c��<�x��\ʮ�]Qf��O���D��@-@[��㈑3�M;C+���W.��$u�>׃�B�p�1�nT�>>��-^ ��T1�T/T��."$"�H3����X:/2��(>�����`�r��Z���<�ҳP�}��[RR�PSZ����7�"�	�@��ZF�n{(����&��>�k���ú
w/h̠sj+�|/zl�=s�PɄ�7>hN1*?�fUiIJ�v���_߄X)��ʭڵq~ݍk���KCM�0�┠�f�����L{�	G���J3��dF*1Ȏ�Df��0{���5�ڹ�g�j��YB9�-HM���.Pz-|��k~����2�����#�"�;*!瞝����|�fڽ:���.kūzUkxc6�+���J})O|ƕ�`9����(P���y=e��(ک���\C�5�T��u�!�B�.]�OJ��G��b>�]9��`�}`���k�k��$�������.F���ZFuE�(1a���sr��]O��4�f�#������(\.��5?|	�c�v���
Y�37e�����U�Wj~J�Z�[�]���Lڕ�X�-!��g�
�3E��Be�
�b�橶�Y��(���y�)���l��d?��ɕk���m�A�iպ����/��Jt�ҩ-݀��A�&T��-3�}��t/pϾ���Ն��WK�j�#���7f����2��sJ�;���5G7
ߙ9�D�{k*i8]3^�^�w<&
8�ޕrK�>���P�Gb�oM�/B	S�˨%�^��Y����kx�_�þ��|_�#����h����Iqyb�����%�=����ZH�w���؝�����p�P[y���y��]�^J����!I��T|~L��+��K<z �w��p@�e�]:_�Ah�s�iD�kP��.ƌ0<ҭ
���5}�a���G �{�ON�ͱgx�^��|������g�
�n�Of'��I���"֤K�T��zAdJg��9��,���^�T>9��GH̌eϞ=3�Ddh�S\�)g����ꚥl��_)f�y��pܺ �uʅ���U��o���\��wR+�=-;����Z"�����	7�ic����ڷ��ߞI��`��O��	d�՟��]�y�̌{�I��}��J�V6��;(9]$:Z�;��5=���+/� ����猷������ �Ͱ#ZD�Jha�E˻Y���ݦ���g�Ii<4�'6j����3��b���ꕪ�&e(7 8�K����w��*�?�'��	��Gz�/
�>*{k�ˌ*a��1j����]�4�q�=xܺy�n��'� |�m1p���{��&���{�KgSr@�������r������M�5m;	[�ʒ���;�+�.E��p���w��蘒zi�ł8[+��F��Mn&x3��p�T^���0U\�4C�4�T��{���K�}o��DU$]}�9��Gh@���¢��|���g*�j/ʨ鳒��&AI���1=���1rV��/�ؤ�k�Δ]�>�t�
�J..DVy�zOܵP��nȵjz����ݞ1t��d,��{�g��1��L}��~L9gt�:�f�^�l�.������؋W�x��A��hu�WB�n��^x�pj^=K���e��(�{Ez�M'^��bN���e�;�p'�r0��֗e8*G;�0C'���kr�@c̾��q���el�e�R�kfG��l���AD�yʰ7��{��#r���ʂӝ/�T��3;�+���^:|�,űӪ
������-[+�nL�-9Ǫ�zL�$g�#]�N��L�Xc�9g9wi��
�H�;w7�=�l�`p����f]<u�i3v,3�k��E5yb�/G.SJ{H��XǡcE:���K��<��ֲQ��}�+Wݡ�S�/%���y��B�R�a[<�ʾ�s�z�͚�C\/���"�U�f���
A^����$RҸ�mi�oa�oI�;M,bӌ����8��
g^�o%e	v<Һd�E�8�FB��N���-�B,䏓��_HYkk�s�����њ��1�4��~՞x�_��fZ���#��y(JՆ|Z��0!Ǳ@<w��6vF7_?b�@�� ��ظ��r�:��O���5�®SS���V)I�B�=#�D�9ɫ3h�y)���κU��#���޺��rC��PY���c4�u��wT0s���E����w����-L�eVDo%l��]	z.-�HY�&XلC���]gH�td�%=���ʅkz<lc른 îi뺝�н��H�����~�4�/2�/Z���Ö��UȞ�6D�L�یs����z�o�!9�&z!6H��,����~L���/|K�z:��Mm`�LK�(�Q��{��s��ب���UyJL�ۤ �,������7;�J\\�)֗kW<�e���n���o�U�R��ěz�R�V�(l�xۺ.���x�ah^�h�l
���ۜ�jU�9�\I�7�.���;'fP�1���WNP�ɚw��!f2�6��ۧ8���=͊.-˧U1���`�g�Nb������oj�g��mr�P)-�p3�e��Y�W]-^���׫Y�6�9ml�c븦l�z��V�Yhh1�WO�.'T���<��:)�f@�I.^!G��k�>����g2b�?6[�x�gd˟�;W�^[����]ݵ��<B� �]�)�!�QA��`L�m�NjS#���Ԕ�p���+	��#�Ќ]�#��d�GRC�[��ZԄ�[*���<���O"��ч�r�sH�d��0�P�ϭer�.s;��~s�z�K]�Q"���ghLG,1wEG��8ػJ�.;��z���|i�{��VLYdbC��m[�rz�c���� �ܮT�6G�
�	��*0�m�QL�/��z�6�f�͌:\�i���8礚�Eⲫ��Qf�c�j�� |�Z�h��V\q}�{�L�:��ܵs���9��N�wE��tc[ב�)�ک�K|%�2/T�-B���*���	�#}�qV�C����(#�.7>��r�9��~�0,���٤%T��sRR꼚*�q��@th��*�38��i=�"�|r��#�[@�*u��
�Lg���d��#H:�N`�J5c�wL�ACɋԓ*D'W��L����U������ՙS)�+�c�^>���{��3U�E��,��Q���s 7d�&;}[u��ڇ7M5�,���ޫ��6]��ԭq�y�]��fE�1��;�N�0�.h8�0e�f����k�.y��]�ر<*{:��6y�_;�Ls�K�����{����׶`��*m�r'd(�z}S���'�F�d���K"�N�B���+��p:��]	q�R+j����U75��	Mb�hu3M�uu��9����q��~=�"���?2&&|{򀊾.~����D��lSm�(���P����s�dT?���+%����m��om�,^,���H��y���*�=j~;�Y���
��N��V�$R9՞��XP�2�� �S.s���k��ްR��:��|f�s���,�Y6�?^ܥnC�y�OD��d�ߟ�K��03:��������E��ұ�XS����Q��҆4���9��[[�\�݅�=���.ʝ��Z��vF��Śs�������ѝR���
c�S}���L�ӐZ��Lhb�o_��LH�T�}͍��^{����l�w�(ԁ{)�ũ �b�b2������2\��է��&��=�{5a��Y�������!�1u��5P�� ��$8�V�]�:�cQ��{�nR+3�.�n\��|�(����-�4
{����)�,�U��a���2�N1��ܬ0q�Gl�X�2$,)�F�w��ڙY�ut�U��j��H�Nְ�ⓕ+���g���A�N�ɫ΂������b��5(�8�HP0d�'�5P�8��8�Gj�Ud�:s�]�-��Cy��f���������S�2��r��8{R�
�yѬ��B��s+��{�0_a�`��mwҏ��V�������2o�g�����9�i������������1Ov�'��p���0ȑ	�@���1n�w_�"�OhY�L$�.�����I_��t�N�0聯^��N��~U�
#�B/(�|z8��۝4%ފ�M�o������$>��E�5�4d���:(wt��K&V,0��Q�5�};ʀ��;~���-�U}��feWxHz=�)���p�Q�̖PΔE�}�!H��.U�*I�(ԅp(�Ó���ϡ�W7�K=�S�=��ԩc����z�eK�Jf�J�Z�VӰ����6L�s��C��wEΣ�}��W
��M���m�]#�6bb�^6�YT�~K+Z�T�<5�mQ0���v������V�[m�N𝚬(�]-�z>�1I�|���(m�M��kz��b���.��>[�r{�^:k�(��i����x�z���N�����N�4A�|mTWFm	�yV����V��^����ua&�j�,�v)��Kr�#�}ST6�&Ƕ(�N�k׏�@cõ�TU/���?g�P}���ս�V�	"G��/��v7Mq��m^���k#�,1�/�J�
7]��.wU�m�]�0����f��e����H��ݹlSS��CzK�K�ltK�\����g�1�}�E:���;���*7� �S4:� g�>�[>�4ۭ0�VB�c�p^�雊v]���Gz�ι����ƅ�D?w�R�h���w�_�M|��`�Z6%�և91&S��;�������v��3�EI�ϳ��؜f=ݽލJ/T�o(�������[�s(
�"�oOH:��֔=��Uye�ɭ�\ϳ�����V�{�лd��~����	�\F#�%b����{[��fk̙������z.
aB�`@Vg�p��]>�清���Ʈ����m�v��rcA��6A�x��6.J�n��L���Ν�̳�6!Ϟ�\F�	�Y��d>�@�b�����3��"��DBt�Q��ӓK�vۭ��ur��Ƭ~�Kw�<v٩�-��5[t>bf�4Mv���[�%Z��껭}tu\��)hZ����+W�+�H�^>J����G��<�0�V�b�{}�ݼ���Vo"�4ֵ������!򍅷�y����1����e���4��LB���������Q{�O�/�}j�.�S\�y$���N.�lF����
ƭ�-M� �sXt�M5���y�5��S[K��y������'n��n��K`�uJ�����-w�t��Z�+�t�B��)����*=�J�����]�܉��x�����(�mS绁��&>�
զHT9R���a�-Oj͉��*}��k�y$�l���r̋�2.�9M��-jz���^��a�z	鎗�F��m�K:ҹ�f߸��kw�m�Gm̆{�v]ѕL����NՅ�I�7ɾ����ў�b�$L��)+�w4"q:�gk���DV�B��a�b�t�j�{��.;���W3�%��j�����v1����Te��]��HF��% z�{0���s����Z�~�z��,
���HU��׉��Ɣ	N&Â`$�MtZ�m�e��y�]>�L��r�`�բ2nJ�ޚ=[u1�|�lk��ڬ��я���SJFŊi��ˮٻ���������q���W��'�_<�6�A�n�qS���]�YF�)@��b�^̏v���y�3Nќ��պ�������]��kL��sBݽ��@�0��N��hT�wי-��e�Xx)�:��\��4#�e�77�M�opac9�`�:��:�WՒ�JΎEՙ��ܵ!�9��X�V�ވ\fl|.���z���PI�|�:7�@s��G�J*�"�,GE�+�p	)�ح#.��*A7�;�	��-U{b�0zcg:��}�/;��!xl��^7�޴vu-;/�Ӱ�\����*,壺�b�/A�7W:�������ʐ�f���,cB�l>�6¶��5>�m�V�>�x�%x����;Ӝ�;/C�x�:�ގT#.P4��u�6Y�bi͇TA7u-wi`;pr|OXWR!��|Rⷥ�	ౖ�.�.�������Y����;����u#8n�j	]�2�k<������}�Z�.kŇ[(�%2�#R篪��u���b]��,r��X�4Z���f�W>A<��E��AW�378d̬Ui�v�M��D��-.G{��Wع�P|Oisq#c��{�a�]��rF�zF��%r������3
��v��µ�Jc�=�AR�Y�1�vvM�o�T�#N������˯"�g}�.���>�\��F��=�&�k.�.������N��I4�� M5�5V���KS��K�έ\jPz/Z7j�Ut���v���C�/1cI偨��zJ�~�TiG]�٭:�PzMJ�.ؗq��Hv�t5J��K�Kf�4�84#�Z�;�����7�Ue���{o\���T������ ���	%�1tEP�Z�뾴���L�;��O�#S���i��b�oU���5�� j�:c�̏�W[�o�&o�b�s^,�*,Tf�ሽ[��;��D������i�+w%�����ԥ�T�GuV�a$K�tﻈ9��>Or>��/1K��b��-�.��Gp�N�r9G��V	%�̌=�A+R�٪�i˭/5Z�1Z���1���4�W8"�*I���e����d�}eG�q6�=E�zdc���[���6a�onV^ݭ��UÕ�9T�V*�"%ּOb�k��IQe_Np<�vU[F��8�z���	���u��O@�N�+���C��$�mV�jh��-	/;u$�o�R��T�3�
�VP����S.Wc�A�*6q�Ȕ��^�\"�diP�����u���}KRPXK�ϵ�Y�J)k�5�S�+�]��`��Xf7u��Z�r�E����/��ؽ�\sP#3J�z$P�=%1+��Z��N��;�Ck;,M����m��Qu#u�K�}��yCv���C��ob,���p�eu��33�F84)$i����1�$2I'}�|*����뺪��k�L��&^Ha����eT5�8�U3DA�Q%D��DQ�"�8�	����
 ��8UBo2����b�4�4RD�Q�¢�d�-OfFE1A�Z�J
�b)ih �8�#�2���j(�����P���15S1QMnr
JF�
J5&Uq�5A4DEUAQ	$KUQSQPIUAF�#y�%IHU35@U%%TE�bPRPH�P�H��MP�FCM�Ɋ"*���F�����Ȥ(i")�a�f%;��B���b��+pd�1$E	He�P�+@Y�a	MU��~�� �JF���
�;�Td#3�c+7w:�2�����Gu�L$\YKU�sC��;b�{1'�2�ˠ�Su��%c�ޚYz�s��_��{�~���<��'�͂[K@e����M�S���7�YB��j%D�cnr#�s��֩Ӓ;���}�<�]��6%"�:����������!�{���^����9����W�٠����}ɵK�vE��vf�j��o�q�х���j�/��k�:�$��R�,d2���c���mk��rq��o��6�а�M�@`�����S	�d�ke1�z���	�S�u��h��Leb�'|�g�:Nz_���|ݨ��bAD+�<��܍w�P�N���{��p�.�Ł�#�U�]�Oݦ�����#����*�o�`Ifo�p�/��u*����g�c��&̇��7*����A���p)q��Z�s�P+�IÔ���8��+|1�SfCe,�b�8uI���ƪ��k�k^��Unw+�$h�:�M�7v�����u�M[�S��m�n�:�ϖ�~�e]��_�r"��6�j�p&k+������+����L�&�ѬAJ%�+4��x���]HvMp�(p�--]OkM�;�mȮ�Y>�\�"�M�3]�f�gR7]������Ϲ�J�52/��R`Bm��*Gf<ߡ.P�
֬r��ԇ�w;{Y��/R�X�#nR�g<��Wi�[ @�ѷ�Ou.ƿJ��Z�r�=U?�*�-���vo�vi�(�B�>��ɚh��?j���5t��N�R
�XP�R�r�o(�9��Y�k�޻�i��n���L���+�j���<��Sӹ�����oR��Y(������\Dt�(8"�-�hg����&��K�Y
2:̛�����,xfٟT���x��FgX;O-		���MP�8���ܛOR8���'���^�;e�M\"o`��.�ɖ!����3sѱ�hs�,�ݍVy�A�y��§��U�y{���Z�J����h�H��fŜ�ds�s��4�pV=N�!3���:�9��e�C)0ؘ`��
˜+pa�Ʊ�q�z�!��U����s��驹��V >�'`���x�}~r��D�����D&�ۺ�wR+o�-��ϧ7m D��r;�1�v�;%n�edLd�:�D\��.M�P'�Z���a�j%��y�a����N���|����o��·q�e������Av�S3W`۝/]�]͓��/��Ɔ�5ք��d�.�o8��Vӈ��/9������=������"��bpc�#<�ỸS��o�f�i����K�CY�/�K0suL���K,��6�.cE���򢆼��!+��b�R����-e��\7l3Fk=-w��\Z=�[��x/ܑ����ތ~��9+R��U�rW��M�j����V|�s_u������\uG��>�O��9��	m��ENC�a�e�2XMC��N�}�7�7��,�M5Ȃ�o�֭5Б��:Ϭ�ۖ��E�,��Sc��<�uY�7�+5�&�O��c6[��>���\���%Y}�%�)I3ݽ��7�/�6�V��!Yͨ4��u�l7�D���xY�^���S��oD5w�o��<��;oR9� ���in��5ԃ?Gn�F�?�7���M�d�dga1^�X��w����M��ۘݛ,WAv�Ȱݡ���tɡѠ��R,�&J1:;��r+qs#�{�u�3��jC;F��4��\x%��o0�t�=���;�o3���5�e�m�i^TT�;�ekb���o#YK�ۋv��W�^'�E^�f���I�Ճ�h.ղ���\\5>����&����n]���ҥ��v+�XEW�	�n���]}P���?�ie>��>{KKfa����{|�J�X�X~S0���,0����bޜ�}�-[I�\�?����pp��p��E"�!��^L�a��VF�wzrj�Fd?}o��9@��2c��x����)��1͑�9��l'�����#���#�#FCr�؋��=�=��} ����~Ê6���^�
h���۳Y���[�FH<� f������.q!��n|is���U���{}4+,���&�P�:���h�xd�*r����Q'iR8�_o���x|`��L�s�{��9F*��7ݞ|7&��KV�N1ע�,���'�Uo)kb�vq��Mv�T{��eLC|X67�1���1-0��x�<�]f�w2,۫�G|�q��$)�l�8cr��Pϐ�Wn�t74Eq~���z����b����j�u�Y���|ǉ�kJ�� �g�����@�F���͈����>�)V�.av�C�����7�r{�91�x�J����xEO�U�1����ͷ�7�ߊ�.U�4��&�zu�i��X�z���}˞�\o9A�'hP�˶�^��r��'[�{�N8_bf&Ů ��������Đz���_Ί�^No��x��_�HڏI��do�aU���	u���Z�C�}p�˵��J��U����wd"q(��bV��3e��Y���C\܆q�Xv�	q���MD�Ϻ�j(�O<�0���k&VC��t���}�C�`���/�>�(����TJQ����KN�>3�0�U��h��Z�3�z�;��<�a����S���%�wLJm�;WW���wݽ����j�fc��sڭ���ǜh�����VDNDɁ���|;u���ݐ:;r�A&|#�>�bm��q��yM�x��U���~ϐ��G�Cy��9k����i��'�R�4)sX�^�&�����<h���ڀ#�dD�z�^Gͷʳ�l����&��#i�[�9Z%�[d�6���G����*DM�������S|R����eD(a��ډ�Owqq�ڹZ�����@�5��(���z+`��[;l�W�p���r<�E�*������50��}:3aDX�����VF]y��z�;1Bx��5��-ww2�Msr]�:nKHç%7�+�+��8�'0H+i���;������x�T��xQ^�%Szk9>�xvp�v�4�nV���p*��E�����x���=(Ȩw��α'w��N}�/>n�[����0r���PoNZҪ�ջ��[-��٧��C�ڱj2˽��Ox�͒Zp��q=	e�����@7v��^FU9�pm:!��V`h7���Q��]��<װ�s˂T{��WSC:��l��l��}w��Y���>�d_(���<Q��Zvm���f6�zcه��ud����:�Ig:&Cv܇{2!�Ȏ$z5�����k<N*�)�w �z^%�����x6������؏�=E�?8��c���:�|�ۆ{�+~�(��a%�n^	���&��X��<�zC�p���T�=>�f��ߒu�&z>Tپ4���{�m=H�;<Z��:���oʂ�|$��LGD{_���thwl��R#IAȂw��O-es�ć�,���}�+h����԰������z��'>�����T�����ɒ�5�"���Я��Yf�z���T�zliݒr�l;U��NVqj7�.�eb��dRL�,Ҽ�������_?�_����	�1�"��r�}�E�֓�m��Ͳη���a8ԫr�Q7{7=|��I�_C�v�7�@Wᆼ0a�{�S�:�	�6�6�}��g�)a�;�d���l�R/e�O��1��´`�b.]h������Dhz8�_K�����%)�9�R6����x�T��n$Z��H���휢�[�k"�9��㤇�
#'Ǚd�h��R/��NKX7͏Z�4��^�v��m�͹)uо�Z���2BW7X����x�KY��d�^f{��bh�V�$���䥖(���}�����[^*���nE�������w7��}4O�ḃ��	u����՜g�kL.��'j)���OL�Y'f�����me�Y�@��M��1p4���.B�O���S>�Q��D�
��xd^W8���9�ݭ&�0ܺ�P��Ac��{�������]��*CJ��C��h:�r|~�V��)��h`�D)HK0-[rܸw���\6�[���$�=���`j��L�u���i��i+��q�l�۩e�ҥ���m�7�mr�y��Bk���:�$��9�u`�^3�+�sm�ɣy���΂n���v�u�VJݾ�ɬ�����/� ��y��tz��V.]=M����5!W=6m�V�y�Ĵ��Н�?����`/�=w�T�Y��3oy��;Z6T=l�f�Llm�U�LH7J��p�+ik̫�7B�1� �˃t͜�ڑ	�G#�[�ٓ:o�VVk�7�s��0B�����B��˽���hb���5����v���6g����=C����C�.�����%A�����$�a��fo�^+v��[�kʢ���.a�_;r�k����ׁ�2�c#��ˌ	<��/{���u��a��)�AY����'���:^Ԯ��L���Η�����y����횇s���s-�ٍ��J!HE�BT�vQ��
)�ޏf�D�ӫoR�\q�ࡋ�{�7�[�M{yLMr�:Tۀ�Z�/���Y�O�lnOh�D�nwq��!욿�]P�Z�B�Jͻv.�GQ�iE��&�C3՝X��쉪�b6�r
�̻�����k�EQM�sʵ�b2&w/joY][�;����A��8���Nni�{c�L�\j9M�'X���4�h_i������s��Q����O*��]�k�<�\��#�+�]"ܠ]�ٶf�(8(������9���� �*�X��~�<���X*QQ�Σ4�tgc�Of3����y� �Q�1J�U7�fUa�S��\.�i�ɂ�z���;q����ݬő���v����fqR����}x�Fbh|؜�jR5�W�4C��1n�D`ܑdUiM�q/���v�Yޔo*	̖�`n���33��na�ݠ!�PE�l���I*&~����-��c�ѩ���hj�ӂy��z7����-��Ʋ:<�ɪ��D��byc��Ou��<�Fo=]甌"�p�5�0-�ޟDh	=��Sv����P���X��t����ŗ�L�jn>�kK��ô^�67�5�Ɠ��]��|���w%�i��W�#�;�9ӄ���Ӡl7�R=�=�1~k�wF����J�dz�YÜO"��9� /����J�l�m�83_\�=`ӆ�ݔ�lZ)3�m��ѳ�!Y�����&����P͔k)k�ô��|'�����W��3#�7Í,��-�m����ZW��*�g>��}^�w1�mo޹JGI��xl���O>O�����[N�ꈝ�:*�EM.$o���x�u�7شd�����O��╵oCa�m�m8&�D�Ga�d>���D�]�@`����;�cI���J�n�o0��k��`�^��?�Fu�H�mL�^k&}R8�;p��C^\�r~���84�,oeeB����b�h������_��I�p�FuĻE!37-k$���nb�o;ӵ|AyR�䲶��mS�����w��\�f�K���|�
�f��|��롩}����Y^҂�]';-l��]�5�m�i/�/��a���ULE�����k�ʵT$2l������2��eo���Q-7Y	>4�A�b�pW/�χ��Vk_�߹��yԻ[��iwqY����+��2�;��os��Y�m�ȾQ����(�`�`@j�!XiK�i�޺ypP�����V7���Ř���h�!Y/��޴k�$�k��[�ھ�Iհ���w��C���pBË4�V1j;&��M4�:v�Ly�b��֠��(l]����Ֆ�P��Q̷�փ�L�&)54�Q���y��K�;A׬�P5��4o���/� �{��g�� L'oY��Ԉ���"m���F���X�}�w5B���i�r*y�0*��Ǌ�5�+J��:�O����u6^��1�(�hPc���̺�	�	J�oh�@�,����00�{e7�Tެ���.xn��rP��R����{O@9�M×2M�ٗs-eĝ��9(݂(`9L��bk�*�M�Wܖ=�\�؝?�tV^fʜ��#�q	zN��|>�OԞVkH�� ~�Ӱ�9I��Oo&�����7�2R݊[�ĴL�n34�ݬh��,�5s�*Үܦ؇[]Y���V2�2�|M��'å�]�Lݮ9�B�)?�kk���[�s��BXwۋ8�L�#T��FH���r�� �V$�c@͕��X6��M�p���'�tj�_W#ۭG�s�\����Q����.#��7�fR�f�7�6�{�_�+��4��r����u�	m�Vf� �4�N�J0!�-@/�����U�ve�P�b�1�_]�x7�����7�5� ��.��ߝuO���Z�ŵ��JyLO(�p�1�h�f2Й����_���E���!�s�s����ҶqL�Y�Fe`�MQ���w]+ˆ�o~�
�iG}�7Uque��y����ݳ�G�D����$�K��O16�ns �d� ���Ҕ�O�g(O�:ۨ:�2�A�](B�P�n,���15�L��컔��u뭼�Y�����-���,p� �4u��e��+m�(_*�l=E��3�y���Ïԫ
��oE�(Ԇ�R�%�󀕄	ʰ���;hu`��3^�f�[���人�m�T���^ۼ}E��<W(�ы��>3y�An��Ĺ�헇
ۼ�:#��[X�^�Ia��ܫ�ۍ�[׼�s;.�N"�/�^���rmG���lz�e���$��[pr��㫥<M0���<�:b��)�e,�;�7��z�N�:ƣ��e�
�~��$^rV+ �m3���D�[s~�88�֠/�:�s㷙k��i#�5`Ճ��Ⱦ��^�*.rW2��ܸ���8م"s\���>��ܰ:[�9�rV0cq�Ӧ�t�V�eIglu��a$�'J��]�
ޫ��:��ڼ��A*�����q�V�ش�*�R�8��JP]�7���H�f�ik�<��-�c��¨S�������ʐX��J��iq ��Ҡ̭#���h�D̑��N��uq����������W�1�z����&_H�26ےk�[Y@чF�f��kG������R�
���ʀ��i�b��#!��)hB7��4�SCE��MB�JUC�ƕ��(�h��@j4TT;�P��m�9-��P4��r�!
h��)E-4�4!�&���h59%U<FH�%"TEk��h���$���������$8�ʗV@j2� \��8��%L�h(
-N@Pĺ�"��ZZ�
H�"Z�2�a RjC%J� J�pr�U�+�^�o�ڶ�4�W�2�K	��H�ޭ��1�F�ޛr��ȗ�&<��Bk"0Ԭ��vD7)���k��սwR�c�	`]
�ѥBb��8Cׄ1�c1~�|:���L �9{Q�<˹ݼYf�/�U,�m�hw�i���\���f�1� aV�Cp�b=��=_nN	��ʟO�������.=XMP�ě[��.�Vtx,il�M�/��`N�MC��rn���7Mogt�cՆDFj����޻�e s^ͧ��;<Z���c�2�tOq���ϮϝT5�&��7*=��k���	����]O�gΪ�ɂ��	vXn�j��3�@����aż��3s֌�b��Z�����f�u~�i�i�P؏�a��E���U`�%����O<�������F߱웠�v�%�@*�1�Z�k}猁�x�U���'MG�<�_]W����z�{�mʿ�qxp2y�N�f�i�Cb��^��l���Cf_s;%j�&bl�_uj�r� QC�}ڈ�<����m�@��ndH���3��(e�w��;�?�X��/݂�����Ypᕆ��)Ƞs�����O���h����X��7]Z�*� 7a%��f�l����/��vf��%�;n�kq��e� }�m�[7xu�{���A�kt�%^���:���0+F>�}`�Oa7 S^��D�����wsW�Kk�Vc��rO����A�|����Q�iW꾲r�~���/�j<�2�M���XQ-'K_���>�f�uUw]J��w8�[�e���e������tk���;W����Zbw�99>OI�5��n���'��Զd)�Dh�� IJ7�5>�5�井�X.��c$U2��Z�*�U׏�P�}���i�����|���I]�|.�(WH�l}[��ΰ;�q�EP{hn�v�g�n2-�i���zW_�� ե�z���lxm�U��`ܭ�\D�ǫp�.�RƤ������Ҍ�W�_��/�`y�fZ�5@w"���uY-�LV�<���Ց��7�_��{4�Knw����o��ڎBn�k��o��x�s��O���d�=�?/^"�0���S�{T8��m��	�Wp>h#�mj�������#$M��!e9�j�鼩�(���Z�?ױ^ڞ=4���jT�CG;�-��9>t�u�[���K�jٺH�lr,;%����9�D��O@j1�-��w��r���
%Gai"�Ҥz���EՊ�}��&���ʉ]l�ǘ�3�s`����qɎ����9l��̣�->�Ӧ(�g�0����i�O�(ͧ�T�`n�
1Y�x�w _[����F�N����
jDom��q�y�Gsv�!� ڟD�����f�n)!�؄�X���-\��f����ζ���M>�>F{�Q5֯ow��<<��ǈ˛����t�I��v�t|��vZ1��8�����_	��\��N��l���=��J�[��ܩ�^�U�JIq񪃝� ��1�TJ݃��*w��Y��D��^IWuB�:�^2�wic��Y
	�mI,z���Z=,p�ǴGOt.�%"p�޻��bj�O���͢J����m�u�c�xua�u��2^V�Y�8ǂڄoit�5��&6�^^C�AS��k�=K��]�f�T4���N�R��ne4�7©�[^̜�(��v��5TڅJ�D��tϽ�×��T��2r��a���H��I��ؼ����4���Z�XQ�<3/�O�/;cGyJ4�B6ʈls3�Tr��+I�1Qnf��ٗm!)�ÏD{ӦF�O7����M$�>���� 6Ά��'ѫz��&��q�w�1��WD���w��J�+��T^�#�y"���P�sDۄ6cs}Ӳ���^���U'{z$�9'u_��m���9�~����]�� ��h�Cý=gr�6�.zT��ӓ��nO����pj�WS�Kx�Y�or���N2�\��9#_m'��6G���H�z�������gm>���N0gHsjA�ܟd���/r�a�x��8A7�3{}/Q�у}�Ce�k�Y~n/�ȋ*}r��x�Gƪ�%���h���N�i͹>�ku�4ˮ�����>��f�!��U�d�/m?�k��������Z�3�W��ϔLx=r�6�*���,ښL��R�U�����S{�)jU�v<{1[���s>�h���Z�7��{p��Y5�CT��׆�Z�j��:��O.Sz�xp����ݣ��l�n����=�)�G��[�3/:+T����
�UԮ���yYw4�v.�};��g^S��|+�Ͷ����U�R��@C:أlqZލ�V�XWN�u�.��۾�[�)k@RɁS3�F��Pv`��V����Q�M�'�k�{��Fж����u���+ɟZ�v�X�=k�=g)=\3�e��Tr�Sd�i�R�A�8񄳊��jn���DV��ͪ��ev麓��E%f��3#��}�l�
�|��#s�X��/-�S�Z̋S뺲7�dW^O���G)�k��4?���xM�`��OV(�l�ٙ�+��ӳ��.�,��#�)�Y�0[ᨲɥq9o�/��-�Y.�Z�� ��s����w{�+Fc�����bL׻��ƚ��X���4­Qb��t�aQ�ݙ��л�����jڬ&�&=5HS1)�,ɩ�a0ג�T��mΝ�u����Fc:l�ڕSVn��<u�7���#M�}z�)�hb���̥/�g��e�z����jR�l��Sd�U͍��veNu�R;��0����r�>�07�vH��/ŏצAƞ���>�Ij���{-�Ꮉbh���A��vڻ�:�J�2�C�F7?,�	��m^����ro��q���OMz���CjA|��L8\c�=d*V������v��&��,>n]]��xN�}��up�/�}-%�Rd��a���1�əWP�ES���	��7�,�[��0�#3�v�l�48��_�ƙO��d�s.�8�Gܗ�H6����r�����Ih�ny�"�e�U�@F�O�b�����-:f���g4�!�]� D��V,�'0+J���#�;.�0�ۗ�:��'���L�r�|9�]]~���Q��U��ԭ()��MFZu��:y�_\n�noe��1�k�cP��|˔��ޑy3���k�z�Z�Zߕ����w�_*Ԯ�
��V�e��M5�Muހ�.曰k�T1z�G��<?4E%���0��G���H7kyU��R2���Z3$�j*UsuV��/nǿV�=��!���q�2�m-�]y^ԣ�7v>���nƫ^��UR��юΐ}�]j���O	��>������nJF�(iE�&�mO�d�u8^X�L{�~~ɜ�IJ��dP�R�A�o>��gIF���!�u���ʷ��K����E�y;c�Iy2���E�Fvm"�����r�7��5��+�4��/f�ΓN���!YJ�`�%(}x��s���]�ɐ���\[��	[&�u��D��{�[\sM�����9-���\d\lV�U��%���%�3mm�Vi�k�h������&ɨ�i���08ksf;y�|p	����r+�'���#,�M�:޷uV��Ɩŝ���1]";�Y�MS�w�<�Y��Z�紝�tN��%��
y)c{T8�m��F.a�j(����;�%��E�R�SO���z��:b��h�x�.�2�9E3�q\Yݶ�/S��B�z��[��sI6#ڍĎT�{e@�Nd�z�_!Wwu7	mk�׏֤D��/0��@�2B-`�ȺA��Wu���桸�i�O���w3�X/E@����z��R�+;VV��Ct��(q���˙�;��9���^���O7H~�1�8�֤���<'S�jgs4�su+��ǁy����{*�X��m�i���j��7����#
1:�Y���z���g;���Է_Rڶ�u��:�� f��V��S��Ք���P_�Vs�������L�M׹�V�Z]Ð�1��&�H�YxGaBcxi���1.nn]r�ؕ��y�O��UgUѣLLn4�����&�J�y>*��:��]!����9w���fW�yQ�׺�,�g9����-�xwB�%.�K������9�9-��y����>��J�c�m��V2��v��V�i�5���r��c�]U�[���"�c2Vk�S���eHj�\����՞�-��H�/�#���5��E��Ωƣ��}�cÏZr��ͻL�̳#V�� W&��q��d�vT�_Cw4�3�ۏ>ją�J�Y�=�o4�v x���ޙqE�|��O\�GWu�Z�߉;m@�dv9#C�bAzsi�].c$�6J��3���a똃����-��{�m1�9>�V揸���D5���`�w�4(����S��ٔ����"|v�s&d�ݙz�s��XwMs�Hi�׌0i@>ّY�}�ql�v-E��N�Vu��=�_�����_�VNÌ��bd`>�[�H:�^J�K��d�����'�V�Z,\k��n���	:�d�Yc-���7�;.��p�`�]�2B'.��vXDjٺF'S�ۮ�1�P=Y���Y���")(�յ׬(y�� ���:Xn"o}9�������`4}�/�uDu����e��y�������U!��TQ,o����t�y�G��i�6˝���p��謉�}���z�j��e�1��Yqv�b�)�Z�ة��e;-�^2)b!����W�nlN��e���ښ��6�wZ;��Tt���.����}�z�u`%N��eQ����R����Cz�Ap�����^Ue���/�v�NC���*��nW��d�Q7�r6x�0�RRT�6�G�\I�Qn{vx�K������??t8��>�6�8疹img����u����� e8{��#8��Y#.���N;�W wvd��g�S@~$V���L�0Y�G�Bp��>-�����?�����ճ��s�^����k�y`�q1�a��w;4�uΫ׼]�������*ߩ�%l�6����z�W�(��T�N�k��>R�sf�{�p$�b��q�!�G��53���IL��+����`�G�4� |��Y��Օ�n��XxiK����k.�p�v�5�]�e��K�'(�V��曬59��Y��3��k�G���*��k ����T[�y��7��p�S���)̀����ڐ�X{�.U.����s���O#�LF�^�����P���wJ����W*ή|���t��A錯	7�m����3�Ab�Fِ.T�;\��:��j/"[g���aۜ��ޮ̹闻@���G�]���Xg�i_+#`e��wl���lߍ���S�=�ru)$��U���ՙ�̔��=H�'�A��?/���*�+ô�o[��[%I�$9�S�ؘ��wW( ~z���FO�>�eT�噒���PLFexU�@F�=��Z٪�W�r�ix�k
�Y/w5�Y���*MxY@���HJ)�C�G_c��l1��Ͼ�dB�g�t��zvFg�]K%�h���K/P*&j�7zu�{���3��U�Y5=�*�e6IM�@{�m��&B��[�z@�  ����=t��f!��w��E�#�Q�Z��u��u�l\D�z��\�6��*1��4�,����g��q;��9t*�v �32�3�|^ngB�9�,�Z�����e.	�k7f=0>+nP�{M����6�٦��66V(3ꗜ���])����+l�1�/f-(��-�f�m�cj'2[��w�ف)V����f�Ö�ll�˨Q
��]��`�*�ޭzʥ�f�G�v`���ܷ����o|��U��`�
ݨK�I��1ݹ��:S/OaK:=����m"��J���V�ǥ��>ը���đV4rK2��f29Æ��,u�u�40֋��-�8d�M�CA�ܥ!N1�[�f���-Hh�aM���훿|m�Nmp�%>ͅC���j8�qfpA��AoYNv����}�P�� n��c���󻡴z�\�8eK���rjb�F�K��W�c���b�᧥<�8�r5���&��y�g��Zi�n�2���m���U��.�Q�����/�Z8r��[q���Y��咹<{pM�|���8	Ū��6��-c%�U:��c��7�r�Cx�����񉾃e�ze��F����5(:Z�w=�	g�;;���x1c9ԖX�y,ϫ�r���cyЧ$�2;4Zү�.�W�fb�� ��N��Kr\��eCG̥�r���y´�R�A̱-�Tn?��#�3�ӕ��;��<�8.�k"��Pˢ2�׉�JyyuI��9�����Uפ�� ���\��4����e_`G�m\sH�S_�6t��%�v\�t������`ǥn���u}��t�,I�W�����Ю��F�5�1Z-�^5�k��u����7�����Y��̧��ɗ�H�L�m²�=����������x����U�乹q��� ��p5/]oX�ܸ�}�{Rї�k'u��� a���0e��F�V�k%k�he
,�Ǵ"�Ik�66�%��Մ"��k�eWe�j�Ż�U�ܭo����r�H�[�� "/]r+���mi�ҟ(�pLh��Y�FѧE��h��ѹ���܃y�.�<`�;c��Sa�{����ַ� S����}FE{>)�j�96-R�������E�QV[��u2˛͹����(9WF��*�;��#�/7*^��|��=���h����F�uB�z��"����ʴqǪ�����%h`Y���z��>�����9�����V�����[��ka���܊�Zxů\����X���#�
e���@� f��sb��8'uB��3C�U��.T�����x/���v2�b�f��%%%n響��n��\���G��]9|~f��:D�����;�F�y��[���u�z2��0��ł,	aA�N�]���{U�m�p�H��Wy���r�w-c�ݳV�w[::Guj�`8���L�%��	�{;�nJI$�N���ITR@���Z�)�M�Ԧ�
"i*�)�(�(5 �� �F����-X�%4�RP҅#M<NJ1�nGR4PPQIB;�rB�f+H<Y4��CO���-EH4H�R�:�%�9y�2��C�P��Uȡ��p���(h{�	@�B�d�QÓY�w��2(�����K�.H�\�PR�!���ox`����A��陷�wݕa����`�܅'R��v�Y�̾n�:+7�$�y!d��Wq���;j���f!�͖������]ά.$���=Go�?Nϒ�� �xl�X��Mr ����w�2^v�F��"lix�>c��K����t�G+|�ِك'rH�h��,�ɚ��G�<2����@�`�!���Kcʺ�G6󻮤�i�ah�^*;������fJ����ܨ��^.������]o�յ�,���{Ș!ջG����s��\d��Jr���t�s=�9��5F����笭	�e�7 ;%���s�s�"#{c)��_�^��>�g�E��N-c33���{���t��So{{�����FȜ�e#~�Rpp��o�X�ze���+�HO�'���<��Q��2;ڠ8�����M���'�=Q��%�ZK���A;`vKGv^3do�0��z�Xwg����n@נ���
ˎ6(R2/N����Z}��2Pcv˦5�7N[Xc@���f�կf�y9�1�h}�8���q�r��ի�8��(y��:�(�g
6�K��nn,N�ai���W��Ҳ;��K����'X6��Wy��U�[E��#�F5b�ˌ���6z,��В��9Xy-w�ټ�Z9&|(ՈWv������-��_x�?�y�::_\5����&�V|��7�t��Lӥ��R�&G\v3�a��� ��.��5�߆�����=�N�^e-���@���34��:׆�!�xr/K��t�;W�!���٩���1��o��C��m�3Y�{�#)%Ǥ[�׏d#S�wb�|-��<�lѥ�,p77��9�|v�+6&{+�J��Y�����:�[��Ll�r�eq{&;#o�Z9!{�@�FO����i�q�hs�����WuB3�sF�:��Xl�}�>�ʆe���L%�,��Zk�#l��)�/G�k-�6�c{�5���uⳙE���igq.9,���E�eڀ��ʮ���I@dJ���Y!,��\�X�2�k�4|�H+ %�"<��6�p�)��oK�?����+8=S��UWw�P���F+m�����B�i�4E7�z��Pe��mSN�iY̪c)��4��^~s%��B�+A,����j��*}�gL��1!X�߲�w] 5�uf��c��[%.�k���]�M����a�ﭪ�����]�/VEt�.��������h���Ü]�޹l,����᣷��#��;��-�y����U��Myf��:�^���G$hy
�M��}/qn4���w��޸L%�0�����ܭg$^�+iތ��n^]�<)�m+���hT�lG+��.Ll,��d��>'�U��l\��K�58��C7��yQ����|o���ȽZ�2z�lz�~�nf����Ph.�����z}�M��*�Z"ט֙�G�~��W9���b8�ie=�=�j��|�f��~����xi����TE�%�7R1@�6Qk�����2�l��x��5���_ic*u	N]����Η�n�]�Tϫ��J[I\�.ǋT�UK��[���[_iܦ���6uHs�A9Sq�;�f�`�yQƸ��:��sT�u��0cK�{G���j����}~�׵�q���9����w3��z:�,���zHO{40���R��$���^�؛g�b���=�kZ�̫Mׇm�7����3+� -��l��Yy�M��$��@��R��y�7��Z8 �|�8�MVhu;zky�}s����ܙˣ��/���ܜY?�U[��n�}^��]t�d�������`|2�Q�np_r��U���֙k��ܬsL/ݘ�nV�䑥�a*٥y�Ujw��S@~��~�;�]�n�̶�Y�����:�W���M1EPc=��]�
Y��E��� �V��'���2���{��꥕������N�W)��|�%[�x�3n+2��"߉jlP�t���x:����s� V����=eA��r�Q�1�ٟ%��*��{$�z+����2��C˄[��Oߏ�����q	Hk˯_{ 2��r�9O7/0��}l����ݳ����Ɲ&���.��"���O`�5�sdz䞠�'��-�w>#���.ٖ!�fv�#[��4c�%�lM)�Kt�S��� @���Y�{Y2�M^F#m��������=ym�X������,�!�W2"�ZcU3u�l�ɚ9�س5�����O�g�_z�Y�]=̜�82�N��B�U,���$P���d8�O"��ɢ̢o~y�;�g13<;�E ^|g^cz��&�:��Fip�,��
^�u�)��z+������dޱ��s&gL�#Ɩ��UV;\o���^����";蛿�r��h+���W?wx�����/T����&�ȫУ �Od�Yk:�nr�c�I�t�xcD�x-�N����T~~#�`��+�oM��+�³�Q4��Ql36��v�>�3��-���C���
�)S�L����5�W*�dVU�N����n ���b���u�7�uz̜�*��Y�E[�^2��%��s$�*�Ǽ��x{�h��Y�Q���	�k4U���+Ȑwh���iv��8��S\΋7D�KE����۾[�u.��
f��~ ��]�%�ϱT��o�l2x��}/�%1�1�F�uU����t.<���J(�Ѩ���Q��<�6UMf]pt�쌠���\W�d�_Z���/��J��b����m�w�}^AD�a�+2o��@� z܎��~[�3�1�_��ԬV�={�1�����^N]9�Ճu�'c�S��=Z�-�jg�5w��a|%vv�\P�+Y�	7�B���L��\Tu��t�{�	n�M]y��h��&�`��Y C_ll���ݸ��j��bn�J>�ݧ��Y�]]_�����]�N�X�߂:�j�t|�v�qΐ֦��oC�m��7У2X�	�?<�4�x�u�l���=ڰ�Wֹ�
zR�3�w�0��k��Q7���p�D�N�VK
�et�D�r��p��w���6g�h2�N�x��5O��p�11.'K��Du��1��f#C��-Űb�Vb�TOv�w1�7�;�(��O��V���Zx��i��R�}��놿b��2<�}ܷp�S��hI�k�������!�c�f<���&��2֢z=;��Y���Tt,֞�����#�d{J��ݱnv�~s��U[⫖T���D�4�g���1����P�b�e�jn�;��b�x-�j�[�7.歖+8]n���
�Ԗ�n7ä^���ڗW�IV��wUgH6�N�!1�R�0][��o��ׇ��@G$G&ɲ+V����t.�%"qNRCT�a����&=t�;�1��dn�f� *.�VS�� )�y���Ԇ^jy��"*,W��9����uoR���t�w�N�k��g�N[�R+�k��u�vn�}J�iʸ��ss�-��� "��8h��fs�ko��/����9�Qcn�P��v��<�5���z*k���⭿Ny� ?sd�Kd!��<�@gv��c��	�
ᮬכt���{_'2���}D�Ѓw:*�@!�>�dXY6��e��<o4e��^�έ�&�vM�r7;��I�Ż>D�u���;%d%�0���Ꝼ���'�	���?Q�^�g�އRWrV��s�V�$o����Q�ڇ.�y����D�w���V�7`��ߧ�ue���\��>���
ɼkE�\m�!�� 4��ʺb9LB�����(%�r����_(�9,�*��^�jT��{:G�Ĥ@��*ܧ�ݟz���	��0xx��|"���{�t�w�Yo(7O�S:�l3��d@Vg���{qi��{7z��Y���h㪚C�����)R��C@�k�~���,3T�غeon-̪�����;�dgS��g$'9><�#�&����v˽�M����X�Q�ܟ~�R�o��.V�84����0�N۲�R����JD��Ǧ׵�:~�����E-�mG���=wx*?~��,�Qv+TA^n���b|��$��=8�,��Y^��a�f��Ҽ�ƙ���k5���N�c�iP�	kI�K'QޝkGS2�}9��D\x����LqHl���L�z�N�aAT��-�g;�2�4۶�$5L����l�69DW!� �w�Z��a���j)��<�!�������R��h���\�S]a<��sx9
PnfnkwY�y�0w$��N+E^Vm���*�7Q��rl�i�R�A�8�Uvf��4(r����p�d혮5K�\/^2�υσ�[|;���ca.��M�)���D�
�F��=iQ�u&.��޷��௷$|35T�؟�2�m�7ZwOl0�"�,2׼Q�ܸ�c�ڱwAJ���n��"46�T�ɤ���
ס�-�2��������ʁ�������cߒN�2�)
��M��P�fa�LBީ���UV�g��4�g�B�
tzude�(�y���A���fX[�?D>��e�M�Vgu�,�T�d���;[#��R*dЩ�wƭ3�\ؘ�L=ɏn�w�cq'�:��!m,_f����W˙�B�'܄�v2��=��a+0��cq�GF�#9�C�E��z7��.̨��e!����J� e�&��Q�\�J�ei�e��U�a���W#w%#}Q��cU�h�ϭ���w�g��븚1x�p;�Qʻ����Pb������c"�A�{m���.�1EN��	�ͷJ���݌-�OW��r�go7}����J7!t�����O�X]����U�K���'B�����/cَC�/�0�ibz���i����D�i�3����Q��ψ�x�P�G��Y������hE�<�.Qʕ/��QMw5������t�#Fta�S�,����:���(����� �etwӪt�k|�58~H�<t���ة��<��TK�����ʶ��-���eM�h䅩[E\�y+��N����0n���ȅ9�����i�7U:��Y�ݨoL��]��3Ƭ���Y�E[�[-�0O\��j�i���L[���/�}DNQ���a�6�@$���T��:���Q
*�A������A��#]%g��&��l��A���n�K�4���v����� ���9�R��(Y�g��8e����m%kN�-�C�l��w*�%��J��qw[n��rfh�J��p����1�V0��:�VE��R�b9C:�:�Ŏ��\��ЩΏ?����[�}�p�s;�e��q��jw:%��[�&#Lm(���`7_-�1���: T�yغ�˹Xm��fʛ[�csz��?���mOx�>v���,�e�!q�q�+R�
��u���[��	���;9��;�����M���z��"7��]��4˕�^����T���*̺s��M�����h����ʢE�=��i�.�C%G���	��"�!L�T�{R���%>���������>i����ki$�� ����M n�oU�1n�ϯe�}Y�n�pdX+�\����	@�
��FF����	�*4_	\��ʽeP��ѷ^�_R��(=.�Du���X3*���oh�6-�9m��xٜ/kB��gKX�4#e�Þx��+������7����0䪢���@D~���T_�
���Mc��q'&�b��҃� ��0t�	 	@ 	@	 P	@� lv ���Qp% $! @!!P$7`0J�J�A� � A  A  A  A A" A  A��4� �   ��@�B�H j�@ 	 	EX! $ $ $ $  U`�h6l0 	X U`�  �  �  �  �  �!X7&
�
��
�(H�J�J�H�B�f�4�++++�#+++� �`����s��}I�7��DE �D�T(��v����{u�>	�����}���������}����Om�cd�<���?������EQEv��O����?y��
"���`�����_ڿzpBjL!~�W��pS�����������ߵ3�� ��!{�������c���3��>	�X׳��4��
Ĩ��H �   R  @#  D�0�� � B�J��H ��� (� �( B�����  $���"a��1�����آ�o��Ȉ�� � � � �iE=�����w����$�����8�O���z�{�@��+����|ߣ��}~�o�O��O��z��UE�}
}��~C�~C�
���"����>�_�=�>z?Ր^v� 5�@zS��c���^ �~�4�v?�3��D�xM	�6*���O�?%?/���*����x?�;���|>����>)��=�����'�qUE��zg���� HH�J��-(�@�҂� �(#B҂4"�
#J�)H�Т�
�(�H�(
B��*�*�(+B�Ҫ��-(H
҂� � 4�-( R(�"-�P��*#H��J �� �H���J����P(���P(�J��!B�H
R"(�(Э*�	H��P-"�-" P� �J� � �B4#J4% ҩJ4*R�{��E8QI3�Ҙ��RK�~BX���I��Y�|~��{�!��zyEQEyK������������rw��_Hv���zBEC���IƐ_}�O^���LS��������e5��*+ �]�!�?���}������⪥B���R"T�J��(�*J U �$�@�Ji��$�Lm��ET��Z��*�Z�P�b�*�RJ�HD��HP���Q0���I*�R�E*��Sw:�E�pJ[(�cJ�٪��hU��Y�J��֊Fm��
UI��4j0��P� IcEP���@SfJ@E*Qe�
������m�*
�1Eh͚5�
-�H�1IB�k&̒�p�e�T)��kF&�2K-PBk--�-�MIE
�[��G!��-4 Q#A��*S �U�2�ЫVP5��l\ ,]��E��i�e�2� �ʦ��֊(�HET��R�� �R
Q .�B��m� �
DT ـeV�)+l�n @ � � b �  k @ ��iQ��\ n  L 0 &� H h��h� �� #AU���� N � m 	� &�� l� � ` ي p     �~@i)J�bhɁ4i�40 �S�	)H� @  h  昙2h�`��` ���S�A)U@  �    9�&L�0�&&��!�0# �I&�L �����z�Q�3����{_O_�^ϫ�9��O��]����:��I	;O�I!'���,�j$�$=� $��D�BI	5 7����O�����h�	���$	 l��< @$��:�?���I	<C �h���T�YI!'(�N=w�{_��|>^���BN����Hx�d:|3�^���\���n)A{����^W31��q�����m��@�u�������[{e@-��u2�V7i�-еF�Y6����ͫT���y��`ڄ���>��Ѳ��kdd��V�RR�.��+�V���bgCX*�M9y�'�Nǌ�,��N�G\�V�l��o5���&eZ�SS����X��Y�&�r���Ov<�nQj�H�j{�Sj�x�F�v�5sPx�@�e(��^ ݫY@��Q^2�_E���Eh;��#fS,���f�u�eC���wJ*k��طf���.��M���\f4��i��Fh�HVE�&��ݤ"9RmŘ2ea�wN�4�7-w�3�"
�3P��9���.f�jJF��jK�6��BbF賲�HYL���&���l������R,��b����a�6��[B�� ���N�T�(<��zv70���1�%E'�KI �@�v]�����$ɋ0}e��Ȳ��Q[1"
P�R�G.� �X�e\J
�h�)��4](���v�"��CQfm�-�P�aR�j%l=v��(I�u`�n�ۛLY�
��ʴ��z�H��Iin�t�wIJ,C��xl�͡~U�ʣO,Z���bM]I���j�������,2]�:+3mm%��Ie������A�V�f�vn���/>(�Ch�t�N�{��E��]['K�B����v`��M�[�_K�Z���
�]CGBҦn�j@r3W�f	�[��.�ۏj\{ �#�VԦ�e������^������J��[�bߝ�6e�Q�ډZ#��GJ��3@Њ��7z݊%�������9�N�A���Yf��5�gKn��ww��2��`��&��ڰ�GN�J�x��e<�[��j�(S#]Ǝ;R�r�&f0Y�����5H�`Z��`�b̛����a֒Mk5����V�j���Wh�oX�`�ڵ�Z�ǉ���I��U�u`K�
��:�)��A�c�L�ji���hZ�v�m陻V���[H��,��G&m4��s3P��GN�\xe��U/j�qT;�Fq��;j���͢1b�W�L�j�Z��ܗE�.F��J�E�nQc��h�� �2�ʚ�6�!aV�42��wf桫@06��/1^����[;Q����!!a�N�YA�[soh�v0<(�B��`�	��,�m��㺶Z�
���}��zn��i���*��BE���SQzC�H,k9�'/7,3K3��G�ř)�(�;���ج�-��%�h�;��X%Ұ����l�r�[&#������KV��e�z�U��2�e�mU�uzK"����V�BM����s/+V,��fYT�1�%�1|�"�m�P�2�d���g3H�m�Z��he�mE����dt-�8�6�`��Ee<Y��&�)�h`�7C�+f^Ö B� v�n�L[�!�q��[4�S5�ֽa��Ӛ���噢���h`�� �r�%����5��F�E�sU��x�]4�	mŭP�A�����)սZ�pm�9o3j�
��4r-uŉ%kQ����hmf�Uƞ� M�
��n��kH;[�N�)�%\�1����M��n ��wv/a j²�%� ��-'�#yv�j���M7C$xSj���fZT%"ضAo Q+���:�&��0~8�G��u5���l��R��`�����i�5nۙV�8\�F����L%d[ l튃#��b��mQ��X$n����#�`B�l<�W�q4�<|��.2�&VJRٔ�����a�j�0�bv/5��%-UP;T��B�^
50�z��T�T(T�b��<KD�GqJ�#�J�¬F�e�Ss	cS�ț{J�؇v�\Vf�T@�M���M�Ux�:��ؚ5�Q[����(�6b��;�7^���<Ff,�:�T�nN�Ԛ�Z���v2���dj�� ho��A\�����5G�I��hR�f)�k��S��;aB`5�H�P�B]/@X���e]�jm8�"[-�[�4N&"gpn0��ִ�G�H�^�B��/(�T�0V�@;�[f�24��/�l3�����n��Vd� ��#i]#�����dE2�&MJ ��2;0k6��X�j�2��;�e�7)��@���@p�wfU+ۃ-��p*��Gj�+���boC�{��6wրn��u!��H0C�[$6���̊�� �J�Hsi\��OYMG�w�ЗW�R��4�L�5bo5��.�wu?��h��ۛ�p����g�$�1�kh'�a����>�Z[a	�� w[��l*�Iէ�T/a��t�6+(����^�de�����X3�U�N� ��V���+���JYӠ=�
4F�U��Zq%�\͋p`��Gx/"*�!�e�	�dt�!M8�V���m�9����P����k\� ����JRDf�q0I��f
���|�X���-�p*B�hk�4�"љh�1A�E��������tX�ǆb;�l�S!��q��o
ӿ�i�,@�A�{�ثz&� 5�]H1��f��f$V-ç,ҸZ�bWA՘I²;"�ލ��j�Pʆ�
�i�/p�m�ժ���B�Ӛ��M��ٳ4ռ������;%aw�U*�y64��Q6s1T�mns氩Bee�t��A�>i�p��j+�ol�YyAJvt�W�l�	ج�]���`ah�	�1�5�lk8�!
J��;ɑW�.�S�f��c�8�f��F'J�S6�[GDu�LB��-z͢� ]m�T�n�Ub�c�2]L���s!yt�؋n�8謸�z���4�B�r�l�OĻ.�˶�Gt��j���d�V��7{�UY"�ue�%Ɲ[أS6�O*�,H�ٌGlK�A�1b�,�,�݉�-� D+3n	�HL��J{RQ�W��Z�D��s`�J��Y��6*�ږ�%�j�2�67h-M��kD�o,F�݆�pb��XUg���n-�``#�S0�$Y��d4 6��J�6�楷=��bkF�c@TUn���GTGj0�Bx �2���<@dZ������>&�D;�[Bi���(�T1
t����K��-]=t��Ȭk�A��fe��a7LW�P�&Xn�����J�MQ6[��0MyV�{�-�K�ȫ�r�*�d8,&Ͱ�"e�h7�X�VZ��-b���6�e�Z��6���iӦ5���\z��j��ʼWB� T�h���Z4�p��68��xSjwHj$(��e�(~�nV�%��C	ͽ�F�*KJ;0��R���vn��0�S��4m�J��:��7x��j۪yh�W���;��/ߪ������@>~��h:hÂ &��on������=GJ4���¥+��;÷b꣋,��Ӑ�4��٘p��y�b��`��go^h�@�j5s��9�s����[���.�i�Ʉ��������
�1a�^�
�q:F0o��OMT�{>N0���rv�^��,|��r�޲æ��9���t�q]�J�Kj,�ˆ���<�tr�Y
=�}X7WW�u�7xW:�G�ɑ�0z��N��wd`�\��0�|���3�c�	K��3ܗY�Z
��[�^A��t��:U��:��f�nQ�r��Sո�|;k����[�C��8���>[Z�;�l�TY���.�q ��d:�	]]5�f��{vhm(�L]�Z�Ws��H,H����*�W��VكS#vF��!n�����hҵӆ�C
�g

�\#׺Ѭ��51�t�2��DtK5`���L�����F�����[��%��f�+����m-{��Y	Ú�jɾ���X�KB�*���Ď��4��O�qy�k���ZV��?�]��:S-d�q�h�ņ������8����9J���1o��(-�9����Y�MJ�˵Y����;��c2s�C�gt����[Κ�S-8~�B�K왺o�����b	N�p��}ѬAuӹJ�m.Qζ���E.7<:��ن�L�e�n�o�^l�Jq]fl �R�t�5-��'�r��z8k��孌n���!���C�L�lc�.+-)v�1�ִ��X����{s&u*���6nK�������+j�}Kv��݋x3A$]��U5
'Uك��AD�^�0o�X�h�71��J�VӰ�:��X��˽+�H�* �� ��'�^S��u;�|S	C�"��u���TF��p蒁CP��fK�=��q����gV�b�|�F�P��h�Sᙕe��t�y�f��X�he;L�����s}�-E5v�w�5}aj,cض�s����$c�Ar�Y�3��{KO]M�E]9��n�&����;�* ]�%�yp	�G�(�n/��W����A�O��E��tdP�7�����8m�7��L�cM��������8,��z�����j-D�Jm�K�o*l�m*�E�L\������%Jc�`>�[A�[���s߅p6h�����ƷE�H�u�b�[K3U�k����7�a.���AHB� U���ZJ۔%�&j�E܊���d^Y��LzD(�8lJ���G�&@�6�K�T�
�9�7֙���j�L6�� �ka:��㔫 G�YҪ��J>�
<�ޙ��`J�/d��a���ۥ{L; ������wx�����B9�}Zi<��	����fq�z^�[����D�ND��,.����c�ʚ&X��2�B5�*ͩ�X�#/��52+�;�mglԻa.���c؆��U*ú��<����묛�#GX/�����Ѫ����:u#;��$ȷ�m�����,y�s,�u��b�km.�"ԕ��s-U�N���ыU�N��u�a�u�\����mÂ
����Y{�(3&(ޫI���:`S:mIuJ�sP��[��urT��h�Z7�A��H6��+z<U՝����l����c[��mr\��r�p�B]t��KJ|�*���@ecZmK���w,�o/��-���͚���;�K���ۖ($�����ؕ*�$���ذH��rjs�"��ãH��ܜ-'E5����aMd�P1���Ѫ	�V>���C���������w�:.�u�_g��F�Q!��q��Х�3�b���H ��=6-�{��JH�V����>ѧ�#����}�N�w��"�oJ�o`f
;#��BRI�N�PK:�Ž�R��#�Q�,��\#�R��΢�]j�#6�*z�ې�m�y�]ʈPZ�|]���+2<Z 2��z3K�2$��n�Ŭ�RC �����X�FR_v�}cF��U2��7k#͢�N��2g]��J՜�\
:6�7$D���)�oi����`��ӌ��(�VkN��e0a��0V�$Ĝ��Y�R�mN��e��yz�ާt��ȏf.�ᩴ$`���f]�m�ŃoY�`"������8�v��]�\���S
22Ěe��w��%�9b`Q� ��;d:��&��t��i�����W�,�7��)�°�&N�T���
��x��`H�{V�@���9��e[�qHD�E�>#/zD�5�#�Z�P� �
�IZ�V�]�2��I�&��mwT_$�˕c:z,N���@J��a��*��	궋·l���H9�L��jc��Ip��Vc�q�R=t�6s�B���zF�j�a' ��h�(�Y8���;*��(=�9�B���W\�F`{���h")�w03)D殲2ge����,��-
�oq&0SNu'-P2ۈzj�q.�=���Q.�M�ⳅ�+\� Nb�6��|�_l���P��5`Ds������Ѽ����W����%\�ѹ������R���Q�> >Z��Z2���#v��iL�P�� �y�PU����t-�b�bg�b�L�.Jqc��&'$�Ზ��zv�r�Oi�M������j��dsb�T��l��쨷�s��w�'L��RˮD��t�Z�a.,&J����	Wz����oP����)��p��Tk^��{R�˂j�|�l=U���3�*�Y�Y�x·��ޝ�w�w�*�r[DO�����-���$Puj��tx�***����wz"��єo��a��ef.=���զ9�`5v2l���W`�LP��,�W�I�w���L�����K��n�\@WPm�݂���HD졲�M4��3)� ���G��5�qh�������=�d���
�z;�;:�)�P��ɗ�J���Uw)e-�Pc���T��B�/�N|�*�ӎ������(�� �ֻ]ד9T��c�����]E5y�%��o���5w�AE��y4�6	,�8�-��:�[Y%HE��ó5�.땆_%y���r��������U�Y�G6��դ �^\yc���K�=;3��s� ����w$�]Zs:�&�:������m�ڵ������m��m��m��m��m��mC�x�*2���ݷY�ӥ�6��K�w�4����������í����5��m��m��v�sApխm�����m��m��m��m�Ͷ�o�m��m��m��m��m��m��y�5����ӻ��Sla6�	N�ۆ�Z�Q�=]�%*b�6�D���m������m��s����{�Z4�I��â��:�'ӫ��8��*�.\�^F�N��Od6�i��[c*^6ιzݱ!)�W��f�8M���)������J'��>��6�hbN��=�sN5bn�oom�c����W��T�����?�$��˴�f��$$	'�<`�T�;�'��DI	=��gY��w��l߳�xo\o|���8מ8u�I��X��(��6I#��Zg�ަJ;�Av�t�H�WX����\�^!S>u�(�o\�:N	ZxݽV��Һq!��u�z�T����v>���YrK�p)ci�q��ׅY����t��X�� �9�:��"��:�[�	�"'���Ϸ�pO�}���Z1��ǲ����͏��� Z�)Ǵ��Vw	��n3q�Mz�NH�ųG@h�����^j����IC�ư�'�Y{¶;�9vy��WCl�]ԸR�qgwh�Rvh�� 9�"���6���L��SSL���|���n�X&�,LE�%��/K����ׇ7�2�f�T]��L�܏D�&��e�wY�F��!��_M� ]lᝎ,�ӝ�M�	)Y����9�{O>��]�TJݺԺ���-0J]o�-5e����5hڥ�G�Q�83��ܙ�!G�YO���˕��
C�Q����C&t�b�V,ʲ�Pd�y���������o�.q$2��r���D�ʎ�ۓ34�'{í&����}m�M3�xNsWW�ԀqU����{in��Ho\�{\#P�yKn���@c�v��VP��6��Mui0ٲ�w<�n<�jRˀ�jUṝ�pRu�6�'P�<�t���E�5��y����L��U������c��W/C����i	&0ZD�,TL��x�^k��4VR��� ��k�%Mi�Ffٻ�1��25w*��WK�5+�,���q���;�N�'y�tqţ���c��<FIٻ�򣽼if���B��D���f�-g|�J�Kn� Z$��uEu:��Z�F�t�׎���B�-a�V���$�\��/��bהGf
3��U�����f��QX{�������?f+��u�g�!ޔ�]��Ø㒙�����R�,�ԍIٷB��[�Vf� U�ˀ�:7��P��I+�`�����$�t��7�mm}��9��إ��敆��}��n��ݢ��o]�R!�b��k"�[���9��@�lw����TV
��r�#2�n�2�T���j�'uy��]�]qE��]������������|��pn�)�:�!�M����S�ɑ�%���m��)Z��&sˌӧ��u��(N�l'�
wM����$�j>cN=vSZx�^�o�5�r���Y���Wyɝ�Z���[9*��ę�F���Xn�2����e9w���,٣�27'v=�1tK%���\�j���P�*	*��;FEH-v`Ơ�m�p�J�w7��Cq�ZwG�^��*���r�ي�Ӳ��ٽ}{A�5��NR�U���J�aC,Er�����"�r��)�H� ���0��rkXR�ڜy�f�X��ٮ�]Ck��,�+����6��$�Ճc��P����t�Pu34v�r*m���Uq=o|q;�Vý�o�>���ʵ�oכ�;9��9��ŕ�XWQ�c�+F�����XՐ)��o]���P�h��t��qL8v���&�l�U���]X�׷#f[V�Fy��Bѣ[��#.ѫf�
�\�0)��r�� �yw@n�H<-$����[��+:�J+mg�x��i�/�g")$���k/�!v�!h�ǹ(OAAX��Gv���6��7�K/�g~q3�,�L�5�sM��Q"�Q	�~{@��<t�P��s��2�B����Tfr`.��X����s��F-�0��&�ކ�)��2�_l�ne��n�ԁJ�/�ݼhB)l��8���I1g-;��?�	�O�&�Z��S����m���L��;s��i]e�:jebg��%(�=���e���VuG�H�G\X�>ŰWTu�J}��������pI��y�H�Xo3�f[e IC�)\�m��1Dd����<��Xn\����ӈr�pu�[I$k,��/hqwx���u�U IdU�.�����+��/��@P':R�z���7c��[�I{��n����J��=����h��M�:ɓ�z6�+-8�:�<�t��Z�K9���h�ٝ��٬�����uԀ�+�Ǽ*�����V�G�1�o.�r���մf���V�U�t�֊�p*���S�0���Z~Wǔ�+0��2v�!5��c��X-���5mi�4�!� /stwK4���m!�X�r��8a9��N��;Y��t+&Q���>	X:�@���:�QZ�D	y�r�l��k8Q[�AP���O<0Ýnl�o@q���	�t�B��G��m�r����:�H(U�h]j�bg%'P�)��jwu]umW�j}�Ʊz�w�l_,�^�'�6�Z���pZ��z����^�F�`R��ZF���J�����Mn�-�'���<o�|v��nă8�ήk�Ag����5�or���[,�+�Wu�i� Sb��|�4���U���G	Su���f]QĶ����z�:�]7}:�ݒ��.r`mmZ1�9�X�Դ|n��m96|�T���dm�
���$K��
��9���y*�	��M˓���*j�n�*�:2�Ϟd<XHԫ!��0��C���K�	�V�<����k{3a��]=�	��A����>u7M>�>�3	R���D��{6��%�o0WZ����l/i.���O��.1���ܙ�qJ�s/�T�,��g&ʧĸi�7��&ۚ��.�[��+��|։�F�$��q�3��S.��m�(�6��m��Ri#,�1���ɣ�+'D�3n�8;*�S��fBdj�/H�d`K4R8��Ju,�Syl�:W�B2P��DV�&��j|�� 
��n@��T�u+�s�X;�3a���)����Հ��ev_T��2v���pD�wj�rA8Y�]�6�M��&��� �x�D^�BA��OG�/4(���y����f��p�I���)cu!o�.z�^�J&�Zi#]�]0H��]C��v��t�ͺ���5��㰵��@u��|�
w�{V�W)�ІT���a����\L��ST�޳R�]�7�ch#���r#�V*nH��fޗX-Z]�+����O�BuC6<��
!�}�dd��V��r�9g�'.wPp��(G3��B��W����a�p+�4!����>����,��T�6��d#N�l��Ô(�hFl�\��E�O�m�M��uWT�V,�Y2FmT��d1a�JS�
+'M����;��;cgBNq�n��tЗL�6i��o95�{��}`^u�M���=9��a&Z���Lɧb��-��zN"�B�V�G�X�߁��b�t�g���-\41�P��͘6��q`�`ek�6(�1-��f��X�:hhY=��o\�x�)t7+
��k+ƭ�XF�i�[�|?��|>���A���,��!�Χ�k��]�z-u�լ���`�*Jp�#�n�/�����J�h�h���2X�$�I��a��OV��X�&�Nq�����AN,���)+B��,�c_Y��v8O#(�Գ�:��B��s��5Je��!e#��M�BRg�[+2N�gM�P�n5:vc�sw�k��p��D�5)��%�責Dc5�W9y�C�f�Q䭰̦uc��*�P��)/�y�)�hV��&C�Q�����J^��-��wK�Ec
����2�U�[�L�}Db]Fو�9����S��v�+�w4���vv�f�����|����}�TX��0�@��̥aXuC���(�V�XŊvBc8�:�p�I�J�11M*HcSHyI1:�`m�`n�*L�ta�{l��$6��*:&���ʺf����6�l:0��m��'�"��I�d�E���hm8d1�AVG)
��ݜ��5M�N2�IPĕ���H�DY
Ɏ�u��{\x����r�Td|*u �q�n�o�Uwu����-L˼�������UF����T���FBv�4k��/��5�$� ��Ijn	B#�ZjN�4��
x�Uh�D��8IGmA���X�Bef@��ɋ��]�Zz��H�'3�F�@��6��؄��f55Yv��V`L�����HӠ��\)���Oc>k*�j�ۨ��41`YB�5�N�!���xE�{[
�.9
wl�t������Yx_����v����یU�\���<5cӕ!V ���)�4��T�(=�O-�GM��pev)��>���:�	�qj�O�:�4^���r*�W�1�P�� �Xu�_�p ��Q����er!L��c�5���t��akY���T��$6r��:�\�ܜs�}�1%w�8����b]n��+��h��[�����\�8ج��T����,3�r�y-�f��M�'H���y�3G�r0��K{S�8�<�!������P4�*<h�XY!��
{�ՑW�(��(���v�Rc�Ȉ�ܮ����^���L	^0Q�G��6�K9[����*7�c�ҳ�f����:Jl���I�E��*�w[�\lD�FKLs�`�B>4P�2崙�Weu����"L�9��w�s���` ���xt�ͩ{���{
~��T��CC����i���vR�ٱ�	�,�O���1�"���9��r��S?�o����}+hAƽ����^w[tʈ�s�$β�J+�e���<����\)$X��u���D���]�{�b�\nw3�+" ��;m���=�"����3�Y�5�8���Uk���C�g��9�x�T��:�e��}�.��<�]���m�����C����j�OP��j��p���kn&��k����A,�=�r�q�6;&[�s�v�=���iY��4�w���%�et.���ے�x�״�}�b;��$z�j�^48�]ү�:}���e�Y�P��Sl|��y	�3�@�s��ǥ!H�Y�+C+�ۗ|l�ƞuN� dq��=���Zޜ��˙��|��ɠT۳��Q{n��S�l�~�g���n�pf��L����E5�\���hU�k U��x�@�s�/A�=��o��n%�^E^�Qqצ3���P�1ǯ�<�ש�{�s�}���}�|�Ӿ0�1]�7�sqZɹ�>{ɩnᬞ�<�'؇v8L��Uː?p�ZP��x��I��/'��=�(��^[���e/K��st�����V��=�e�4� ���<ٗ�.c @�厠�r劕���%����T:Fu\�2��y��G$;ΜL�vlr�;6���(�.FN�hD%�TX����f�Ck�T��7}��Q�l���|3�W�=�ip'ϊ̢��
U�����m\f�ղF�K�l�*$��MzwNm�>��G�˙+�=�lI�wO�֏{�QEY�A������Րw�N2}��]+�W~��"!�o���]��G��.�`;fp1lB�e_[�x�{<ӓ��`�p�c�[�"�K���3��ѣ���5W�u����(w{����b���[쭳�^���^��G8R1�Z�틢�4��a��z�.�,�ݚ���3+NGoN�+�Vx⌦hK���3�u���@H�LN��&\����u���[G�tg9�ށ������˚�t�q�����9��z{ʓ� �ηB�W��=�o�:T���d@��X�5�Ӯ�.�OK��;}���M���IG:d��ӗ�C�U�^˳�zjLg��^���y�;�j��]�=cn����d+����R���=N)o����(�mD����؈��=J�9�[/�E�h���閃�є�c�]K]u�V��tDjm�,0֠�lN2�eN����	C��퐤p�r���0y3n6����O��v<0>�(����Neʷ����[��Ge&pC����ݢ40��^W��B���^pm�Ttqן���5�g�W������M�z:ϖ�����;Y�_��;�ї�=.8Ǥg�Ջ����NՔ��jޯ�bV��V���Q��#g\����~��9+N��W�M�L����3� I���6@|
�Gs���ۑx7C9�r���S��
`¢�Ӵ0��3(oC�j�,/2�Ԝ�m��\��uxsB/(�8	EviUk]N�r;=|"������5zʓ��VC\�4K|���g�a~l�^f5C�"n�|�#��b��7�c!�;�o.m { f���xrkܽNhwݲ7�إ���̍���nx����Z��b�������\7A���>1�OC�;j�^�n��D��)�;]lV�����\�{b
������?/O2$�k����_+QjgO.�qݸ]���c,������շ=�o,����Kp䮝O�4sr4��e
sgu�N�J���Ŭ��:*,��a��S��f�B/��Y�o������%Ϋ��7��D����*L�]Ḑa<�
�٪��뻞��W�Gb�qW%Gw[��G���l�\�.�ŷ1��u֕�g�y���s̸͉LS�R��r�Jxn�M�T��/���إ�{Cid�$����;^�ć�C|���8-�Fgz�8�!�R9�V���� �=��qd:�i=w�{mh~�5��1�
ɷ��[_�Z'�ݷ;�栔H������n�hg�?<}^��Ȃ�5��D\�YjU�p����o�d��L���I��U��8���p虓Q�f'���<ằe'��B���g7VN�Ȑ��)?
�S����>Gl�7/|�4ʹ�6'x���<�s)6wfՏ{��Ȁ�v	��PL�t���
�G��=����5�O4j�󥸝�y+��$�]Px��N�m4�K�Cc<����N��х,0vr[B�}{�a�����2�:-� *�{�b�ɳ�Q+N���[�á�1h����u�����_�9�{���={��ۻq�V�rH���"_���[Y+�s=U �5�oPJ�q��>�8�vi�"���P ]�7R�_r��W}��G�qf=��̳2,��@8n~r��,QcwF�#J�wE�*���)��LG��V��3�Ew]tὔ�ʁ��Ǩ��ć��ԭ�G��ʄ:�TD���5cK�������7Y�C��v��vv�tz0U�T3��u(i��6�I��F݋.A�s��U��MM�`�W�2sy�E��z��Z}$m�-$���زw���3�&Z�~H5 �ۈ��ъYs?y�]}��H�L����+H�õ!N�*���;�µ�N��lc����1<��W�.=����n���Ʌ��������F�wj�x���x��뵼+tXT�T�����VT9�ڎ��Z?W���'[���t^�o�����3JR��vRS{Vd�f\��4�¢�i��n��N�s�����Bî����(ik|#j>�7k��G�T���=79�ވtiu8[ZgC�C�q�b��5��;�&`B��\#Onз��
XnÈ�zv`"�G��K�lQݽH#���iƚyl_������Z�WNA��Zھ������c�_`]��?��݃3�Իf�>*ϳ)�h���6����^7�ȴz�njR�vۢm^h�-�a�ݭzk (��lG���)!�t�8KǺ������7�5V`�oC�k)�x����)��6D�HB'b�v��퉓"ɶ�6ͣ����hI����S��v�+�[��g)���l��o���D{��>	$��yLgd4��/z�P��l���IF,��m�kwl��D9���m��9I��yLJ�R��M2t$*�I��f*iY-�T̢�E��LSTP\a�k���֤͢^2)9B���p�E�7�Q`bT��%E�j,(�ٌ�%M0�d��P8E��*V��v����'؄�lo��[�R%�4�c+��x@�ӛ��:v�}d�a�r�NRtH`�L���
�e�,�4w��Mo	:0�n���l;�9d:\��\�+������#���q�~��Q�>�.y���d��N�ќ�*����@�rkٶ��Mw�����������ծEt�Ӫm�ǨV��F�g��&�
�0�N��:gNdP1�)�7P{����5����÷ݿt�w��C�׽]�[����G<��^�gԙ�=��q����T5��,�7|���qq�닩Ky�L��4Dۧ�<���W�]y���A�W�c;��A���h�{�<TW�`߱~k*̓��v)5˘:1�lO^"O?���P�o��,8�M+-r�t�5�5R��������m��Y�����x�ˋμf?W�����ߢ�~������7鿕Q,.�Xg-HOXy�v�F�vqP9�s��Vp[ ��[.����}=&Ҭ둅�-��}��t�p�_`��:'�s�y�Wa]�pQNO�X_6M{-��1������*�Oo����ʦ��Yw��{��	���L��L���,^9�7����f��Շ�渽��=��q�#�][�=����6z+o'�}�@]$`οN&�'������A4ݕa�M�0Бv��26+0]	9��-�������Q� ��F���}UZ
-��_����10��c��v�(�����)c��y=�������G{��ec������~]��h��^��K�~�ë�\#}��X��^`�Ǽ(�yR�?b���y�9S/��Yd��=�R�J {��<����4L��]iAzϯO������A7�^��L#i<')U׼� ����so�9ے6kT��3!��w4.�k��W��g~��H|3�\A܎fAh�!�t���{H�j��m�t�"��$sU:.K��o���:b�w��W6��$�Yy�F�������=��kmƒ������{ܮ���AEf���Bͩ�3H�9�[k��0�y��`˩��9�A�"5�w�Yo�Q�6W�؀��>����꼕�|��oh�w���W�'��+Fe��\45M���B�B�]X�����`��ǯ�y�݅Oל(p���]S�CeD���h��t<���~]��R�mv��Vn�3n7�1�2r���g��kҀ9����G9���d��u�^���ƢÝW�V�k��S��-�:"he��>��:OuO�sو�w�b]ۅL)#~.&���vاAn���2�XK]�U}U_U�~\?�~?)�_�8w�l��Aa�:��_�4��a�y=s)������{ri�r޺���;o��Y�D�Oo�;UeG�A������|3a�;}<��o�>�̟���wdN\N=��\9r}hE٫��S��+Κ�ǒ�gC8�vgUz���YL״�kt��	'gv�׶��t�)s��VY��
��v8�k�s��Wҷ;-�{u7[����z%���c��o��47��#�6 �����6�]7;�J4�N3��Z8�t{���yq�-�u��*�xr�+�����+Oqo������4S��O��Er�v�Cɜ"g��}�E�sV����g7���{ƒ�~�yx:!U��/��rR�]��Qo�|�O.��CG�)v���>��t�i�&}޾�)C��d���=(.�_��B�.��>�2z�Ƕ�e��/]Y�Ii�r^Oo�9Z}g�#�Y���Ļ�ߝ��}=H�W��z?e?pE�K���9����'#n���B�{����Z��D~���=?{�:L��r�6���k����	Rt�A�G�<�.!��6"�K�D�����w]��x��U6�dI���C;����_�������y�����*�%7���{d�+Q�R��S�־�UVۛN!,�}���*����?mb���ad�zt��h��I����=<�ԇ)��Zl��}>s��r7�,�Ʈ�6�"���g6R�;˥N}4�N�X��O6������r2��pp�(����|���s�!f
�˱�~��p������@�X��W�����gu���e�jYeeM�A����Ƽ�4ltK֪4\�3("A�;m�e��>�N�4d%K�:ɉT��ޝ0&7���힖�.���}��_UO���û�l�50$�'ݳX]��{��y����U���O�p�{��yBk3�F>��/{ B�i�Of�"��繼�^��K�]:�].����`���kH�Z޾p珫�0i���Κ4�h��8!\��ܚ�؄p��@�B�����tf��>��>�r��]GY�i�"�I��k^Y兩�/��1��N�Fm���j'n�b�a}&ok��C��[�;Ϥ������R�]y�E���szE���!�5�t�ăpq�yMoᯎFo�f�p�c/[�z�UBk![�{��f�`6�ϫ꯾��R]���~�Z
�3�T�R�����}�G��n�0��S
�Ү��rl\�|�υ+f�ݾ�;[zQ�/a������+���(o�����+�\Ƕ�5�ǖ�Ǆ�9�ex�� �>�S$�^���W*��py���^��Ysu�5l<���g:[��V_u�ksyb�[&�_d��YhΈ�ܳƢ��k�5�"��K�os"!��35�$��tOJi��cF��בaͷ��Ok�wV��LD���bA�wY%#���
v�TT�?�� �fU�WunE�O�qַh
�YJ�B.0��O==��͸�b~��]�] �n��_V��4{����ܣ:�/���ǚ�^b�/y2�\���-C�ڴD/5f҂K���&�y ���"������/�����s�My��߷Xz����j,����x�{��+BlzL�]B}�����V�G3�/�m�-��g�oￚ�Z��"�}W���gw�*-��ޭ��oc���N��2녙a�(	j��ٓ0q���Q�2��1.pK����:�Y�b��B�L{2����Hi���̑LZQ8+4�EGC�2&n�s�Jwn��0U�*�rԥ��#�X^`�n��QG�Wܤt����q��RH�YR�l���̥�1�������S;VQ��#E-`�i��Ad5�r+�_Jz.qg�6Yݜ�AO��3k���ᐋ*:*�NbX��,<0<�t^^H�U���k�>q�9�Ʊ{;��̻��=�����b��M���젲��0�M�6Q٘!U�G�a����.毮�X%r)�-��/���ɟ�m;���x�O~'�D{���[o�.�^� �Z��ae��i"����(x��}5��fr����:݅�s��B�.�Z�=œ^�n-��]�����H�\&	�'C4%,>�1���]���ۑ�3�oi�¥�j�<)�E-{��@�KQj�|μ�\o2&�&Oʮ;���_!�m��K�J3�48}ϖ���-��Q����G�C��[��}Z��{'>�f� �D�Z�:��M.��S��k
��!6B��pp��/w��k�wM<��u�밶��L�nVu�r���1���lP�k�Ѥk<����h	I����S��v�R�ݹ�6y��Gkf��~w����@��^"!"$�cmN�q�&FdX(i����VL\E+��%E��'��C!Ť�TPim�	í%���1�ȹh�KIX.��I�n!D���@ݱTU�Ub�"T�iW�q���
�ki�L�Wj�Ed�l�-�U�R�����
Ш�,R"��x����*r���C �%<!L���*��kj�+��6:l�u\�ܸ��:WÝ�ſ���ʬ�w�϶N����B�m+������R��>d���W��V�{+_�I��ü�K����MG��}�B��j���¨����z|��&�n�K3�.X-���zχ��'w��]��3x�\���m���������e<���e>vlK9�#*�+�3�`#e�+��݃�c$1J���H�_c�A�m%S�/ )[(�;~���Vݲ��2��^����|%ea���;��7c�L�З:�z�:OBY�u&����3�R��K�zWPx;(��j<`���W���| +���bd7Ӵ�i�a�6,Iu�{���3+q�;���VO�����sĕE1�.%[3Ά�*��`�fߥ?ʜ����S]�9�rң���E8L�.�7ٮ�Z������W9��Ź)4RxV��c�6��鶽C�w�f�6h�k���3�m�Y}���xk�C2x�@u��QGo֦��8���=�9�{�cEJ��7��~f���t��J(������>Ӣi��( �3'$$��3
�,Cd�&������ w!f�7W�sW7r��?�U}_W� ����R�W�6S{_�^#���!�&˦�������x&��!O1^k�^���	諝*ixs�P�:��,gff��\���au����}Ԁg�}�^��]��T�g�_eU��i^uĪqF�7w�0��e	���nR^�=W]#�G��w��"�<��ƯXꌍ��n%{���2�{���7��ޙ<�sT힇}ǟ��.����Q����k굍CFs�&ǋV���. ^#
Z}M��*X8� �����q=}���ګ��SI��r�l���O���W�UEMfr�[1���Cɞ�η��X��69�=��p{����Ƈ��MԾ�8�v�)��;+��nОA+����;NE�>Y���RDX���q�C���t�՚V6����FX��+5p!��"U��y�w���TܗՃZ�Y3��e��">�r	3�k�J��o?T�u�Hmt�B¹�]�ȓ�yy�3ͦM�b��=�k�q�f"�l��vo-++SBYx+J�8�cF�˵l[2܍�)N0���U��D�𦭣C_ř����tx���rI�y��Gƿht��n&s�nr�����G��ᡯ,���X���Y������oau�<�x��2���p��Xn닸5.Ԯ�5�[�y}�}q7�ql&��fa����uߌ��y�*	��yDXԀ�7�/u_��g���mz��u� \�v+�=�y�۫Ar�J�OY2φ�L!�6�ˁ�ܥ�܎c��Hm�Mt�5���j@����I�9˅{��-����%Pu'���W?;)K��V�'�j,i�_%��n��nR�m�6Pa�;�yA[��W9����Svyq؂ܶ�V����1s��W��S	��:=y�ݽ��
��u�+��g�c���9�1�Wa���܋v��8��{*(��tK[6�����&�G�k)��V��$&z��퇝GQ}�N��ϻ��f�sxz��	SK��j�?��<}��g���3�"a��[���&�wl�8��0׮��������s���=�O�u���Zyz$;��O�o���p'A��v����Y�,ߞ�**�b-y8�58󻚟hd�v)H�f�E�ڻAWV�+`�:������+��r���TK�OZs��n�}����b}_J��mM��N�(�+a#�/Y��z���xj�B��������=���lU���ꋔr���!�|�*�l7�3Κv=~S�O���1^�㞭��׏��r���{�l�9���t|i}�I�"��}*�8���L���[�m��Ì*#ՠt;�����_���c!H\*X^���T͞���B���U%~hﰲ+7|��P�yLn��e���\�v!˝W�뚫�g�D����pP��6 �����V�vE����G�S\N���O�}�}TI�_��Y^n���T��̿��c���_k� �H�ړ+��[�h�s#��7I�]�����.�[�����O�ng�������Q�����q?��S�<����R���T'��(��Gf�p=�|<��*?��W�6oA���ť���E����/��nI�ϟ.=�=�&��hE�=w��\Ni��E��jV��Z1p�{��2�^�{޺�/�����*�qkk,Ω<Tš�cs��I+�r��c�
h�f�[�jP#�|D+���u*[��W�*�Gٹ]��-1��UUW��I��~;��f��+<חoc�$Z��(T�n�\Sjq���Ȯ�F�^��64m+C=5l�⧞&_r
��[��L�^x�&@��L�$�c����R��D���Fttn�ڋn&q__C�x��F5<q��-\�E��[�-*=�qj�8(v���_bS�.�0��v�Tk�A��#���jrR���y���Țp�Vx� ���z<�����h��;��C�W*�3��n���
��rψ�=<��n��C9Z�#@�]�	��2k��\ϥ�q用��u������������Դ{=�2&�w���+�r�?�"�o(��4�8�\�z�Y��}{�1餏/��W\b�;gb*��ꭼv�e�
}eu����Jp�47�{�Ӹ}�W��{]��}��/�ϟz�89��5t#Q]�ݹg��t�p�����G`URc�S��古���7Ƕm`�pv�tx�o�����׶��AG�Kz,b�5�y?'��{b;Y�7�נt���|5t�[���/�%T�a��4#8�^�7Q�VmЉ�㲋��E�h�n����	�G̾5�g;�9J�&��c\�.�
ϋC�M�����狵��@m)�������m�ؗ!]Le�=��)ж��|��g0�0�ʍjo;�Uě��Q\�i��Wy��v�F^�>�Yڜd�G+�µ��fR1�b�u&6P��y��5�����hj�C��AXT��ea�#9�Ƒ
X}c��M���Rj����,1
����{R`\'0v�ޠ��J�|��)b�mv�ݫs��@�7Y��k}��:N�n���/��\-���kHb��V!]���k��Յ��ի��x@-�͵\�z�f�֫�9���H��{t4����ќi���ɖ��<BDe*):�f�]�
\� %���y)�ι�˕|e��ʆ[����!F�riޭ�ݵ���w�0v��p�������C;+����V�0��᯸��X�}�N�+�&+���QIi���7��5
��|�hҮx�m��~�2�RRvJ�*�������S��f��o��ܛ�ҋf��uPjN��n[oPy�7�ޚ�׶� R�3��H�#VWH�Ag"���79�����O}�.���vT�Z�,`�{v��N����he�yt���wwwiE7�ف����݊.y��v�}� (?�$�I��'�J��*�LNR��G�Q���*"���fXT���G�^���Wt��j°�Q�Eݫ8�r�(�Q�DDQb+P�v،�8�P�j6��7kmdv�*�"/�o�LE��TUDX�	F#Z+�*���*ESY5�9��X���<���QQ�ETt�H�1���!Q���A����C��]�a�q�s�����v3Mহ^�[�a��Eٷ��?���ѥ��q���qk��w{����i��+��{;���(������h�X3zwD����uHҋ|-�oN�P|�<J|��ugTK\�5W�3w��3:ش�z����&Q����{�"�W�*uX}�����BH�V��z=�4���>�ڵ�}����s&����ڸ�U����s���q\����z�*�ޮ=����n�׮�{����F��x��iF���:��I��m�
�iv�]ۻ�"��|0�'r�lu�n�n��ٛ����XwK�ݝ7rsE?�}�� ��_����.��O>�-�Y�������Li+�j6��()��^�25Ѩ$�-�x�z�w��Q;�����O�O��}�Pk,R��0�v��^�{����F>u�+f��۾�X��؋s Xu�z.����7vөg�>vHLo��M��]e$�y!�t�+s��ị��W=G%1�Ǔ����C�E.]����x麨|�|�I����*xzn��ݔ�~[��2�P�� �N{E��Eܽ1r�BRuzЯ[�5��P�s����6�խ� ��?l�k3r�H9�v�q��Y;����P	6����R���1ɔ�ﭜ��h�ݓ]w]�z�M9�s�אh�Ѹ|_�j�S�[Bpg=���c��'6�<.���b�5Ro��y�9��Cb8��+��)�����ኗ��^���y.�5q���s�TW\v��ν�s���RC��+�a݄�(����/9��1M3[}}�^	���!�;.��u��b��K�����+}��k�OOUu��MyOq4J!m��d��.na'�R҈腹7�(oX�,N���u�*~�������Q��>�{��:^W��#�6���,�j����>Bv�yv�.(���d�)���J�O<˺+`~�^]X���2:�9?	��C3}��穉�.X\�x[�Sm��wW�u�M���E�r0u�Ҳ#�'Fe[�^`�}����Nfc4�L	�R��g�D��ջ�k��ty����ٍ��{iV#�bq�Ҝ��wǺ��׻�����HKݧ�bl�%粖��*�G7����Q�2���(,J�
Wt�\9w���`�G�)��A�sv��ۙA5/���[}�� �l��S��}��ڲC��.>��E%�u�i�[>^�c�`�.ɬ�uQ�7#2
��q�Wޘ���=c� ����jѕ�>�{3ܵK�L~I�OM��N�鮭Ӛ0<�ܽW��Kwԫ,�j٣�K)�}��x��Տ��\�ܝ���mOg���G���#~�qzWw���	yP�r����n%z{��K��9�01�Sۭh��,>����4'FD�� �J���{wh�ص�FR:J��-�f�B�����y���J�=m�̠����}޻	֭�x��W�V�K}�󟶦��'"����Ѻ���N�&��i}Ѳ�M��XE����t���q�<F�Ʋn�CT��3]ԭoG_[�[.��U��O1����zH�6�_�}!\t�f���=}�R�K\g��c��bh���T�ǽX+ �fu���;VZUe2�l����K����hݟ���a��.�S�����в��&Wtj�z�>�-J�RՎa����å�5�J,1�l=�`&f�}DZ�=٫���WLL��Jq��A���jթR]Z��l���n�4�6�Ne���(�2W�〺�U��~���8��s\�z�/y�/0��=�*HWj5�|��d���$��U#�I1Rf�џ2Xrwj�o�(��ʭ%3n�t��Ǥj�X�,��=7����3�����g��Ӑ.��������h��g;<#��`��9Fm>yW���!��7{3l���Wz]:{�A���1��-s���{O7��M�l�="��'��ٓ;T���;t�m��]��я"5%�0���@����w¥Sq{���cTm�������~�8b���̹KiXw�ˀ�@����F�����ͧc��n��}3rF;٪���裡��i�;!H�]
�jY}�#�����"w������ٔ]p�.2<Ф�:��68�L��a�G������y0�,�y����ѫ'b��5������W�Гy�cNc��(�r}֞V�h�Ѫ��Nk���ܙ��<2V�Wx�ϕi[����&Ԕ9E�yUԾ[{�G��*���
){<w����\��듹f����X��o*�Vv}5`����3���Ύ��m���Q��O�<���ϑ���|�/�ud��	��䊷ɦy���o��$��n'�V2�9�ଊ��h���$�^*)�EB�D��\�0n��9��A��1cT=��7�W:{!��+|�n���hȦО�_P���|�\o&P;4zu5��d�
���TN���Hߕe�ٺ워�H�
�8�t3R�|is޺=��*�i]$����G�^ll���|�j��1��-��sasNeۆ��;��4s��C6g;#X+�Z�-����2�͟���V�g|����Z�&�}W���!�>n٣�b�{�.3��v+��P�zvI�銞�ho�5�ڼ�'<F������1̦�Y̫^M��>$�qE���L9��Ƃ�%��9�`�eZ{A�^��s�e��FөO��q�0վ�!�	�oY����6����W����b����q[��y�(*�E��#�� Q��pN�l�Zyغc�֎Q���N�)\�Yzz��5���ܦP��sb� �mz�Ժ�YX�s�����B�f�(�\�^vڇm��r��s��<�}ʥ�0A�XUJ,�[��_[7f2>ccB��[������l̫���>g3H4#Ỷ�!y݇U�b,$��>�:�-w\5hk��2���u����ي����*�=��<ݓ���C�},+�7�i:��<:�{�k�o`�N�Yq^�9��:޻�hm�x%�GN�+@�X�' ��f�&]��+X�fЧP�t���#���CE�Y`�)���{jR[uf+��r���l��Ι%_>�qp7���$N2=r��L���#HA]�kj@a|9Sӻ�`R5���?��� ak�s{�%�٫����H6�$�|OOE�F���N���:�fX���Z/J�|����Ps�;%����jq���	�[�ά�O72�p^Y��|�9v�9�bdof�)�[hSyI�8b.�e�*��o��[���b�PDR����^<�{\8	�B�5yc5H�Gy%i�ܹ�эջ�{��V1bI�>�{�m ��O^3��a���b�x�麹Ul�]z���Fˠ�\�s�p��m�ٗ��ok�=�]�bj�)�Wd�x�X�.�78��^6������Ք���*.�;;�6�ث&�%�h���n
�������c��v�#ԖF E���6�ss���M��6Ҝ��˶�D\������ �DN��zP�g[�QdUQ��ETQ�*ܸ*(�2�M�8�LjKB�R�KŘ̌lq.�W��h�U��,DH������������(�i.%Tv�(1G�Nm�Pb�����.C-N)*"��h(�7v��AiPAQE��1c���*�"�U��ST���`�Fv�Uc#��z�����^����)TQ��Md|%��mhM(,UY٫�uH�1H�ۻw`�J�%C�t���X-���o}�u̩.:�f�A��YZ���6��/=5�ɯ��
1�}�O4*�n��Y6���37s�^6��]4*�c{#��n����ż�"jk�~�p*{������ާ���R����v�^�$��9�k����v��ɗ���o���qZ�W@�~��;Y�BH]��9�L���QQ-�SH..��yj�����^���
v���J�K���_��si���^�{t�*�&�x{�hn�vC����>c�v�p���ܴ�U�|56S_�@����J+���������L��,��$�������ʝ����Gt���蠧o���\�ڗ�Տm�S��'�ڳw[���=ة�wg��p��a�w6��G;�nq%F��}h�X#�6�/���vf�{��7��^��*m����$4�I����H�\�����-9ڌE�o=�i�ѿ|l�cau�c{������=�Z~[M�^��-�v��7����n���l���r�nv؈�g{\8)�u�^���	R��wX��.����g�ʬ()߾kKO�/�E`�N�~͝��Qk�����C�S#��1���]yХ����M��z����/`�-��Rڛh�����|�����4�CϞ���>���e�"���|� zbꍉ�J=���rO+�^�ʆ(8�r�G5ž� �-7}	��#M���W1���h�/�w�k]���'�u)%i��\�7&q��s���Z�dvAJ?Z���1u��I�o�Հ��}�6����[��eV�뫃����{�N7�����������ow����� �o��<���'�ߩb�(�x��D�^��|��6�\��;�އ���Aɧv��͊�U#�+������6�f��/>+
��ة���
�-�OT<(?���yi?d[�X3v����6}���'w4�z���T�;�+�Hf��U��kB��59}��=�Fp���5<|�z]�Ν������ms�#������z#��� �㚟8ӣ*)�j��
��w_=y�� N�1��w��o+<��C�z���h��'a����W[սX#��%��P�WaN�x><��}_j#���������GG�Z۵�����Ģ<=�;o��}���߶�>!����#��_&}I����>�4��i�k��ɅE^�:��Dc[� 5�N�]�������M�0�>�=��:..��\է7nTA���2�:j�R��6�6��ۺڸ�+2n�]=��{�8o�ʣ�zy����^��B�J����W23�P�1��ze@�MJ闵���f-��t4J
�bGt�v�e����b���{�������@m^Y\�svóݥ�O�;,�F���v�`��T���Ͼ�ߏA��z�W��k�f�m��xy��"{~�Ȼ~V���u=�43Ճݡ��QY� � _m�W�$c���ȵ8t�q[<.g:�;m���F��0�����`�Ws�R��#�7]B�\�Ft�}'���jy�E΍=���V݄k�,��f�M7�g�ɒ.�e�:�LWG�Sh�Ω��������Y=Rj�P������i{�����q�̄��ȘA��X��?k��s-�Pr�i.��M�'�jӰ�+Ym������y�L�
��]��k!�O��^慄~��P�{u��kI��u֎�b�_f-�dm���{b���u��.�<5�����?9��.��	�.������f��Y=��Q��[�pw�����m����$53/���7���X�c�ɘ�!q@�_#)?c������7�U=q�/;�y�y�0��Ў�P9h o�wZ���y���9^�ιq5��tm��ׇ�ksD�P��OW*E�W���cȼ (���S�WL*ʝXdۉ)E���\��uu�vV}�%� ;�V�Z�F�瘳9K��﫷!�(�絛�i��ei�����5���,~���	��:�B��LWC��c���_\w�Qۄ�����^T}�uІ�)+���jI��-���x1y�zO7�\��ō�8|��X�u�ϯq�z�q�K�9tI�r���܃�	a��m:�A�<y��W�:�z:֍�[vc����;�6��iy�;���mlކX���~Am���tma8k����y̍��D~����4,|���֦��F���؆bf1G�%�vڤp ��4���K�fޮ ���e��S���n���7����iI��ޞ\�W����S����0ً�V�eЕҞ����V]Ys��P��x���������b��_k��-�1�����z"n�<_�q�h~�)9��6*޵Ig�����]��§K�]J�I�u���F���^p����t�I�E:�uG҇�sɬ~�5+�n6#�Ѐ�BMJ�Qś�GtOn�S�ڇM��u^!u��AY<e�Vg;�P��������ʖY@��E�D�󶉇�$r��g��^�C�t'h]_%�l�O����]|V3eG�ƺn�z��#������韛-����k�sy�_���>��+p���w3��R��9��ᠪ8ӡ��B��{�v�4L�^BW"	]Hx)��������eMGq�i�u
�zܨ�K9}�w�:gv�"�{3�a=�Շ&׈�����Ľu����Ut��+5@��O<W�&���K��]�@�{�����ۓ����4�������w�z�s�V�x����z����Y�P�u��E�L+m�V�i``��c���/�0��!��EL�0r��X��02]��j1S��]��
��`s�cM-W�b�v)���͠JPq�`�V_�I$n�ݍ�Ż:��7Q*�6�;���U�#J^C�b��
��%i���n���hn�&���nQ���t���Ã���'\ �7�'�W����%�p,�*wݬ���k*%��m�����elP��l3o��ك�КW��M�����gFo'�K&��W^C,j�jh#���6���0nٴ�%J-��]>f�	#(ޫ�x�[\��nvJ�EJ�z�?z��5S�`�<Ws���(��,e�DR[ke�mQ��p�tI�nf����l�-e�=vnAK�'r���'_�%]� �׀�;Xa��Np���wP��ӥG32��Fj�K7[H�{vI��h���X�P�1L��8�5d1&ᯝ�ލ���.g��j���?��R�F�3(SF�4�H�M�M�Mt0���ΦR�otj��p�N7wmT�U��#/6Ki�:$�pX��is�uvF�8���ѝ�d݈��2Ue��t�9.�n�G/u\��7]�+�r4rC�X�k�P.l�y1��	��������߸�\xv�^��u�-0O:A�m!�����[=YA��"���;��	Nr}�'�����Ҋo��8�˦�E��̶��,�h�0����mQQb��E�+�U���U�����"(���F(�)]�A�(�{%U�J��j�Nm�QY壺���#�i�UX�e��TB��Rժ�X�1MТ���o*�͢�,TAUX�
�m�*+�((s��X����yl^iUb�Gv��EPx�����Z�"	�RT�2�DQ�VcS�)��Rm��QTd�-+Yi"Ј ��/�|���Nl��{�څ3�ݛ���a��Wלz�㻣5?����RM�}?��?S��[^�t�k�k��[�6ۋ�{����{�:౅�ٛ�#~���ǣ+��Y�B۳ܵ�*��Z���հia�����9���2wϞ�<��+����6��`�(�iI�J��|��<r�g�ŵ�����֭Gϯ�Y�^W���Z=|z�8M�J<>+p�D)7�3�s���{;����'9��)3��|��,N��O��ɯ���^!Mm��~�q�h*�:�S.��	�Q���}�5<:�Y�]�q��e�E!7��K2��}���2B����Gk{�U������nݷ�!���/����"���@��Y������)�6�缙�����&9�|��?Pz��2-����ǘs���K�Ӊ��q���va��E��^3�n�z�23�݃#I3]W�R�6YfGf�#YB��{=篯���&Q�9��y���ר���(Y�ʥ xl��K!J�iocNS��7����������Q�^���=o�S��P������ii�J�v%源;C}��[�3����ܙ���;��Ct�8���4�����h��C��3㮷�:�?���8��x�tyZ�*9V���ܽ[�w՘���P;\.�rT��q>��v���WB<]h#����q,7˓�q�Gӊ�L�^�5;����`�O=rU�x��iS�"�9~�c�R�;���{_�^�6+z������r��t��:t�9���5�پ����?���WŮ���9�n���ѥ��3uܰ��.���չ?7��ںlE�d1w-�����0���Ts/�g����I��N�vɵJZ���1�:��7q�cy���̼���1T=`�.�.��`�k�K�'*;{��.��:Z��x1��X����T�u�+�ͣ��)N�ʖ(���N����ĻpN�2��X��^R/xR��ƪ�vlr��]�|7���vZ|}͵.�6*-��ĺW�Q����e��FG|��:�������^��e��=���x�Qs^�%/�ׂ3ݰ��X���͚�hS9C����Xǯ+���L��k��2�m�0��Y�]p�#�F�Ri9�4��V��,�����KNoR�ʇ;'VX�զ��똶�i'�� ��sq�� ��3�L~9�|���f�sU�c���@�k�&k�S�,�Ӈ�햇�2��%��r��7g�CX���c�y��z�.�Lc]'�-�{�h�h��T�HS����M�yJ�Z�ٮ��s�
�ns�h4���0H���궸S�ދ�<�J��h��[S��z�_u�_U���Taz�;�z)��]N��!C2x�ʶ�c���f�
��*��{Ձ�}�'Y��[�)v��Iq/?
�La�ڰMY�b߈3O�%r���fT�u���쳄�߫����?7?�k���mm�o�U�O$� ïn�E�=�I��U�h���p\�gl��fW�8�q{j�XKDWڣ/kN�X��O7rh�I>M�:>:�G�����~C����r�	�|w�
 +�ѩ՞�$'8ꋀ�?h��H���-�=�!y�#��Y��njq��:~���Y�u8}aS���.�U���V����Ϣ�*��gj�u�>z+b�=�;6��QwY|�3A(�X��L3��b nڶΖ��ѽ�C '����wGbҖDc��(A5��b��Ȗ�3����?X�.e{6�A����q�s��`u�����!����ղ��׾������j
{���Y�ը�w���Y3��9��w{|BlSXڝ��?eu���R�s�ֲ�62����쎆�v$gu��c \��s�()5�+n*Ԕ����`�!��N�s���퉋���;�ل̾}�?qz��H[7��{Ґ��N7�t�I��^""(t�����z��:ҵ%���Α6�}��`��yw���w�Wz�J���]��f!��EYe��u+��znC)�+�[������a\�}VJ��W�MP��R���}����r.~��h����6�k����S]2�5evG�����w��L,����-b���W��S�g�C��hڱ��T`�P���{6��7��:r�A=�m�5%t)ڕߛ���2�5����Go�"��Wv�*�u��.tj�;o�C���w<BV�)WdؑЦ��\���oV��"��(�O}�Ӝn���값����q`�1���_���'�e�T��j��M3�����]�3m�g���Q�-?k��o�����p�1�[��skދ���)��8�\�SuX���zOm����hs5��ק{%u����=�Np��qծ;F���|��{}	ث���!Y��V�u���WO ��윻��yhOm�L��N�{'J-�>kw��P�.���,Ҳ��0<~`�Vo����S�^�8�%H8�� s��Y~^��Š���`�a�B���&e!r.��06���r)(���rR���M\څ���F�ڱ��=o���(M��v�J�H��x&�v�nALͫ@�:�.��LTջJ*|\P�8�E�SF��A9���{YZ���8�zǝ.W��L��|�S���&�[��S�e�Wo�>)��^�y�@�����{�t?v=;��D��X��ڎιP�:�,�݂��e,:(��Ls~�m{��}�Z�=�=��S9�g������Ӻ}gƼ="����	�K����R#~7���=n����󩬨����ma9t?�0=o���AjN���N���̜2�l0d�e�ڕeաr��!�u�eػ�|����7��n)KF�t��l ��ι�1|����� ͬ��48kS;1T�,
R��k���wB�ɡ���"��Xc�헩��t�r��B�YH�"��+��1��s��ٓD��6�[�q9u$y�Xκl��=��K��y�)���+��ې`�	�y}�L�i�|x�]u��s+/�ծ�� ����P�#2��ų�ӤW�̵�*Ga����{e���I����:�E7rig;i��^*"g�C:%�e�����gQ��M�������V�z@������hd���>LҪt����'{5��k_;��%���λ^������q�+o�u*�C�m�b�恫5n���ys�9��дg>���6e��a���?;�E���M�+.e�-.�&,]��pta�����������S�H����	+��@dj�G�:ɗ��l2�-��p>n�$@��B�Ԩ1i��Z�v��K�W��+\�B���sw*tS��v�"��4�.�*�4���f�u'
����l7���D�3~�DԮ���yN�QQT�r��	xqրx�ӗjH��\3�����e^H"{�cNu���������7����+ۈ�
v;a�2B�;�$1;@�J)wfA��R&�%@��R��BD�%·%�-�8ۦ휇��8 �rs�O�>�I���m�+#f��y3o2�nt��E|H �ҬF-�Z�m��8�M4��o\�9T�U�啙[U*���((��(�!m
ƔPmR�7e^�
3��uN`���0�Aq*��NR�@Y4�D�Sl
"Ŏ�b���`"9J�,���1W�D��aQE��U5KxͰ�F(*�b��c�i�[�%�� �E6���:��Ea����+1�!�5�"`���Bq��tި��Q6���2j�<��a�9����ŵh�`���@�������Jn ��]ln�Ӽ��{~��Q���*�s�*sӭj���y(Y4%uܨ�OASy��M
��C=���B��o�^���OƘJ�]Ύ���ˎk��]א˾�l��X2EZ�\4N�[�}�v-�����8�j����ҙ ����a�S��Y���ׁ�C�̆��[Y[<�wʃ��\7��%=tc��ɤ�*;�Wvb�����4,��u:�A�N�ݹ+ܬ�p���h�9�G)�pv�efK�[T'��p��N�Ś�y��1O~[�q��|��ɡ����3{��I�ԝ�Z���{�l�����Ūs�ST.�z*��y������fa�\�.���^�NCاU=��)CI#x��q�R�S�y�p�9~�4{
ӻ��v�	���2�� ����:\�8�w���o�ob#������L�_�H�-�t}�6<knf�&��Q�(�h�8b�C�@=�n/C�W�w9��-��X!�ܞ��&o�b�+�������b$Q�}7��J1��vjL����������/��x��ǺT��xV�̬.r����i��&'�[Ǒ,m,�4�R�����`�7ٛm�7)��F���}��@�Ѡ΂T4�yS�<�懕��]w�6�ِ�y �g�>]6�~sKm�<s��=�=�7,{��� �?p9Z5Wqү�y�����Ny77�F�ʊ���G�Ы����O�kL��\�̼^��=D����F�xmǒ
ˏ�ٖ݉0�A�UH0��n:�W!;�<4_b��S�2������Qwu[N�T�Wհ���Qo��~s5=��9�8Һ�s>���n)�]���Vv����/���t�����M�!Ӆſy�MT�޹�AOPJ{�(�<�!���҂(o}��OY+o���چS<�q�cuݩ�[�V���B-�xܕ��7�����牽+ڮ�v���g)��n	YJ�;�53�\_�����Fdݼ2�W���ioǤ�h��y�)�W�{'�^�m&g3��LӔ��f����֪���÷s�n��t�fu��.tF�Qj�B�ZŖ�˥y�y甆�3�o�b
���]�ziî��<�=��C��LR�]#�:�j��ʮ�fz��F� �Ƶ����R^~/����,n��2G�6��>s�8]���q}�T�C6���:m�2fU�8m��5���std��j8����D�Ǯ�(Sx��p���	�֓k�E�z�V"=�ۙуF�n��9�Wu?z��Έ#5qy�w8dr���発1�h��
��gw��K��d�3/�*ߕ��]tr�t�0��е8��$�\0�Lv�0�N(�x\
�U��ѐ����]�XXR~�c���l����^zb�L�`�f	�8�h�/	��Rw?��������r	��کp�]^��T�͊{(g�l�Z�Q�_W������Zu��c�fu�3^��+�8L�.KݮA;�s}���w�o�e��Jq �LX�G��m�\=��1�X�f����������zz�*{LĦP�����h/KO)�;�CՇ�V�k���Y���~���hf�'�q��Ez�F=P�b��T{���૬BM�'��225�0��K'#b_���<��c�d��;������E����Б��b���vk��_�у���}��/;鬎2�:>�����>i�F�S�op��{�]c�:id�Y�|;{"�W �.�]�w8~�c�D��{�{3ĩ�'�y�Z�k�q	�d��l�9�̅S�l_>ȼ����y�V�����5�h�n�V��Ϟr�����6�D擰�4�|�A��7���`~sR��y�ѾDx;�N�#Gkvn��������ׄ�Vg%+e�l�VТ>i߹�H����L�����[�hj�s��=	~���x��9?���V���
M~v�oi��ӧ��r��9���~�P�ԛ����'+ʳ��ބ�S�d�ԧ��J��pz�xWy�=�{�(_ _�x��\��4oX�ys��U�U�	�Ӑ���x.K�y��)^�%u������ڷݰ�&�{r_�]��33��S�?e-"O	��\�Ζy�Ǣjk����r���P�b�Nܓ�0KeC��ws8���i�������6Xv^���ूE蠬��z�kf.��R�U�Jx�v�GK������%���ѓ������E��O��<Y�m3Ey��V�}����6]���GI5�ꁨy�FsŪuʢ.��<6���u����r�?@�<po@P�~����Ǵl+�h�ZE	�{�!5��Nt���vO@��t�J�=7����&"��* �y���麭�r_!�B��5p:l���A�c�����[��6+����<t���HN,(T�>�:e*�ˮ�wʈ�����&d���,7���e"|��*|��\µ��`�w"�ѽB�=�5���-�˯F���"M�#N������G���in&�!��¦t���xн?�����*E���u�M�g_T���S�1c%�\U�E��wen5s���� �)�>�Ywy��A�����?u���z0�J�	X}�dr�	۳��羃t��<G�������|`�p������{�4��3��>�8�:�,Ը�"[�s�W�v40��H�nIG�b$Q�lыC��B��Z���'=Ȕ��;.���&`d@���6p�����]�m0[TjU 7f����fo:D�G�^v����7�g��G}�i���,�)7��4t�\EB�x�����u��^�@%�jԠ�?��?j&r���aO��f�g�?E<E�p� ��,�!p�+���5�g_	>&_�@�g�7�%�f�p�ۨU}��Qu3?~P��A��ќɐ�����2��sͰ������re8��YL��-��W�<*�7O�]�½�m���)\�T#w�(��V�ů^��r떗��h�jQ��l��՗0�/��l���+����t��rQ�,n1�����謬���j��ɣ�i��╽r�kM�k9ΦAh� U���&oWi�a��9��ԇMD���1Q����Jw����Z{�&<ط����+�ǝX��0[�wfa��}�w6MMLb�m���B#Rb*ȧ�DD=�I�O���d��i��}����;Ѵ�FJ�oТ2��GPs(�e\�V7UA����J���Kb��S�ǣ��'��ى:��f��|�Io�ө��Z��p�4���;��u�w��^�)9Y�$���e�J�4Aye�7X�E�qؑ2H�0���I�arT��ְ�'�}��j�8�^�z&&p)�.��d��Mۻ�. h�K�.�N�*����`��Ӕ����j`�(L
�j%��7����t��VI��V�U��N���(t��,t����-�z�%�f�u�8����y( 7V`��*Y���{���v`�ҕ�wu�pkh���p��vV�"��5Z�pȐW�L�j�f��t���D|�\�a�I���y�v�ƫ B����e��i�++C�b n|(���1�=�S�v��n� [�nrI�'����JM�v`Ű�zsӡ�ju��ws�{0�!�+dN��;J�z�C�16�V�I�QE��,�I�1�(E֬SkY�bb�FTR,* �m��-"�&ڪ�`���� �Fi�$Y"��*ɴ%E�F""sh,i
�*"�Z�T��0(Ȫ,�E��n���TS��j[Cy�"�V�ʆ5R�6���W-���%aE�%e��0̬�aRJ��0U 5A��U�@}b��܆���i���>L��p��n�+��%t��;Z�������dǃ��~ŞXE���0�cv�KBN3X��\�l��mabS<f���G5�[^"oz���^�͋����,�$�Y&\bV�C"3� N���7�VwG��j�V�#�s�x������o-O��+tX��%a�>C^��VP#|����)n/^q����U�\0�!��#��C�})�H�FR�*wք{�>ʫǘ���K|��]-4dFls��	����{/P���	�[�J����"4!���ǵXH/8$�ߦ[>յݘ���)
�6(�T`R��}|P�.1Y;�,3�7Z0J��Yj��RDr���~L���7y�7n5�)ڣ��#4̸s�:т��R�IL#�Ҹ�Gju�[]���!�J��ge���{��o�_}
:���A�P��ADę���/~���O�S�N����i�KkH�0��#�jo�����t��r&�jփ0=� =��2d����??�����_C6D�zFb�ȝ[�����-uo�H��P�P<`LC,�����"�q��O ����>��	^"L�%z,�6k���c��ˊ]��9�ݞ�Q��t�E�?UX���	���<z���V<�c���Zf�8j�>�BO�"�g�v��I���;�7���B�Q上��t!�F�6�%�]g]b�-/6t�-0��zDyQgK7+N��l��9�]x�P��{������Ӛ���roh=�Vv��C�\���3�`s���� ��vZUfe�b=�Q�˻��C���a��Z���i����6�B����e �W�;1�d�)���B�/�<j�B|��hG�׻��\�������2�>��#ǌ�<V�+�/���6��rK�8��d٨C�9����9���7����@fӉ#-8���z��F-�.��Dz�.�Ơ������s">���9�9�e�8D8����z��γ��L}�=G��T��!X������.���E����j%D��OJ儗����Y��Ng�r>퀻b��B�!�Xe+<FJDp��(���f�����=L���_6~s6�3b�{�U�4��������7����C)P� �jwg$���Է�Z�C��_iQ32����& �aX�a�\���)Z���rr�:��ii�~�3��i��,��O�5c���n������C=�"�0hjg���d!����x&Mx,%��Ĭ7.��"GoH���3ݯ�o�E|~�H�.!��p=(m��-G4!w�w��_wk�&�#=9?G�	Y�X}�����s����H��=!�D�J8��.Gݽ������{3��j������'�
kI"�!f�ͿO��GԹ�6�ǂ
�s�p�${`�dY��tz^{=�hz�(�������8��;{
�{�m�g����ފ0%Q�4C�L�o��Z�W�|�af�u0Eh�Ȉ��
��{��k�fΔ�IL���ףf�V1�A�+z���P���sK��r��KOqo��:~��8���s�ڻ*�HY�R|Y�ZLmO�ޖ9(�_��싔 �����DAx��;ډ�z��aY�����e�,<`�\Fk�������so\��㷖�Zi!p.�8�4�h�$a��F�&ׯ�w�R.j4�sU��+�3>W�ig%hJ�p�Bp�t"H�|���fR�#�:C(ל_(p)t�Ͻ�]��QI�@�VI�/8{�#s�1w�����vx4&�ds��U�\A��8��T�g����W�p����S�#��7����f��z4��>/�rr�����!�@��@��8d�Iih�<�ms:���Bb�����ty��f�{ ͸�=o�/���dt�ب��q��Z��f��su�nZv\+��U��c�_�"�n��3�֙�O�W��i%��pM��	�波�)뾶(���pL#��d��m�G�j$z����Ϻ/�t���k�4D�@�\Q�*0)a~__)�\Gb�MC�ɷ�_�q�4v��z$��"�����3ݓ�x8�h��Dy��Ȓ��[����9�������a�
:MLj%y�#��ʸT_��)v8ڵ|/=��^�/3jux�{�x���Mz�fb���Ժ�<�Gm
������,ί>�]��Q��z}���C�@�b8���H�ּDz����4y�����T��DY1�$ٯDy=wqM��g��U!�WCpM���: ?fF4�����!�ۦ���ݢ�^�;շē��g9RAu�ؙ�s&�8f�����";s�ܿ8z�>��ia��c���	���~�{4��]D�<�(���V��!'ܰ�B�b�'�!�暯W�Rǭqt��e ���ǈ�L��ֆh�F��;�o��H���ܼp����1ޡ&�:Y��k�Kɻ~�<h�:И���Ix����!j���{&��[w�|=���$��U�!E@�dq�DP�#L��yz��|=�JOj�^��G�q�ǡ���`u�V/M��s���G��G�	���pH�0� ���0ӗ�=N�\�ھh��|Y��fQ�4�b��!�N����NNnm��P �/�0Z�$��ZD��8>���;����.�N��NH���fAgv�,���C���xU���<z��8%ݼrk=�'pt%�ܡ|����L/9�݉�U��y����������~�ԤR��"A���\}��wd�:���{Q�x�{��s�/Q=(M�4��7ڻ�ϯ�:ORoP��#' �4��f#�b��ϧݗ��l�Hd�a���<Ej�?8�O��;�=�לϪ U����:t�f��$��e]ej]�������ܬR_���I�3�F����\#ݭ�"	,�.�'�f�@W�=�!#���{���ZIvb	:C�ゐ�2j8�R�M��8��~;5��{`A��쏗儚9+����|{s6�6;Ha\̍<C���_:R��Bˁ�}���VmH����6��q��Yڙx:��:����G!���͝	{}����0��1��>}�ɑ�h���Ͼ�DM�r�3�5�/����52O�B�-&�,��k�q�uU��4�R�BmI��B|��$�j$Qvo�j�yr9a��;HsCai�B����F}��,�Cq���3;=�Q�$�w���DG��H?Dj�
��:H�u����؂���l�u!f��̜'����H�ZN!� ��-A���G��=�"<�A�y���z	�Z`5%��5���F�e�.��>�l�2��p7��i�)1�,ɣm�Qݛf�|CS�2j<Gk��q�z�jf.�Gzt�W��=��h�}��Pq��ᤇ_�dTa�o���m`"=L������b29k&��B���>�P�N���S`��[}4�D�7���9P)�.�����?�.���qo�U�Ywx����rI�C�MJ��c��NO����4�F�^ތ��?.��a��/W�i@,��㳈q$�5���À�yY�+2p�������7�޿{ƣ��ʺ�K1Qlu@��!�<Ye$�Ӈ�zcΦ�cD������$�j�!t��I������n���Q$"$�Q��f���tH�L��J{�����mw��
��� �SMb<�ca�����Kȧ��z�{ܨ�w���#�\}�H�_w(#g�E�3@~>��y���g�E����Vʄ/T�hf>H\�u�5n�2x�ޘK	�4�&��2p�6W�4��òbw�1��4�����kXR��n^����)e�U��j�b�)����"�U�H7˩)��.3,:]c�P݂�[����7W)�}g��6�< }׽PϬv:C&5�&�����.t<�GX�d�5� �팭Z ���@�ع.�ػ��\����![O{�L|z�h:�S��J*��`�/��L_WM��L�i.����n�]�����k�,�t�M�@�Lʎ�eڮ�����ۜ��`*�v۝����uJ���8,�Qm����+C��{X���u�j3Y�'g!}�[����n9I�%L�35��h��Y{1wN�7h�諝t�����ZL�8,�#�ڀ���h���Ez�vQ3��Uu�}�[ Y3�XѴ�<�i�FAe�����.׬�(�{p�c���1*��D��@�AbrѼ���S�����Ec���(�a)�Wxvh�mj��tm�NK�e�S �I�%���I������_lϱj�[��!9Cn��"���h��q�=��U��F3r�&F��^B��;�	
�{3�,�3v�J�j`v7�N<�JmK<��r���Shm�j���ѹ��d��)\�
4�[�:�}���̆!Ղ�A�%էxuQH|e�+cwI��T��Sz��8S��ν�|kC��VvJ���I%Av���΂S}�NiN������I��ͭ�gh�㾽�O��P��(�H�fkZ����&�1�cm��wN*)�%q��CT
�k1��f��	�n�Z�IR&Xc�����ۦW.�P�AdE%�d�IXr��Ci�л�N�'	�ST^S�
,uJ��1�DA���P(°��o)��Ӎf��P�H�̤�5aPX,բ��Nf�1���&�Q�+��ݤ1�.�b�3E��Vژ�zq��S���y宀���U�uo�E�����pu�9�FM_�}�3ә��/@�Zx�ɒ?��	�juK�<E�-����<�G|�=HV/"}�Y��V�6j�
5:�6�J�(�4p��}1>6s��F��m�my{=L��߮=E����S_d-#�%tYl�!�+�����W>�Y�,���r(����}�Dܼ��y�v�wևмB-3;�(��XoWوI��6�O^���3�0�yP7B�|x��Ώt}h���󈊲�=�:N$�lA���Μ2|s�f:DyQfF�Mp�m�q/���E$T����c�Zz}�j	���U�\�_g�'چ�C���P;*h��"{cƨ�;��e4K� ���.B��?�åN[��˓�V��ee�]�ݑ�qڧ�v�V7�m��Z���D�.읃����~|Tv�x�ye/~D����;`Fq�P�B6���6����g�>__@��'N�EFM�YiK�~�fJ�1�L�H���D��4��`����n#��x��Ԫ�?4Ι>(G�GRd�%�hK��:��f.tx���"(T��O���֘ށ�e7�R���l�Aw���zC_��O�^�����;c�kי��I��~\u�!ˏ��C��	a��"�nΉԈ���C<�y�ˍ�-g�M���h�k�Dh��=�9V ��xѽ[K4Fm@�Xw�y�EO���D�>��%�9�����5�߲Z���߿9P�Î�@f��-�����w��-��V��A�DU\�\q��NrXZ�%wܭ*3P��f�M���#+xPUF��L�����;SW���D�d��=�%���i���3�dJސ��s���oq��+��	i�/0�r���ف��9�����=���yI�Ҿ��h�3���F�Kqd�U�g�+o+x�XG}�Y�.e@Қ�@�o�\.����38i� ��ś���p�&��	�&���ޡ�O��^�a�D�H��!֤�#o�u��#�Y<w=CG�9��BL�"��*6%���$ {����h�U8�*��7�0v����F�"�3PL�{����4��q=P{W�>�?}c���&���3��+|���_�$�1��@�4�\�X������YX�{o�y�@~����zZ�z7Ʉ�mb1eL1���R���P��5@���}Vt6��N�fW݈�1��;�~�"��&P�K���o�ߍ�L
�Y��$';� b��	�~Tu�8<d�y�.KY�x���A����D5��b���桚���R�z#��Q�h�&:,���� z}"��LlGz&MO���e��܅���Q&�儘o�>��ONj+(��k��'=�g;�Q�D,��6�X��uZ���t�ف��:,�>�5�ఢ��;�NT���'�N%x����!��3�y��%2M���Y����H���ز�̒w���(�'Z5�9�w�j�&�o�?��*Í�*�ڼd4@�L�Op]1���*L�W�^�����x�+�������Xi�]DzL*�z���I�X��(��e�eŅp�:ڋ�v�a�[�rܭ�6G.����m��3�j��F��M�u�3���2t����[t��`a��cP'�ZF��ܠ���gE�Z��f1��Y��F5���,jò��C<����}��^�$�.�gI6�H:J̐�I��iT���������e��#�Q��t�,�w�>C��
1yBg&_�����Vd�2|_-0}�flq�&���2x��ު]|"�+����0��M�t���"��q�o����C��k�\
}Ad:Zp�&,��edc�&&}�{0���������qg�+2c:k�*��^/�|��n�'ҳ�}�m��"�3-	<l��3'u�ٕ��yn�備�FCo�
�L�_�M���ľ��1�ʼ`�r=�0�G��L[֧/n���\�U���!��k�5qQ}y-�4����=�n���GL_�$��鳻q�4��@��wX��2��o��Y���8�F��Q�㤜7��>�f`ӽmVb4�'�alq�!�A�$�^(#�deȞ���0z=wn��p0�ޏK��{���`*8F]9�ygd�Ϋ�ne�2^�,���B�����:�	d٧�Tn�����|dՠ�NDyQQ���^,�؄`yc"�C��s���r^:>"H��R}*�3��v��d�Qi��'sG�x��<l��q1Ə��GNo@~��(O��WO*@⣞Ax{g��m*����%�z��1D��7P9�]S2�ɓ�hΓ�9!��fXUd��ޒ��#�.:���.��eţq<;�6��F���.v4�9�SS��3V撞�'"��U��M����>�����D�<|`�5ő�;c_��=����F��gi���* ��}��Ӏ����Y�\љ�A}�~Q7X������џ�^W�uifF�hOEzj���5�
�J���OT҃�Dy��B�3&ukS��{�ʅ^�ΓZ��#��j/#	�7+M�ކc=G�3�N��0Ƙ/�p2y��)i���s�v��Q��H�t���mƖx�'Z�K�di�i􍟔z4���B���]{��/b���dBy�hv�He�%҂��Ua��ݻ����t��̂=�����',�q�t�@���W��j<�*�<}�4RcBn������;�ϲ�V�F����?YP0�Xҕ{}�*�K�|�*���P����->��H�_��l�!~Cax�BR�e�,�z�3�n�޾��dȆ�gH�Zp���D@��bjnmI{��Ş�@��k�r�3�*�p0��Q��[�w�i�Ä� �/ i�4�6��{+<����0ߪ�[�Ҭ�q|o
���*/�m�GL:w2F%���3o�B�e�B�Vt�ˈ=� VGHN�����;�^΋�y��E��N��J�<oU�k�KY�"}go��m�������Qf>�8O������@�|�)~ݗg���4�<��.c��B�5hx�&[�:�8�;���v�c�߾q�@���u	�i�q$D|=/؏
����^t�t�������$����¼�Ksj�vݹ�m�}i^AϸTM��}��e�����yS�6ʅ�bnk?9�����g�_�R4�V|h��Ό�H�ϕ��^�����esPalx��3|�lǤG�,�C�Jg�s�U˸E�Q�0�����>0q-k��ZF�&_l���M����#a=y�
ȏ���@���@ݾ�#�c�z:H��x%��;P�Ebnؘ�G��X�5�ewWQ��	|`G���:����H���a��vy��q�z�a�C�ǎ��GI;��Cua�f�wg][��e�(��=�ƀ/��P�
�PӠ�L��FmvCSwm�� �끒�Z�2t�"hƭ��y���4�ʀ�Y� �=}bWb��Zr
�S������21�����4�7>9��>�cr�3Br�K5��-�_`����G�B3j�۹�Ы�Ӹ�6���xRO�����X����Q�i���U�f�+9�7�����:0�:}��=p+\}bS!ڣ���"�3WB���cfR~�$a�q�śkb�/mȺ��lW����=y|$��	�ܤ�9/�7P��6Y� �,5ɞ�	�謼�\l����㲆Z�+�K[�H��9�=]�޽��f��|6�G�ʸ�O��N���6�C>p��]�ƌ�'��ZF�$��Q��餰ĭ?���|t�Ύ�MZ�:m��$��G�yd#.Nϥ�W��cg��q�\adrRY_y���0��!�sj�*�W}�H���kM ��=ȜiŰH����׹f=)A�Qg�74�������G��6h�z�S��C�
���d��Ч���A��j�S�͡w0Ωt���,���"i1�	]�lF骃zܸ�@e�x��h�y��ײ����I�^.�[(Z�FN����t�&�J^�WNR��9�yK��5[�%w]�&��lC�����I�X���f�6�WcP�L/��r3���ftK8j2�p��vY�p+=�>RL8��H�J+��H}sd7f�o`�n���i	ʲ�k��\u��aӭ$3� �GgۮJ�Z�e6�jӘ��(1�got�KΠ�*S�����P�����J�2��構E0$ԫMSp�EZ�Wwő6�����^MA�r���M��aW���uv�L��1o7S$��I��F�jE�<���w4��<;6$Vs
�9P�|�67�:��Y�lX F����b�eByw�������r9��)!�6��8Ǖ�w�J��在�L�\�T�H2�;c�k�O�+U��.K��:���I�:3>t%ά�C��\�I��Uf|���x����h/��we�;ȕ��9I�m
�q�jf�D�e�9��&u=p�l�7�:��w�f����zulH�I�,�܇�j�T��т��UM�Qw^|�-����\r)+�Fқo��u��pJ7�C��7B�V�`/��\��֯:��:��z�J�}��V�_v��w��ԛ%vQ�8ANNjs2w'��;4ro�-ËC0���w\뎼t�׺gDX�j�;!*Z:J�[U�:'M٤�Yì�*T%kW5E5i��
±
��e*��
���`VE�c+$�a1�v�,�1
�N�*H"2� �R �4�H[I���	11��&�M"�]�)!���b�"����i�c&�b�,Rp�Lf2�Y����`i�����zv��X���f���F5��s3�e.#<tNh' /+_��}|r��Na�S�~�:<�Q��؁�x�^��]��"���)*�兙�zdu�I"c�<Ovdi����cH��c�"&�\L3F|��:c�ݣ�[��V�/���tq�'^��Q(a�-";���<��{��p*:<Iæ�RrGGjȹ���1���*^�l�4�4G�QOtZ��c}"�"���]m��y}�>��Q�1���f|�T�ZY���{�S7�W71띏p�|��hq�ށ%꒏42��0^�������i�q�N�D�!��s�<d�&y�3��4z�.�3}�I�zN�d%�웈$��^/j��/����6@R��$׺����7�˖����fB��T$(�>;W�oD&��'C�{�ᖩ�)��=��,�e�I�{`n/6<��/@f��d�������)�^�U�]D��&�}A�$s�=A�횐�|�Δ�Ok��0h��#�k\x�ˆI㥒k�=�;a�^A;���P���Y�B�ІŹ�N���
�c��^������c��������
���~c���� ���Hzˁ ��m=�M�*��L�w_UG�W�Om���:G��L�>pȗ� +�C����{��r�ܯ�ɣ'���D�T��n�OZe�RF��mZ�R
މ������r;ș���&����c��z���߷�x\������_н�Ν8. W��qs�+RY��𪬾A����hƻ�m�Ω��+�Gṡ0,�ucU�#��+cb�b<!�$n�F�󾼠�=ŷVI��_�u4Qf���\���<D,Յ�����Ȝ���L׻Oj���,V ��Ĭ8|��;~�!6"=W���Ye�&���ZE]C"���7$�Gm�w۹o|���=]F}�E�q�!{�a�A�#N6�����G|��$Z��̩s��8%af}�8Nzߕ�x�u��a�<��0���x�R}Hj��q����f�,�N����"yqx�:�b��W��w��.�M���e����<~�=��\}��(Y�"lB���B}AK}�;W���F��H,��#�4W؆[���Q�:E�y���}���$U�ܸ�������_xDZ�N��3S��4M-�CB}z��6����pB�.���Zˎw]�Fw_޾�K��΃R���;��"^��r���t�dB:I��AF94Ű�Byۮ��B|��B%A�\ԋZI�L
:N ui&(O�5㩽#Hf��.S=���R)3�NhɁ��~���@[�*2d�=�ħ�Nlq��
ʭ�so�&視��fG*�#� 5�3�i��t�J�����A�H�ؼGZ��L����?Id9U��w�r^����VMOQd�\@��H�m3Ŗl��#�܋:| �����~WH3�������,>~��9;ѵ����E��� C����ki~�>;�fzk^��v�B�y�y��N�3"%��Nˏ�7��`.~�؏]؝䢏uã:-��,do�Ϙ��'��| ���&���A����4�	�Wq:�nʾ���_]�{O"���(�Wg�`YݘZw/�����-o�m�i��#=p�$ٙ�p��>��W�]���S:C��$�JA�H�5��l�{��r� ������fR�Rf=��j�^��at��X�{?CHϓ�Lі]��Ĝ���`����z���|dɣ��u�@�%d�֧�1���v�:T7;un��f�3�H�g��r���>�U�P��^��I��Z����Ob�"P�hϓ�ki@����s���X{>�:��C;�'��P`�!�'�F���;�Tj���ʶ8S�jjGF�`v�!��񖬋g�7����7}�նy�KC�Z�B���qz��@��Y3^�������ܹ�v�SszA�&��KU�@Uh��M�h��2��R��X^�k�`��ݝ�PǦ�Ҏ������ ����f�ب£�3���q�%Y��r}?q��M>��43�ϡ
�+ށ��(�ߜ��yyJRc�޾���r�Z�q�'H�MJń�7+Mߵ7ީ�����qQ��=���w��s���3��٘n���s�L�q����ڣ���{#M�	��{?_����[RI�R|u� �����v�YǕX�<��_���Q� �nD�̂7�ǎ�2�x�d�`ܖn|]߰��b�Dy5	����!F�2��(����8|��D��C�"���^*�(�G]p����UEթx�bĄ=�<��.>äm+���	TE�[��]v��y���r�"�#&\����iz�q�ڼQ��C��%��`6<�5}�T��f�N�b��[%<�3��p��9�-SP}ˈ����������q6���e�U�
J�X�[z��\<t1��ʕ�.�Ր;�3+��LZ�\d��q�
��k+�[�j�l�!6����ج�ӷ*}�����8�^�l//j��̚#���W*��x�(��<r+�n��د�3��T�r��F^�1+gZ��O��1k`Q㧚��Z�ڄ��dT��M���~����u�}K1Qg���3P���Z�ߺF�hY�F�6���9٭��d
k���R4���(�e�r���X��w���9Y��N�0�i���8ߪ�t�r���sWBv��3c~��g��N���ta�#h����aE���[�_��\A�{gݻudE���w��gz?��F����i+��q�g��ql�=�FE�����k�u�-��Q�ξ��+��(r'<���������T+#uq�T>��oN�/#��j����`�����l�y�wS7����>�A#��r��Me�0ګ�;ў�{�¢:r{b�M@f93�#:��Ȃ {`t�'[����z��EJ�t�*:I�>�t��Uz��ʔd���_Σ�M���$D�����:��L�i_�L��۟{ޟ)VE�{dD,2D�����lq�w~�eg�X[0gN�:��fH�C#e;W��n���4o��rd@�.���/��,�K���-f#�I_V\�����*8�pB[��kE̼4\նz�.R�ɠ��dŔ�uw=��d��q�i��&�ˁ�� �+�3�W%W��F�f��fZ�ƈͧ#D����̓�MD>�L��1�dfȭL͸w��y3��`��{�M�0sP��"���};5qQ~�3����Y0�ݽ�AⓏ�I��M�ȃ/:p�\x�y#{ѓ�=1����TY�ZԊL�q~�H�fHQ��l{ia�u�x��س	W!!l3�<�Hp$�K�(A�R����3�5Č�-3>	��3~L�ڴ$�t}���I�*��D^��щ{�-3FC_!>�'`n"uw���|H���F�>�7+�4�P���L�H�{�O�8����y<8�D��<p�l��5�~��Mes��D��=��������%YfQ��g@6��{!�sL�rgܩiK:0ֱ@����!�EؽF�l��JR��cmM��*b���8��Q�=ˍ�!�2DRba�>�\�?^[�,8w���-?tq���(g�Ă
[oO��i�4�}|��Ӝ��9C��qdL����^Ղ����Z����de�A��x�C_�I;sw���F<i�>8��!}�p2����z�+�=�3��y���;�p�*�Ãށ�����9��}�O?_�0x�/5wC"I3H{=Ƨ��e��w����w�Ⱥ�H���1�r4�KO�IQ��ˌ���!x��B����-.����4|�/�{���=:6~Q��)v*!�EH�����ΰ����y@��*zR�UUUU~�[	!$$r���!$$���%�XI	!'p�?X��w�C0�,�.�B����O-��|C]�Ivz�0��Jk����g
 @ ��B@�	!&�I ���B�C�xFf�Bl,��C���BO`�|^P:�|����yo��$�ܞ����v֢a�7�願zH!���Rs?�t,9�a��h�u��|�d0���;��s�xI	!'��?�����?�!�y �BO�D$��BO�'�XY0����I�C�?�!���$�w)��2t��������{g�|�#Ow�	!$$�?�'���ޑb}���:��p`��|`S���4�z�Y�~e�$��Mj�3�D7���4�w��*Ώ���ǀN%�����d$���뷳uˇ���5��! K�}�C$�@� H{���V@��
ag����2}?]�Bz����?MϮBHI�	8DI}'�'����i��������YԛT��zD��sP���~$��B���?q�i���<}�� I!&�P��c�=a�!<�����{�d���pjS�'����;��9~����=�{��<�l'�xyt'�<fxB}>��������BHI�Oh�����b����@�t�)�2Rv�O�g���!$�l�$������M~h��� �I���C��Cp�����I	8	��*��;��H3� �S�I$���&�Ò$���	�5�u3��Fq��Y}����d'J}da�-���ٮ�!Ɂ�F�$$��f����_bC�	�BHH�~'�C��g�||�=�'���?|�v�< �!؞���'��@>_	�'���}H������|�wX}���O����>��9�����$����|��G��!������~Н �!$$��O�a����?Y?Ru�s��b|����y�0�	�����ܜ�8$ ���р�0�>�>^(��|�����>D�D>��z���i�	�:�y����;	!$$���@�|���OB9<o�G�'��Q<�P��	���(��9��}}��!C�&��y=L� HI�0�a��󓠐G�Y������	$$��{��S�qo���7��C���9��>y�8!�Db�A?̤�˿�!��s?�]��BA-�