BZh91AY&SYx��ժ_�`pc����ߠ����b7��  ����$Q�UP���-�kj�M�+A��I(J�@cd��"�i�R�m�l�٪"�� e��SA�`���Ѐ�}�UD話��6l�j�f-e����l+Z�T��V�ԁC%df�[j��U��)�ҙ��5lP2�mFl5%4�uՆZib�)�Vֵ�J��2�",i5bIm�ZYa�Me�M�f��ڋ2$6�6i-�f�"[j���6*��0	Y�kVʚ�-��[nwv�J*-��p ���ѕj �T�j���t�S���!�n�D+\�n�;gmN��ݮ�Y6Z��Z�[:Ewu)��[i#q����:^�՘�[aeT�TZŶm���  o|:䭻�W���vs���)�/Yk)����Wg��K9��԰avg��mb������N��anO\�մ4n��=m�/m��n=��m�R�+ry�"͂�J��Ŷ)�  �}'V�i�zR�$L�O�����}7ܓ�T�[c[i��Ϗ|�����W�zI]zr�k�O}z�l�IO��}���Y󳲷>��+��eE%��\�����*�o{*͢�"���D��+Q� s�Ӷ�6ك��{OT����޲���UE%=��W�ݴ����{g=KmR��<��[cJ�{��;6�v6�u�j�ҰẊ�fu{�^�M�8�ڛ��6k`i��hk6���Z�� ���m�TT׽�wxҶ�J�ގ;���omN�x���MU�6�=�¦keM�{����5{j��+�S�֚c^����m�����93��E�n�^򪼫P�\%�f�mkM��kL��JS� ���)'N��Z��9�Wm����Mm�h����vw0�(�{[�<�g��)c��׭4yە��=⧫-���{ou�J�=����j%k�ܼ�{ލ�m�����m� m66je�@[�d��UV�>U�O[vݥ��ޥ�U�Է��\��ʒ���ͽ�Jm�[KW�g�B����׹��M�;2��R�S��ݪ��P={�k�zU���+6���Z�[(e�ѭ��������w�kM���zE{��꺠��p�)ݺw��5�]����ZG^ǎCT���sҊ�X��Ӫ��H֢���E2ڵ�+T�� ����ӪW����EޯOz�Q+Z�<�x����'�^�q��Uzh<��p=t��x��^�t{���(�^��=
U$�{5fbF�T��J٢�)U� ����^�oN�(%�	����ۼF��{8{�Z<�k�A�����뮕Gr�==� �{7Q�@�{ǁ�G�  t     50T�I4 4     Oi��Pd  hd   E=��MS@M=L�� #ML�5S� IT� 	�&`	�O U$�M�a11�C'��A���ST�F�h ʛF���j0�i�=�/���|�j��}�=s_@�*�/0�k��N���޽u����Wϟ�����f۝y����ٶm�����fٶ��a�m�x��߻�~�������o��������l�Y�<���˦��6��-�o�6��w�|߼��C~��Xo����m��������ۢ?qca�ɰ?y�df�0=��|�����[{-�=���lc�c��=�lɌ=����m�� �L��m��=�l�6���m�6��f�{&�{-��l�{&`�Y�{-��d1�d6ɱ���g�`{-�=��{#0�f=�͛�l6�[f���{,m�dd�{#oe�{&o$��oe����f�L{,�e���C{,��c|�7�f�F����[m�od��oe�{,���}u����G�ǯ}|��������9�8^a0�~�×4�J�Jfa%Öޢ�n����Õr]�\lh�JT�]��,�G0�A�P�U{Y�-�im`��-�7Eܕr�{���A@v�d�oK�����5�R[�h9.\����n��4f건�)�Ѽ��	����@lé+p�N�*�׃7��M���f!ra�IVU
��E�a�����9�A��ǵ�L�7O21����n%y��#[`��+���ek͢+���v�"�H�4��k.��t��jl�����)���Rr���)5�Զl;g~�ng�f����VC��PU������sX��}5�VRT��Ѷl�b���Qɹn���&t(�(*�H��yhޝ���h�m�	�,\�v���]��@��c:X�3�z�
��.��p2&�)�*avi�
V�+0ZȬ��i^ٖ&K�p�,���1�xɁj5�h]F�JA�Fe	p [yZ�k���r��c�{z�Oa*c�	�IO
.�e��i�T�n�����h�'X9������8`Lv��Aa"���{D�v4H��4#�.b�go7j)�yII�f<Qf��[�wp�XI��f�u��`����5Xd5oq�ǒ=�m��{����4�݁�c����^��
di�%��[SVc�M[�����w,�t��cp�;21A�R���s*[�D�ȵ��a-,:,�X��Eګ#n��8Ra[�#D�m��64�G�5R�՝�]�n��u���[�ۭ�-ݜ�x��Ca�^�����v�>�P���NK�"[cNi��|��ܶ�=�HӬE�n�j`ʏ^��ɴ��&E��n������lY-�)�d(h"�0;6o�CT&������(R����s'�j Zt��V��)m�WD�Y���m�|�ZBavi̵z1��73mY��6�|1�;�톎�;"����KO+i�/����M���n�e�q�:�*��K	�V諀��0C����d�۫vpH�����Gb��7u��1㩑�©1��ɍ��4�n�I�Y���/^�0�Kgin�J���`Jt��kH��FXh-9g�3LRx�8�ĭ&I7b�ڌ��n3H�w��n!SV��0�&�7���Xv��7+�w�6�V]#r�$�gGr�(�e����׌u+Оi�Z$�2��F�u"�ҭ��,%w���V��Q��5�&�M��/M�{�VDK	G�5U�P5YI�!Y���-���ن)/4��YFY]�J�ʫe�
AuVn[�2@@Q�V�J��1Z� �^�m�-��u0YL�]�IAz�ٳ�ֳ��a�$f|JP�xlI�(�J�inJf�SaÔ-v�)Zzx�}[�sǃl]_u�U�&�FsV^��Tk)9v%��� ��� M���h���!�]�͡+bxC�6)��I3*��7[�wA�4�Ch�p�wWK�Z*�13�yJ��<X�t:�nsx�/Z��Vp	�lQsb�́���œ�/�x�̕f��K�6Mfka��vޘoi���"T�Tꀖ�����h�VÔ�0y��F���e[�|ʼ��R�s�ؽ�:Z+(�ga�"`zNˢ�Gb��U�:�m��w3�[̄��M�4VnF�ضL�-���2&-�&�&w)Zl��b	Fiw���R�f����r�ʕ�O����Z�eYr鰎�ƫ��ݤEL�g�7*t/p�6�ٹ�A������Ú�W3I�0QSq=���#���B67��3��X���i�Y!���im#B��WX�Y �hVD�Z�94��:�ef4�n�\F��eU��iea6��n���o��Z:6����.Y�-��f٬�b�[�F� �T�T*f��p��P�N��_�e�mi9
�&L�?Ey�k�,�u�����V��V"�V�I�'7A�[Ɋ|���|y#�&����]��u�Nփ�����&�fM��(D.;l��[��&Ո�^@���(Zh�ʻ/(�pn�F띵���� �Į޽��جth����Uw��u��.a�kN[y-�k{��wݤ]�q��j̛KTN��.�Y6�b:0��F��	58n�K�S3 O]^ڲAF�n� Tw��^��Ӽ��E*���y�r�K��]�oK�7�t"w$�B՝	�8���I�vVC/5ݑ��Y?O�e;�sP����T�ݝ�,
�ێ�fT�e^̹Fi�^eIe�KZTݫx�ͬ�l��&��{SV�*�ϞX�{LcW��sa�d]���\�Iy����c^رV�*}�ե�UcDWg&�=ǖF�P�lK:���.�<�-3�*�&ȉr�f�Y��Y��A��y[���O5�3q������f#/݈�˪?�e	��;�W�1x �Ͳ6ڗ��3�V�F�ő���+5Y�!���I*ԋr�� ����i����J8�HxKj�k֍�D^���y����9%�ך핫K��ƄjOp3L�@�@ԭ����l�t�M�dŦ��6�e�˫�ǘ��ÙgJ�,M@����e] H�葆���&�p��{�R�X�d�@��	�fM�yYR�Oa��o j�Ee���:Ҡ���f`��b�T���j��0[)�RU[(Jj��B�E��Cp��1��̤fdi֕y�������4��Z�(L�d(�6�K1U%�2�u�ҵ��lqfE�I$�jl�X̫طE������s8���v��uZy�<�fEl�N<[{��0sE�5�1eBUHj�&�C�N�1�K�n^�O(Ԭ����nޭ���%l(����\ٶn�e�vaЉ����ڗ�o,,k�+���nI��NV����͔sI��&R��S�OAw�Kq
*� �xn[�H�L�H��N�F�e���S`$���Z��)����ae�?�
�cU�Z�4���-�Z��.J�e��f�b�od˅��^g'���S���CB�yt������#�2j��b��U�-�\��V�����7�V �	�6��٤�����U���.*��傍(���/�gl�2�R�Pb۽�K��z�Ϸ+1i,Z�U�WG_��^�n�����]�����q��*��׶��ue�+S��Vh͔���࿖���K��m7"&��.έ�V�m��Sn'e���ԭ��Bf��W������I@�A��	ڻ;+u�$6J����Kv����K���2�X�����C4S��0�T�&c��J�*��/���w�C�Oo1�C�!��c����F��y���7.�d1E�:��R
f�.�tԙ����j�<ð�
��dI�bݠɣp�4هf���\�p�ձ��9wյm�m��^\F�be�ږ�f����6Ӊ����̆�a[����a�J�B�H\@�̔ ��+�+�͚�8+kӹ�����$"W�^�j��c9[�q5���P�0P$n؎�L�[RJ��!X�Zq�S�&�%H��y�:�Fa�q�aQ�5d1D��W6��]�wIZ�g_��5޵#�h-mɕ	'r�n!ͥ�V���d�K�t��5ALF�ߚ���Z����� ����W�x�P{���� �V�*��3[WeJ̵�˄j�W�vX�u.����\+ph9v��Pbѹۈ�\��E�]�4g>�4�J�d�3����j̫��gd��J��R����2W��M6T{eb�����ݎ��|����Ü���*)`ⱴ��M�T%^�b�q��n��zG�]��rk�����%J&�
�:#��B���u�/a��S���ʑ\��M,k���Ȗґ�NP��t1⼅fD��
v�en��n�d��10ػ��!OsR�LCPz�]�(�E4�	�k�ձB���%:�X�j�_<����DR�7�. �+V�"�̍%�������������
R��I@㍧�jで�Q.��rt,�6��ڸ�a�+6�
<�ܷt���b�A4.12��P�*���Rd�"}u"�]e��f�Tj�h9���k u�c�wR��E�٭"��ua7Xs0�b����[psH��o&�y����4��Ŏ��.�<�ͧ+.�-l����Cٵѫ6�5�j7
�$[,���0֜Ƭ��3Q�a��5��}�6bR�TZ��i)q�l�XT��}�Z\��ۃ�6q'յ+�k.ܱgQw�`Q�g.H���(F�f�[�*�@�`���{���sO:y�v���v��Ÿ��,��m$2J`�H>r���˵R�[��ov�=���?�Y��,�g[�x��_�1v2f�hf��ر�5��	�mvr���嵂�k��R��Yo����h&�:;sX2�b��x
�6іJ��$S��J���I��J�0��b�����h:�*�'A�� �Z���d��@��q�H�}�X5�qgS��f��˭�n��ߡ�։� ��4iTZɸ��Md�N�%r���1-�L"�m�-qY�Hn�l�m�l�IT�D�H^��˨� ]/�[9F��>1�.��{z'�z�:/p�ƙ֪Iz��h���k	�\��d 1SR����E������V�WbI�7q:os�b[��$ƳG]f(�b	Z-6�@����e�^n�A���c�+�y��t��@�i`�o�u�Z�X9CD�53e�%��+��2��2�e����Y,n�V�S-�RS��ǲ�"h���X�p֐wcQ��e��EZ�[7[��`|D)A�B�<��ޅ��Ԇ�mc�u!�#i_��ުƘ��N� �oD;�b���((��5L1�u��C�������u+�N�ͼ�rjKrdѦs5Ҳ��J֋"��	m~Il��hf ��^��'b#��f�f�`�XJ=�`��V���C�ˤ���n�4�&PƱ�i*�ہ�Z%���"�t�YL�%�pmf�����Z�t��=t(�X4U�3i2l}�(��aP�hi*�U�cF��E<��e����Z6N4�U^�U)���B�4��R�U�kh$ƠvA�yPd�t���B35ˎcWt@͢cm9s\Lmh�%*��q�a�6$Z�����j�<����řQ3�75
i(��Ya���ͻ�Q圭��lђ��[��!/C����CFk�fː���j�ݹa6vX+�8��+�K*kR��4Sym�".��tN�Ә���0�7aڸ�oS˽���6���������r�yz�9T�AH�Թ�1�rɻ�����V`el�`����ٔi��T2��'N��7�
n����J�9%���Yc
�q�[Ytv�[ �w�a��+/7%�.]6Û�r�;�y.���ⵁ�ԠhJ$e�r�?\̒,L
��v���Das.�ӶSy�:�V��/i�\X3��w�OKoA�Ov:��#��Kt�q��V��\�f
G6Ճd��]ۛfY{�VU�����pm�6�{R[�-mGN���f͹�\"������?������N��Ct*ۤ��'�F�`^�� � "�m�W�-��%<D�EY��H����V2�
�#����D����vw�n��p�)�4y/6	ko+$�-Ǳ4��`�1~� �;?6s2A$Q�����J��sM���- �f�^�����{[�REK�����R��[�;���wz���I3��-bkV��#A	B�#��
Y�3	�7BY8B�B��o74���9�Sw.+��cX)�'DF^Z�P
�5+:�s�d݀v`&�6�ŸdI�d7�A-p@��.\Wa�k2�*���r�NL�0(�1i��g.��puI^�0��NPt�A�n�B�Y����6fd&�d�L-$i˔Y��F�Vf�Dk͛�D޻I4o,��ІIe���ښ��X�pw�R�jM�Nfi4!���m٬��@����@d[7h\��liÔ��L��y|�b��q�HkM�2���]�"��{>���R˫��7iԥ�P̂������;�&���Mܷ��e��[b���&)J�QAZ�[R�$��y���{���hђʢ�v�@m��p`����K.��&�5���:�����V2L@�W]B��yƴ�4��V��=W���˽i�����)�C�X��MgM�b�Ive;�щ�p��Z\
��6T��_�b��n֌-V
6�0�K1����'��sI���J'3+d�.]Z4s#KIuh�b��Gk*��h�1�Mj�	�8M�[���a
m�$��d�"E����W���v�)�.�kz����Ù����lYh�j������� ��+��e�C��Y#��%[Ճ3��!XV��V`z���˦��P�H�]h:���mH%^ɇn���t�-�+5H�L�օ�	��:���;��,�T3V=���j�U֕���)#5N6�[�H0�� �S�fMxz��.L�ΤpǇAlH��M&�H��7q�Y��qH��I�䣌�6�*Q]
���ja"`�z"�Ռ�X��)D�L�j��iv�?-[���է��`y����;�췁V��,[ss%��F'5�n��)⫘aK[�b�
��-���E��ۛU���W��L3n� jN�m��k�� ^f�y�;Ur�I3K�YpIVN��su�.�l�uo�u�YfL��*k�La՝GGB�͊��6�LL����TrTa��1F�eY�A����Ugo�N3���Ez#kI�I�L6p�$�o�xB�G��;,�q�F����Ӥ�^6Qq���}p�~5�ii�r쵖�Y�D�.�d�4Y���4fqD��ZI��:ae�$�G�:��Mힸt��&6|_@XH9Jq���T�Eٖnk�lU�7d��p�|r������x��Җ�����]�m��B�pF���e7�kQ�������?�{�o}��#��_|�=��'���C�Mc�;�u�`P�ۚ��G_�յ��貜�����Y[г�j-��l�5�]���7�F΅n=�:����G�����u_N��]��k�͹������+x�&��E��ϯIt�r�W/����Y�̙CJK����l�=؉��ŵOHX>��2[Uǜ.�	��֑�e*tIT�2Hs�Stx6]�y]�6d?�t�G5�0&Ϊέ���m����m٬�OL��z]v������_�O�˵Y|uu��:������L���n� �����S̒���讙��oz��j�Md�o-�ڈ�5n�v~����Q��*��3���r�)�/H�m�)���d�Lob]���KP��Yrps��W��G��7p�DY������Ƕ5t��;�[Nk��P7��vpٙ38)�+e�r�����n�����G.f���+e��m[���4��&6>�rI�x�l,*�Y:GԮ�82:�R��D�<w@����z�S�z�^�T�������IQ����@X[m>ƶ��J'1>[�1{�#w���j�eeM��WY��k��8:Ո�w��#[�����-=igCouJ�Ӣ�˰�
z��eۙm�u����ݸwb��_��M`W�k3gU�b�ϳx���;����F�cB�a<3�C P�,e�n�uD�t+��C.�5�.�c9U�GmN��3o'5g`��+*�VUm�=��RKg ޝ�CU�%\��j�i-1��녮�j�����b�ځm����`P$l�x�;i�lƖ�p�K�)7%2�$�FX��v���X�F�)�W о��!&;�f�a�Cݦ�Q��e��a˦�_:*���17�����y�ͭ�nJ�.^�����z�3*I�X��k3�eƴ4�̵#�7�5���Y��,p<�9�r��t\[R'��7����u�<��҉:�-����6�rUw����z�|�C
ܢtJB�����V�ܚG}{:��1��!Q���a�G��Iwvz��m�રe8�oP_�91���I0���x�8V�j��'o�=������C�%����Tr�1vU���8�c;6�T:�؂���x�Ȩ�mEi:{ya4Flȁ���(/S�@í}��ջ�j��X��C�spS�+%�����3!}.R��3Mu=��/: Kd}��Lt�PS������+,��2�9�W!��4Zf�W�R!n��hSn�K�օ9]�2�)��ϡ�]����;K���O��Qb��c�c�(VP��T�E2S�N�$�h��#���J�|�j]|� d�5{�<nŰ��
Q��1ϗSͭ�rD��c-:9r<=eʙ�8�yG^������FwWv�L�mI/Oy*<A�$�1�%����J7�7��geeX�I����0H����;ݕE<�|���ĔP굶s_�1���r����lb�׋���Xc�BPv�o(�՛P���F�Ÿ-�AF�$��+�E����r,�����h�FCC6�-wG;�,yW�e�9��
,�� �"
�y���t�I��n�p^�L��Yn)����G5�]Up�`���d�ټq��v����y`���U�u岾]����N��7��<�L��f��1^�[�:�(0�P�<��f]\x�L�r�Ꝧ���ܸ��:k��p��˔1�z|��z�('xrfY��9˕h߀�[��9z�����#��I�����%�NB^�į���$@�qd���f[�V��C6t�J�[�Mz_t[rF�8��h7b쎗�e՜��n8�尘�z��A�2�G�AQvk���\6ۥ1���a`�s8����@����S��`���Gue�V��t���DE�K�l��m�p�o]�MQ��^G_�Jh����i�l�ܭ�m�B�{�}A��]fvn��J����R)�s4d��f����%N^q:����/���[��8�=S������KԘ�l�WVuNQ�:�ֶ�6a�j���7�h�h�ʁR�i��:/r�4��#ފ�F��Y�oh�EX��o&�.a�itQ��	�#WN�-Ǩ�Wq�E�:u
�r�������tn8��v�кp}dg@�˪pn��0��!�
��:�i��Ԇ�fÊ���P=2�����[��mC���1�^\�ԫ���cr�����VY�� w�۝���էa6�cE�Up%���y���醳S�o��K������儯n;�I�3-T���%6���"Ă���Ba�؂��-;\�c�ԧk����s��-�JӪ[콧7��cM�NM��,N�D���#)�Tp̬�t�θw����t���=�Tu�n�;�f�]��c�����3.�e�e����{7��;wC1���'���LDX�E߻C��ҵl-�ZٛZ/T��y�ݦ�p��ɛ/-��w7��5r�.�\B2�9�]��$�w)�*�$5��rGۻr�wWv��8Na=ψ�	B�f�3O�Du�v�f`X�u)�<�W��uhR���2�� =n�YjJ(q�
�2u^�,1�mj��j�l�(��D�<�ln5#�o-C����4�m�a�m�/9�Wu�tOL�7ۋX�����T�Y��Y��kԬT)H̽x��>�N߬7/��׵�f̍a�^S�B�+okm��g6SVP�c�0�+/��R[N�i�6��󨽚�[DK��b�a����"����y�,ul�EBW��"��4�	e|R�r��Rn�uP���˧-�o�Q�?.]�e
��gʁO�����)Yݷ�x(��]-P�R����=��y�_@n�|��P4���2�m��}(��t���/I���C1g$�Ⱥ-�B b���y���|*�9�k�"��][W���0EX^�1q ��������l�o6{��s�1eM��:�����h�Ʋ�\ȋ2`9NEv{��-�6�6����7���w�;�'�˒ ���ӈ�{9����'t.�nnz-W9. s:��^�W�S�y϶�m��iH��RO�4��� �-Y�����Z�٦j�[���6-�B��:�GWd�v]�E��m_^�2H�7ի��mZ����/M��՗Z�FfVfU�,��rV1CJ��p�k�h4�n�9�R�Y6��Yֳ���Q�C��ƽ��)���uŻ�ث]��k.�)K��ChI�X�
���f�Rv� ��C"a�K���׸�K�g'�,�b���Ǐ�5�5"�Tr�#�d��Vrhf�3K�eR�t�e��ə��ZD��9�nj�ķ�����Ϋ|�ǗG��u�D�V�kO�g,����{����@n�8�� V�*�MQ!�j0v�5}iا���Vn���e8ݧ�л�T�,=��N�|e��R(1i��J5eac&���c%t���ނ>M��Nm^V��άv�Bn���{��Z5gvf�Z"�Z46��(IlX��nU�zֺX�K�3j}s΋��X�{l�G���VS�J�0�����h=�Ou�)Xz�VJ��,($G���`w���tT��!J�&k��QT��jk]yw�R���6�"q*�3[Q|o�S�:3���Ď�$��i~���yx�㛯�rh���e �m�`�Jm(9E���HM?��/�]�:�W�]�A��'(k"PL�Cے�"��LL��8�.C����n�\�#��G��a�y���e��Y���L�%vXߕn�r&j��c��X��h6Ld;2�C��M�Y�b�y�ƾ�%\��+��H�h��ݙ���V���q��`#�mf���Ն�:"3��0��g�U����k0)j�L�Z�n�s��u�qZ�X/I���Ǒ_LY�����P|,≽���vͫ��l���Ʋ��Jf�iZ�2��E�(:tnhv���c�=��	�e���Əp0�d��0��b�3劳��^P�g�}�Y7ӳ����]�m�Kn糃��Ц+4�U�)�[�ZW��/��B��n���.���	C�^q����f�@��"���W�/��U��lޗ.����ҟז�w���=����f�l��}�䦅Êcr�����67-���[ɪ^�p�W׹S�(�<�W�<y)Ȍt�9Pj�]l��dKJzx=���I��!bї}v)���p��}:�nus����7`�T�ޜG��Ã��V&ѻ�V�qD������s�[y�w^�^�͢�Pu�q3S,1]<��G/{].pIv�ha�OQ�]7fŖ��#���*�|��I^�V�<.j������!*�c'&4��ۡ��,�*�N���[�)����B+	�����/A�6�l�ᨘ�1/0�-l��m��;U2��n],PP�z��Is�F��ꂁV���n"�>V�-��Z�_K4�+�Ɇ53�ul��t�G������y٘,���_i���t��]W2^��Bڥ�u��q���`ϷhwQ���6�����ܞn���X-�xSlEK6�Q�r�S��G�[�k��+P��3w��ԗ^�5ʵ�{Yo6٭��3��K�t4�Kv�ے�����I
���rK/A5�⃦��0h�C�j��{�x��."�B�=�7���>)���tv�޵ˡ���g+n�򐭫Dޗd��:�R�U��ڱ��4�f��6���沗Ɣ��ۘ�����0�FEM	^�*v��hKk�<u{ǌ%r�[�i��]�n��T��%������հ�o�[{:oa{��5���]����R*���n�y��e��3z���] �϶d́V�I�y��iKc���s)*ʽ�,�Tŷ2��A��_,������^a�+tӼ��tM����bo,V#]��� N�JH�T	��Y����#;GT�ё�W^�q��h�_&]P�ʻ�&U�u��f[���1n�̠�k��N���
Ɔ�)b�4NP��3wV��H}e�һ�|���7��5���J�]T{�K�P�Q�X��+p�%���l`���gb��ҳ2� �'���vR������k�<��UqͥG��aX��{z��T��[���c�*e�.�l�nu�6#��zŧ�:>�@�dgq��lYݷ*����q�H���z,G5��m�ۖ�f��\�Y���S�s����P�k���ӳ�@/��V+^�x/�������v�|7/�׷cCl��.q��+��\��t	ݶ膙ݚ�Mٰ�J�rf�]v���xq��kD"JRӻ�*�i(W^�Kc��)�,\��v�f�n�4&ַ�����嫓�Kj�%�N��'3i�M#��V��y��a��T� �T ���5�����W]Y����[ޙ��)0_<<s$�st��G�ٖ�8�S�J���s%"���f�`+W� ��V-�� �
�[sMMw
3�g+;��̖ݤ��f��t��'vڭ�jd�M\/ot��o�V�M��Y�S����:]�����z����m�x;{��:�P��p c�z
�M2lV`�%fnޭO���:\�,�iid�X��8�$i]��I�+�ӏ.������0���P�3Ɗ�08nb�S(�a�TD4�"d���w���8P�*v�2r�'P��ʀO�b�s:f��I�a�*�q����-3ʭAL��[1G�X�Z����K���[5�ir��)�"ΔM�z���4N���D����F��P}���'J�Y�r����ѹ��d������vR=!��6fw9y�ݚڭ����(n��������"B�4��ae�KÐ�d���7�ܐ����I�N���&��F�[W�(��s��#_%��icf�N1Q���WZ�!�ϋ�w�G2n��4�����LoV�c�+��Z�����u���o$o	rmKqTZJ��|�� �W��oϹl�Pۭ���Z��p�nc���.�N�ݸ�R�Y	��۔���oZ앍��8u8*��xV�.�X�m�O�74��3��aipK��YmM�������%֗�w���W�Kc&b0n�q�y�D�6�T-t�'��ݴ�7�T�H���ھ�vc"c��B��˅U�b8���N���|2#�$�wH���VY�)˷h��l'����[��8W�ɲ�)V���:�9�����'
/�4��4��k�����<��fՊ,���9"o�u%N�0rxZ\��t�
��P�cI��e��5�O�o�07b��u��D�4M��o_���ѥJL8���ڹ�-�%�X{�:�x�{|��vIr�1ٱ�^� }��s9�31�����+'M"s%���Q55Ρidf�L nYCf�^�Y-�ͪ�*��5��\��+z.�O<!��(6zM�VtX�C�X	}�C4f�1��"x�h�;�Х�u"ût-��85يΕ�h��:�ڶ�s�LDI�C��ٙ��FB�]�y8Xa�W�r����:&�Y��M�FD��(�5�4I2*�c�T�O_?���[�U9�Q��%��:����wiY�P�j��/r�|�wf_I��C�q�����nM�v:��_h�s�{�1�'�IG�~�%�2-�2��]V̤̜v��f2�9-	چ&fd����J]; �onm਌����� �w���?Y��WP�Mv�Y������=8��F6��'^CYi�:�nqи�-;nK���7�R�`X�%+�I(�/d��SfI+g#�/��$�.M�$�$3���d�I9G:I��*t���C:js[89���ZRK�oc�G'l
�*��;�V�U��ǲԔ;'D���G�,a�rI$�I$�I$�I$�I$�I
����<�
 @ �$�A���n��7O�G^^����U�N$��8�|��<��7ź�~D6�bgMЁ�����,Ԉ�jv��:��n��oO.�<I���o噳�����^�-�ϯ����y�g�lf�m�������}ߊ�y���}���������:���&��}��4[���Ϻ��dl]�1\��h[!Wsj��wNb�To���,�-꾶r�l��d/d�=��QMS�}y�1���6&	C�٤�M>ٷ��`���*�f��uךM�+v=1���δ-o8�*��u31��.5���<�_>�f˫G*&@TM<��U����>�z;���B�Fޫ�[�y��v�&WDw9��"zN�M+"w��ǣ�7+W|5��0��g�����L��O!�{K^�G��[6u[�3��3K�3�3ƚ'(nEY�K-�0A���$�"��3��ҋ�|���f���6��mT(�t�$��	'��b�ȃ����h0�X��.�>�q��fU�w2��,̣��G�%z���&�ǲ��Y�)��/��b-����+-t���r̚��%<K�{��hͻ��(u)�5��r7���0�q�lʼ���y�ҽ7�B�>���S�X�����ws`|��O6�UM�6,�n��BΜ%a�Cf��a5��g.���2�B0��1�iQ�ok
�o�R�V]hU�_<�oz=���7�,�J���31,��A\r��Gn��X�M0tgb���Cp������1l������l0(�0�tf_n��®9'��1�!"�ͅM�%�GC�MW���&����G�H0(�v�
� ��	wW�u&U'���oFƼ+t�a͢6ZN�@�7j��iA�a4���'Z/�&ܹ�!0
:�n�&�3&�P�ed�@־[�u�SO�=Y]n�1Y�����й[R�ɐ�+�W��|AW.
�9�:�`��D���wߴ���ۻ9��t�C ����l�mn�O98f�[A�m��w\�����e�Ϯ�蔆�����e1:bǨp�f�����J��QdI{�l���6fǱ,�Ac��\��U*D*Q�F��9dL�rsF1�jf
{W,�ܫ��v��)��޻W:�Lm�խ�҃�9�PD'�D�/x�N�5P1R���+w�gr�}/,�*L��[���GM�gb��1��˧P���kx%����j���T�t��:�'I��QE�P֧�N�d���,�	��̈́/ <�k�I�j�u����:Ln�}��,�<nīñ��=��P�� ��X�s�?�㔩�U#GmSUzv�d<zJ�%L����\E��^�*��r�o64�Y|�9�;Ffk$m����n�л9	ɼ�c��3���gP�*g>g���e�;�`�{��4fWK��-�+���'8��9��gz�G��nk�t��L���B��88N'��]5[�J�B+C���梬KH���V:���������d|����%8e�;����Q����/lZ�+)��OY�-�� �(��;:-|��vr�R�j�����f��u�	xa4	g�����dv��;��V���1����˹V2�=(����TH-��X/[�}TaeJ˼�Wgm�U���������c�%I���*qX.a�˟>7tk<�3[�ؠ#=$�� X�n
b�;܄e����R�u��lގ%�c��7���g�ŵ1w1Ѹ9��.����Ԡ7\�8�WA�/~��\�(�|��-��Yύ�7�����h��
�xp{Ӫ�Ȫ,��s����Ż�/1���j�����T��U�D�N����_����pBLm�4�����P7���FE�vV3YX%F ֢X��yBL��X���qy[`c�c���sP�P�� Ԣ떭�+gq;�Yd:�K�\�+q�q���ŐB0�Y�q*�sͫ:��e�1�(���zW7�M��$7e�;���|���9�nZ��r'�-�sAe%��c�
x���q�
Fۣ��{\�cÐ�U.���#�[�ٽ)�8í�}����QJ`���46���^:w��O�B%;� "N�-�����D��ڜw�)`RK�G������k]�Po9���	3���eơ������U��M��h�͂!ԭB��:���a�/���l#W���wkT��'�@��$Ztjn0�ə�:v~��t�f�	y¸���h�*�\��*!��vu�j�QG��Bٕ|��oB#�"���Y��
�����+Dr1䐫�N�Na��$���~�{�nav��:�W��3v�&�6R9/+/Q��=�o��ӽWI��}z����K !6�)�fW\��v@���G/���q$�.X/�I��8�M`k`ei�v�=��+\��5.�Iuלq�:ꝺ�V��8N�Q)v*�CT��[݃�E�2E�W���Ν��O(����vR��3(f*�'.鬽��v�pjr�An�j���1V���ņ�h����f��/�V���X,Ӛ^}��wHv`��k,N�d�s*����'���s,Q�٤�]�U��X�#�$ۣ��6��J��]C,�IACaY[WZ!s	�n��wc�7�	�ئ$'{�)��>��94>�YN�jfq�)�[�q����zi���SU��١P9PY�ѶnZ��<�Ǵʎ��}3S�q��՝8T�e-�ұ�����t�r[4E�\�<���j���\/i��c]���峨�Զm�"��{�lW��4�p�98ٶJ髶���7�*huu�x��/Ze���=bs1aQ��{V�:����h��&�H�)�;�ZAQ���h��K͓&Xa;=z��U�DɃT�V�P$
+�Y[n�qq�ԥpP���kLAɭ�˖Zxc�6$���|e��7t�J�L*e�{�.x�q��U�-�-޴t����^`��:3*�RI��h�����O��P�RK͔�J{n����Rhi� 2�Ghbђ��_*n��wxb���Zu8��fP�̗�^R|]5���F���x�M��f�ڤ(�FpWQǯ��Y������b���H�n��<c	�h�q7�p�m؇W�p��ɇ�&�EI��|N�1�JѲ>�->�}�`�w�J��LMZ��vu^���הr��H7w;3-I�����\�`3�v�k�B�
,g%��.�y��U��T��J��\G�Z���ec��6ڹÛJ��r�tZ�����yz;sp%�)�i8%@��N�UX]8�-��V�ǂ`5V���=����hu�\}�5ke��_uh���ҍ����G:Z!�`RǬJ[��ҭ���z�\����)]u�ǉY�Gl�`�ʝ�2݈�%�D�W;�i�]�{N�9���q6���%�9?$�\��:F�8s ���v=�DVR��aJR�̻:s��K��vզY\�g�ćv�k�#�o.��>{n�ͧ���� M�FÚpN0��9yXm�/�lP�*TwJ�Mvig�>��V�G,E���ök�}u
�Q�]9����%'y����8�!� �/����H��r"�fŐRØ�X\�-���-��[v��tY��X���8$�֔�{G�ut8�{�\��]%8��ƪ^�7]+�>�w�`9��ֶ�aj�[D�[�me�E�m��D����tR9N�&H�u�Tnů��;|�a������菣qq4��GWz��MṯP�����D�y�p�u��[�7��nVeaK%��VI�ă��:t�{U�t�.WhX���]R�\��{�*�ʷ-��v:Z�k��\T������d��N+�׋xh^v(TO�r�F-د:s�H��n`�j��fg
���X���'}7q�����Af�c�qi˽��n��O���J=v+qGx9!����!���P��c��:���ك!a�3�PR�6�dU˙ٍ���0i��@�M�]�0��le\sj"'u�j�����Z��S���}rR��I]b]ք�p�K[�|^mYF�[�)ņ�-�J�i��o"�:ٲ,�8u��@������S�FHp�z��[Ʒ���V�fR�U�f]�P�Si��D��g\qw9����b��Q�r�%y��I�Z���ʵ�aU��餯Yy�-[��n�$��J�*�1�ӕխz㔦�<��9���}+5M.�?]�P��{�:������n���E˙V�ӿ�&��&vH�2y�Ru_�0ɴ�]4*�9ΝP�%����G]H�L�?�w.�����zV�Yn(M�!̬��f��˂:4� O�(�վ;+i��.���]h�Z��[[N]K?j?+�k����%���em�Ҏ�ܜ+�"q`(�6:A~�cU�'�v՜U��lD��3���!Z�F�%7l��ݘ�v*�x%ƭ��?du^��O;�����Kzu�;S���4\z-�V���,�V+�8u!��{��ȍ��0�36�΍�̈(��&F ����!s2X<j��]���vk%��6��p.��C4GQ��k�N�u*lLc���ڋ���#v��{���T�(�XNB�"�{w�U���gR۳kr���./2�1Y���6�.a�wk;,��9}��Ge��S�]\�f\�y2�7�w>�Zn�h��Jt�%�Nl���w�Eܣ�
o��Co6fUM��wC��M�0�51k��V��3,ܮc���6��J�#�[j������t�P�76���R����5�ي6B�;R11�z%��-��޷y�o+�����r��!2��� b�VI�uι�9���7��Pd֥��p�Y�6�'+Hknus)�u䒊�X:U(�����;f���]��T�&����9]�$'E.9mc�U�́wC��
8���9,��^����yA恭7�F`:�&%�8�\Ӧ`��rW\}v0Q����^f�4(r���Uhr��n���:���2��"Jj��GP'r",��ff�[�6�T��.N�z w6��N�ee�e�Օ&�ж_H��kg^ɲƻ��zL&�O.+��rh�'�)1���Ykw�-�Ob�����{�֑�\��C坆-����v�
�U���bEkeF�jX��d<ȸ�5�j,z7/�8*�u��ЙK��[���aǘ47�� �y��?�_z�z8�+8�|R;/�V��cɔ �C�9Pa�4仐��7%��D�pG�R�c'92��\8�000�t��#^����"���A�&��+6Y�;�K�j��SYvКc
C�л1*e�$<���cZU�����3�&�|����z���{��^�}3"�k�6�����)�÷*QWjг��|4H��Xc//���V�}&Ҥ��x�E���
�W�5����x�(@�����,Xg�1�W��mr��A3�)�����)����Jm��A��-��s��C�J'v�AD��̄�Q^ar�j4�����E�B�o�ͽ%Y|�s����M��-u�9w>�v�W���z���tk�u�S��[�
�2]a���saֵR&g/�+lTr��{�@�`ئc��&�v.d=��:�^����0ɲ�����V�j�Kk�΄QXv����Ӽo�S�hf�iŭ�d{�oN��-�:�ܽ�/�q���-��� ӆe����::��j�uq��"D��j)�oBt/m5Y5��:���2]d�Y��]:6x���)%���ktu��<��3r�Y�C(5�,�'0�U�m�F"�ݍu�^R������X��9�so���O�_3�8!n"��,�'�Waw2n5�!N�z<m$~q�}]��,���\:�};���A|�=�^�_v�gheړ&v��co�!���]��~`Ջ��cy!2.\�f;�੮��b�we�<��]fj�Oh��B1�J�5��b^j���ͣ-��K(ET�8M���,�N�G��b��.GYhK���{�Jq5JS=�Y'�@�+긫j��Kn`�,"��,N��ɰ�1�}V l�CG_ܕb��V���Z��6M��X'v
J��"�y`�29a]-�C�t��%���p�E��Q�ev�����1d�e��e�;f^2�o3H����&�g�{{�N���z�>�p+y�%ݽ����
tf���ƃ��̩�Wc� �U�˼
i�B}Ք��2ܫow%AK{�;�r:�_7���/)���w���qW���L�E�'�t���ݣS0�]�>��jv�G����YIH��8�UZ����K�b�t.�ݲ����k��Nr��Lb��jZ"�
�f�Yj�It[�_t�ěb��j�ٮ �'oT�;x)��Ur�Cȵ�٥���V�BsE,	��[�n���]:Rd�$<t���S��K�gQ��^��9!�*Y�t�(����[�Q�Z��]o�G�sk2�[`ӟI���F�ZXޭ�ڰ�j�j�_F�u�-�0����r^f$/:���c��IΊm'�����Ɛ�%e��6TI9�ڢ�V�����:����5xO!�>�S*��m2�O)BF���-%�4&-�M�Tږ!G��i4E���C:�����p*c&�C���CT6-9��g2bF�"���P��k�vr-,��3��udc���,�tQ�f�oV�*��ګ����\�k/�*tMkY��N��[cuw��]��Ce䷱��ә���G/^.��Xb�}�Lj��n���C3�1i��w��%�"�-��swv�ԅP�}չ��%U�w��6J|�_��^�����v�я�`e푦�峇J:�(������Hp�έ�R6���p8����VΘ�6�>ܫ.ж�����[kuۣB��G[�hOĺ=;M��Bu�J+z�s���U^%�6Z�\b,��W��H��vģt�2�9)�m����s��V�
��j�����7(Z-⡏��W�Np;�!���`�,��{���m��S
�����P�庂��u��+��r2�O��V����{[�2�<��x�9���e�R�c��7n���,�U�+w��e�f:F��r(�	G�Y�r�O�6�����^�6���ﾯ��Y��?�����~G�">�����O���_���zy|���O�n�>#�v���@ B,�J�3F��ʿb�sն�`e�'p������,WX��u�ޥ��a�W\�ܩ�S���r.��<na�:����S�K%�����@h���s�N�5��Zc�K\�shh'���j����W�t��
��a����mr����"<E���Ԗ�+wZv�/�j}!���<�0��O�7�Y�`u�eD��|������VX�Idc�vLVu<j�)>���_)��p�42��e+�p�YU�r���|[�{�ZY:-
�3E�S5�K_3�s��|��*�T/��!�d�"�Y@5��y𡙕'
�;��c\&9:�cm�沶��lW���^�!�T�����J�.�kH�P)Y\�H��]f�fe\y׆L�r���ӄ�v�֪�����	K�/��Y5.K���[U�OD�Kz=�ս�y��Xî��Hn�ʺ}y+J<9񥗣m�q
l��d��{X�R���G��;)�Y`�e��$&c�3Ol\ݺ8+@�}U�Ze�������!Y4I�K���K\�$��gT46���N4��sZ��T9IJ^�+�[��ߘ��Y$R�#,�N��j��̷=}��f+��áI}]��Ö����p �J��J�kX͸ɥ�Ԋ�WAs�c�Y'NˌȦ�2q��H�ӾߩԬ�B�� a�(@� b-��AS�U���ݺ�:��p�e+H�9j)YB��T����g��I*��V�ը����qJ�R�j�%[R�)JR�R�(���UR�RV��Yո��9�U眨�Ij�J+K)Z�Z�U�e����*�K*���^yȪ˗
<�JҕR�O�ĕ���
SJ��,�"V��իQUZJ(��V���*�*�x��ʥ5oS��jۻ���nUR�ZZ�9�eZ��5*VV�����T�U�r��5���J�$�U+k�7$��U��J��T������/���|�<|�>w�8�9}إN
�^������,����^��)�:��o���7�U�mM(N������D/� ��T��_�U�wz���¯����m��u�|U�=$�F3w6�����rw���՜����*t��QӚ�����ͻ��kh�ݏ�-���x�������{���~��C=�T��s��S�z��o����@���?_vU�q�z���v����&{r}�/w��!c,�O_���br�Ҳr/F���j��6�{�WJ�=��}յ�n�'��F����p����G�tLC��NX۞���̥픝h�7��W]Nl��^����Wa.`��^{h8��ܡ��T��p73!�d�t��|��5<�{�l�%]���j���@�y�K��jw6�3hz,���%��<�<ײV��>����I�����C����W��m���ܰK�9R��z��#�&uzL�~�Wm�_�5���X��'�M��_�:(p����!C��-�:�|^�u���z6��;[��H�w-um�俑H��0o7b]��Ǘ�7pË*R]�3����Z3C�hy6������w���5�35�F�q�6�<Ħ�u9��5dnsg$W3W�Z�[K>p�W��-��o5�����q�#ų3ޗ����ѷ.��Q��1{>�뛻�s�o� ^������c��<�Ї���>��ς�r���uw��6����5?Fw�ߚ������ ��r�<Y�,�C������;�½睚�7�p��<�|���Q�����˽=���x�k��Y�U�;6��S0�H=��6=������%�qM����N��^ۼ���c����J�۸n�8d5�;SGk:���#������7��b��/G�����_��SX+x�����_���x���:}���:����nٵ��jL���X�~�%�o�����g���ߏ͏�����O��y�����㚞cu�rJ?R�yo�G�ay�{�7�{0��~j�9[G�xu0�a�y�Æ:۷N�y�Opc���:o�uo�8�t������;O���Y}X��]IY�D�Q�{y��8!Lm5�~o2��]�mH�%Z4۷p�D�ە�
�L\�,���m:�8�;.�2��_-.;JK2U�k���;1�{r��\���r�ESsg\���Wu��t��&#�9u��� F�b�����R~�۞����N{�~�k9������q��]�1����72z�gbS�x�w˟�����?-�������;.��{��������ӟ7���'�Ϊ� �^�����UzOJ>>�k�s���%��חƩ����}q���f?FO0��m�;�ݲ� p$�h�k��!Ɔ�6U͛%��4���jl��W�ch:}�ۈ�Ժ�_��;V2?i�����_��:��Om���:���4��`0������ʇ���p��;���3���I���H�#W��3�Pmje�Z!��B���-\���*�g7��yJ����oK�\:m�u=��)�E��s��]�v{�T��h�����Oޮ�B߈��VO��m����>wfc���8j�5Fw��g�mf�}J�gT~N�&#l�?h�qbkc�868��9���{�9�R����t9���,��$�ҶbVw�8so2���i�x{srm���JN5ҋ��xw�ʵϤ ��K-u�6nBq�[����U#��m9)���ϸ��4a��P��hCubF3�5iޝ���s�yR�?j���s����%�|���:x�ӱR�~�P�AK�JK}����+���=?���y�kU�U�o��W�Cj���ŧ{<����g�x�N���=�G�k��7�������LI.�zwl��B�e�}�_P��Ýh�U�����o�k���جW�'�]�=�2w;�,�%�����ey���\����g��������(�_N�p^)�����U��=�|M����d���/�u����ȩ�w�Sޏ<�r8�����M�M��������9�ݏ�չ�x\��}��O��E�/4h�=�MLy�f�W}���gd`�˞�7t{i�?z�Z1x�[�t���&!�7��y�۟8�*P�*7���k�ӹzP̓�ٲ"4�������9|c���y��g~9�I�a~�5��)x��*���_^u)V�PЎGv�V0L�CD�<�^�3z||$���oc��e�7����W3��j#F�e=��c\���՛H��{��u���F�
��-���b�cTv^0M��r���Ԗ����X!�g��w<�.��9����A�o�<�����D?��}���Ot{�;�,ԋ�t�f_X����P:K�w~w��{���N��H\�.��囗�W��ε�J��8�����bM;(p���&�_��UmU��A�����ʖxx������ǝ�2���r���;�ނ��zk9�0o�W��=�d��7JM�j�jyGW97;�:��Hץ��Ϲ٧��Cs|"��4G�M��};XY���G)i֧���z��}�~sݫ��@�n�ozm鯶[��9�D��jϚ�<ݕ/�� �o���7|Gad���p��o��L��
x�x	����A^��3R7���Nϧ���>��4<�L�E��!�s���i��^e�mjO�����f8(/�~�����'P���擠��H��y%�;?O����~����Y?_f���FI�=�q����;z��o]���\�zK	�k%L�L�@q-���[7iɝs�(pmh#���"*��c�隆e��A�)M��rY�d�B,��+��V�DƇP��ݕt������ԇ[��Hg*�޼��L���V�BC���ۗyYjj�Gu2 ��Ɇ�nP��{=Ⱦ�{�S��-��O{��V[(؉\Ue�^'Ť�9GeB�������}&'���Ou�ܐv�gݬ�oIn��5���Awj�G��l�3ٰG��_���y��܇��~]^Μ7E[Sk���/�����)5��`@�{z7��&E� 	�y����1xgieq*]�W�3�U�Se�����9�NY�ס�}q�|7rzk�u:��~]FmA���8{=�γU�wơ.���
B�2��r���xN���a�n �7�Nv���������hx�^PWz�¸}~��j4y��fr��o_�X6P���7{�'x�s�E�G�y���Zoф��X��z�]�F������њ���)l�,����"���0�3�䌓8ӧ��,K���zo�&�x
��Vv�}�FY{����xg�I�g(��*��TW��d)��X�75K�+��U�SL'�;�ۥ�e>���7Z&�o������:SU1,5�M�d�`�y労�Փ�G���2ɶĨ`�z1fn��@��z�8K������0�ۅ�s�4^��_ZӲ��1������.^����~�$7�hE�o���}1��a�^/���Jii��,�����i���yTw�vڪu�ʩ��w�[�L��m{gxC��d����rl���q̉�j|�t�4o3��Pq�y����jY��C_A�����9�/j;�F���#�Y�75����#A��Xs�4U���;ųr��8@�f�n�t7��ZNf����1����^{��t{�PW)�������좝�$���������|�\�S��w=ޖטzz-��N���\p[`y�
�o����R�^X��T��:�2�;����۬͑�:�z����:��*b�^��{=7I���0y>�Pt�;�7�kV/��3��v�y~�R�ww��!b�W���>�/#=9yA��;��{;�PX8[3�ey������}�D0u��Bwo[�Vкޚ-v����58����ގ$�-���k/4�����c�J�#x��sa+ql���II�ژ�Q���C��})��ѕ�;�f�jFe+y5�*թ�KR�.u��q�˼7M��O�Y<���F���{�~��#^��y���ܜ�x.�=��},Й��4]�M�y�ݷ����=B���ß
�˫�sX�Jj�e��}J�A��"U�Q/{�狔#q�8�#bo��z ����NDUL޿T�:�X)wW�^��v�����h��^�~��]Q��p�?j����[�vG���Uq��v!�=^�K����8����o��� ���8�n����و�-5[-����MQz����9}�����1��7����X�~�ys7|Ԋ��L^{��ㆼ���ۉ�$����yU�8�W8y�88���z�����V�f�Y�Q�����x'/�ޠr����Yl�D�v͹�d�ݞ�Vk�C��%y�R�V�Ok9'P���rI�i뮞��{9ZV9킏s��;!����!�{ګ�պ��:�$J�sZ��[q��M�������՛[#��g��y��3xV򶒣qIm�F�8It�p{y�����x;>����,���*��iW�pO��s�WbP\��v�6�Y�����c����r�6�5�!v�����b����x�����]�9� �������}�kg�ӏ�'����3��y��{S��LWn�9-�F���]�h�����o�`�4`�a~>�S���ge�ӯ{}�T��DDV��[�lo�G5�}Gv�q��y�۟9&\ |�Cj�)�o+�yB��C��D��)�����K�^%�uY�,۱���0�#�S���8���zZΟCX���&��N۶��~&��Μ�L�E+�c<~�K�)
�A����r�mV��[z���p�`�}Sgsz͝����{�ӗ�
@5��U��;OY�zG^h���yֳ�{��� �P&Ei�#���>x�s/�+�Q+Aw��C�)�K�Wv����I�*N�;��vW��>|/���['NΩ8X�I#q��k��L�\��q���A���Ʀ�����4�"�K��[ԡ1a}� �xD{�sҮ)w����;��깷]{���WT��%���xh]Z�;��d�otJ�[�w��β�d[����*r�D{NEwcޒa<4�aVi�<w�u|����͉�r=�O��]�R��V��V42OY�/�r�l5yM���D7���zfSo|����=�l�Z��G|3�����k�����n�1޶��U�|�7�Xw-g��;=����Q�էĚ$�7k�����Rِ�Ms��5]+kӳ��ζ���yy+� �ގ��k$���q��Q��٥��*�P�.��O����R�|��������y��P��øI��Y�=zՍT\P�9.Hu��������G�ڪ/}x_I�~�~>��1����dtv��4�����/9���3�Q:��V��m�uK�7���y_�y.�0I�g��1Ov�P����~R�ؾ��N�䬿���c�x��)�Aq;�L�匏j��t�N�D��𜡥��{����ᷚa�7��>E�Ϯ�z�E�L� ���z�>�W�>��~��'������A����?�8`, �������=����ޔ/q�ǫ�WP4p�X6��wDQ��ds_0�\�9�]J5r�:v���8��f¦���V�]�{ut��N��w3gM�oo.��ioKR{V��;���ٶ��sn�͡Wݯ����rg7��o[�U�d��C&V�ٺ���{�R�zu3_'O��OI�p[�W]}���oze�آ{Q=J��
Lλ�I�k�xb'#SM����T����Wɑ�(���}̉�۶�����4
�7de�R�v\��w6����=�]��x��d���Lj���ݮ�+:�2'`h�q�l�R$TD ��zŲ�^�C�|a1=���3���I|W7*:���.�+�bl����k��Yxo�4������Y�1q&���FEK`�V}�q������gV�m.S S�XD�5?Q�I��sݽ	#t4�q�]���U��]e��|F#�na.Ӹr�mt�[�92��_l� ȶoT�V��M:�48oV��n��R�4,��c���F���d�Dw���\�ʅ��L�<n�d�R4��T��ծ'�
���n���ݬ����PXU����l�e��3;"ɚ ����<^�P�vk�E+q�]�_i
v���;z�ǡTыc|h��8���n� �`���Y�!È��W��w�2u��GA��eJG2���Nuu�1M{�1�U���t73`��]o-h�)K7�3w|B�(��i���O�vU�0�/�oucH+�Aaϕ����2^�;�(���Uo\6���Dt������A~�SF�����v�g\e�^��S��-��������M8�*uF�9�u.�gJ8&�#f�ǞEb�2e2s���CjY��Prl���	����|®���5o�PO��"e��19��)��ʜ.miő,SK�.�n�Cu>r\Gv�%Ǐo^�mI&ɲ�Be%^i���͘75A0\{5Һ$��>���-ve��:�}l�����΂;�T-;�X�ct�^�{.������j��	{tm71�B��F�!�Ȏ��X8Hl=�tk�Rft�kKWv@HZ�Q��U�·�Xq,�@	���˩.�E��r��|�펎a��%
eJ
��V�zt9���ޗ�n��Ѧz�D����nM/����W6�\�Fv�U�*B�99q�f�����v�;x-�IL��L<��.�ϖ��_Ry#'�:]�N�����ű�)z��-C:�k������z��e�0/_>�+R��=��iN�+�2t�<����WV�^J��v���A���3Q%���ɦ�M�V�@��6�d�PκDظ;�8[O9��Y0�b�s�ْ�ic�%��9���ܱ͈�rĚ�jW�{^Lܘ�θ���N�k����f�Y�7��U:x�ݹ�ML�N5J�3xY=)ا.pr�+���]˦���:7-�4�jt������t_]��x�>s����έ�u��z��u$}�� ?~$�UU�%�$�)Z���r�U-T�y��U$U��s��-y�Բ��N�*�N�KEI*��jҒ��%*+�rT�*�#�%-JT�U*Ԫ���I�9R�&䪪�s��r���8⵫�qYJ�*ܷ5���奪�*�JZ(�%e%T�o|9J�$�VU��j�Z-*�V���T����7�j��Vw�d�dW#��R��Jʕ��5MRJ��8�*Z���j�V��UiG\�Ww)N��SV�%Uj�Ej�J����[U$��T�D������ZU$RYEk�qV��+UeT���j�#�y� P��`ýM�,��;A�o�f�ȷ�hk:�f����<�J0ۍ�	O���3��d�X2�V1bg\��͊�|Ɖȗ�'b��#���L�d_���E(UI��Pha>؇l�vl���3$*����;s������&KC�F;6,�[x��ca<{ɲ�-#��Ӈ�f����La3�b+NgT="M��\l5�6\CqH�i�����>��i';T��0��CPoU5�|�>+�7w��1Y�/f[L��>6�"�����{n��m�X�}��#�k�1<#x�[�Em�GLsI��I^�V�v#t��Ux0'����=�Tg`��R
yu>��V�w=؍}PÓn�G]�b�t�&�f[k������3-�8Vn }s��#�w�^J�Y���_t��)������ܓ�Z�,v�Y�d���'�67׎B��ϋ�r����3x "���'���v�ײk�����)8�����j�{B�cjrr�R�}���[�هש�|��:p�KUƁ� ���%P��TR����
�yꩺ@ٔ!�w7^�_!~8��{P3�~>b��x�̥��0ѭE����Q�]i��x�TvW�ϳi�P]^+4�4n��i��tD)�F��d*:[�V�R���G�ضI��y�;��?p��%�4ib1�*<�nc�nQ��it��(d�)���b�8�C���ד{Vf^@�H�Yq��f�Bo��O�t1k�gd:��E�E���:��MO���{�\}U0��M�
��5P9��3�i�A�/�\:;��b�T��zis��&]M2r&k����8i�Ŏ=<�p<yͳ�]�����H^[ɗ���y�h�[e�0�~��)U&kg�е��y\�}����k�a��v�L�i�4��xqʉWOL�./�P͋.=B8��m&�qڌ�m�,�hJ��TX�B[�a�M%�g�xuՏ]A[�VKH{�-BC�sC#ؖ����X��x�w��]'^'|+�@�%Oo�񦇓�#-9tj\CsѰ�ݯa�qb�5�P�-p�����s�9-��I�=�� k�$*�L͓Ȱ~̹���/�r�o���z���#��|�L�A��3� �A�@��Pz�MY��TY��g�����ܪI���Kk�bxs`�CT�d�ə�Q�D�P}>��W]�/��w<ؒ��>Ր�((&�ˏ���.M򛇆���k��T	�*�\Ib*żի�U�7�@�Q����0��ҵ�c�m�m
��5�)�5L;��\:`F�smt~e��|�eB�e�/�Jsz㓭���5�C�vy��{.��Q���PP��\L���d٠V}�;�>v#�[eIXx�_eiӃcvW����2�;I�]��J�Š�Gb�YE�� �E3
9�e��r��xUw&�羙��F/���3�����w8X�(.zY�l�B��U���Ev:ny�J��j��v�I�&�r�zv�B,KAH�Q�6���;=\/��q�d��V�`��K^^��w=��-Z3:�4�U�a��oU�Kq`ѣ`��jȰ��œ!�{��ꆝ�"S;�b�D�ݼ��3kt�"�7�Q���Ɏ�m��EI�.�!����A��ã6*�)��B��}�p�L���RaET�)�EJds��h{�� �\ZX��`!|xk�y�f�Et:�A���O)�_sH��h�i��:.~W��CG�9�pN� ��Fȭ�;�����m��R�;������G�=B���eJjޘ.VGs�)�o����o��*�5����0���wlga��;I�l�������%u�¤��Z�k���BW�o=bz�;V6�vϨ[ ����4,��m�����酈�}B�1�S͡ɛ�	.�=tF]�z�"2y4ĨStp8`�SƹЌ�0N�"uR��8&��GC51���m��iM�b�d
����w��Kͧ�
���5�'��|�d�驳E�ˆ�yԼ��7�D�%�,�o3�[W,'�Ԣڤv�>6���͔^'����C��^\�ۛ��+U����z��Gv��/�;�\��ެ+�#�r��������y]3������������3���Z�vJe0�ʿ'�p�>ƾv|�Űټwh�<�nU=���ٻSa��M��9����;�وA��i$%6����*�֯��wt_w�E_\V��o'�ݴ�s�݃h�������O~�|
svdKP��.��پE�M��
�p��S��>�[/5:س2�o4�Fh.9�i���Q���fDSRj���&��ɍx��� �GJxg��v���W�4�����z���&�(Q�m�e�7�����q�!��'���C'!f��1Kp?��{t��M������7�uDf@;Ve��E۷0��B[��N❈1�i8����m�xΛ�%��2��TĹ��m��(5�{�v�%K牰��\�; ����Nu�Ѫ{j+w^tv.�<���J�^�b%9a`����M6pY'_�I��Ƣ��G��ѧ%���5sj^�֍�ׇ�Ae6!6�ݐ[@}�4��J�.]�Y��3�+<:-ۜw@h~�E�qH�+�����t�Ɂa'�
�q�e��)�T���bDk`Ur|
 �G<�Gk�ym��Ǜ��b��z�w����Y����Ի���N�XlM��"�kV����:�h�6�c  ����n-̺���f���Fe���ʈ��i�i�N��t�.Q��n͋e�IdV�Aב^jn�:$�ffF����}�k��`U��`�M)�v��ֱ$Ϙ�]�|��,6�;���9���X�bQ�Ylt�r���s\���T��;���?�5���DƂ����O�e�Ɣ8�M��44�begBaR�L�A�lzQ��#���(��&���y�x�Ɠ�a_ylG�yQ���:]�ȷʒ��l�oSR�uHM@>q���c�L�(쎊��<nZ�pv�3Ͱ(,7y�ǉ�n�kle��[�F:}.�T>:��^�H&F2��0��(��P�[���F���4t���Ej�<�9��gR!{��8jI���s�W��o[������jkfJ)5[ėq��6��W�o�[8C��a���p�QΑ����W������M��FIR�hʥr3��O5���i�{N��-P_Vlg����S �f�=�:R�ږjț��D�^���ܢL����ш�隴4�s�R�sC6^�e��w�i�{/P��.T��C�L�l�S�	��Š�ʝ���
���:���,�J�{�k߷�3?n0~nR���:N�&��\F�؋���P	q�E+��x<�:���>=��©LC���ՠ�* �{�玕8� ���Jo��#��
�{��IQ�ol�n���5ZI�]�O;�.ê�yG����L(]�+)M9�/n�O��c�6�K�d��k�ٴ�� u���U�ûO��	���v�D�{&+�\�S��ւSx���\k�2Q���CDl���j��������d/z5AgX]j�>:�qn.���'�w��d�)���$���ާqNƾ	���_��H�"��1�~[)�,^�F�Q�X���F�,�SmL�0%�5|�4��S�ݔɺ�����-�e}�^�����h���B���&"��9��x��i�3�:�YCع��t�^�m$�8�X����`��C�髉n5�ƃ�T(T��X�M���\�U?���e�ǟ���7-�d�و�̟�P����.��	CmT>��3��;B�R�evF�F�?��D��6���ä�����d�S����Pw�������Y�c���L;���kM�����n,�ܜ�i=3w�/���ā�1O�=U����9ܬ�P�C�=˿,0��r {O9&^'/q� �j.-O8@�	�~--��LL/0�]����d���O�7�5. �Dv^�/�J|U>*�J:�{i�o0�H��U6pvI�;�|2]�|�%ڑ�e��}�tܮ����5yk3��y3��1��)S��:e�%��[�oUO�MӠ�9�,���Gw=
�{�׷oX�L���c�(<�����-tb����W�V�V�׷Ơ�q�g�^����큉�-�"����jbj9���M"~q������n��	 +�0˕c��:�ʧ��i@Y�e���RA�j�r�_��9�0k�C�߁��uM���H[�&���+,�gm��U.q�n��T ڌk��nƨ�.#e͞'ԯ��(u����QS{��6�b��p2�Tm�z�)����k� ���.l�+o��qM�b���|�����;�X��*�E����M��?D��()�
ʝn�#�ScX&.zX�լ��Րp@yҲ����N�����o��v�"^4}�Y��������r�����-NeRm~��" ��{Ǔ�ɘ^ɮ�n��������QfA}&|ݹ��K�2����C�FY.�;��a=:0�ݣn�����x�Z�����#v6��d��&˽�r��,�y�鶾ͨ�y���+eMsl)�����Ά�<7��y���i}<�[x���9�y�%���s�D�s���W����#��Ҭ�1Q�K_0�ڭar����x�C�>6�g+��%�a�n#��F�/#s74LR�gM{W��	[(��;�,�����K�����[*nVV��1{f�c�I�7�Ygu��|
��i�s��8f3wQ@�1%V��������1��8֘B|������b�nS,9՜��T��$S���rUm�`͎���? �$ ' ml!��4�m�t��1�Պ�tz���6aR���Ψ/Adw8�N�n���F��� 9�+�LGS���A�@���+�%�缪G�/]:?K��-�mH�*y�6څ����긇APZ�rC�>�I�e�}�d�6��l&���%�ʹ�v(�l���c��Y�{چ;sJt���(���8e��<hyЕ�E����P4y��SfyT!�։�w�e4�f�^��o���:l�(I�kLv��V�>�v�#�L�<�ʖ܉����CD�B�O }�f�dl��v��aYڮ��D���\��m	EڢC�;p������6������癯��"~gs$ǚ);��୦͘!�n8lI��O��R�m��؀Q�\ʜ�E�׭itC*�#zX�H#̆�"����)�46��L���KBI������!��ֿ����lI��~
��ǑU�쨇�zw�f�6-�DP�r� ��nQO᭻
ll��&�-�|wS����$����K&ǳ�Դݬ�sl��I�1.�+2Ð7��<ҟ��I�ۯ}�Pu����B�5�||_+�]��**ƅմU?�V��H���}�=CO2��9	������?��M�S�[��U����^0 ��4����}�F��j���m^�a��v�fC}le镽K�C��=>��< '�9�<T�5U��dJaIL�;�U2.s���ʜa>*,����*������C�&��Vm�r���"9��}��<��E�%:aet~�����W轃gԹK��('��ҳ�/A��B�f�N�c8��<��c����@M��<�Eŀb����/��?6H*V>�;�U�f�7Ð�gN�WP��(�N0쵼��ǧ��r�=�y=�K���q;�"�P�wJ�z2�P؜�k`�k��S�}3�i1�<;Ks�����ͩ����
��R�q�Ec<(x�����Q��C��xq��v0)�����0N�Lh,`g�u_�_OE@E4�-r�0V"Q��d�LT�����y�T2�RNtt�U�j�UZ��v5�>��,.�j����\3�q9��f�vQ�BK��S��`���W�U���=�c�p~-x����F��s�>����{�ĸ�el��}݁Ra|f�:;yX6��/a�rw�Q���M'����
f/(�k�Cg���3��>����Z�=�/��)�Fm��x��-#C�^!F�+i�q;4��'F�F��*���#�=��=G�#��2� ��N�Ȯ�X߹���q�B���yg��S��{��������*罔lBdy�����M�Ul�Ɋ+�L�]6����.[e�v�X�s��y��b�"jhv�� ������U=�,����Tic�����i3���2����)��]e~�3$fVozЊ�3}��c'��C� *X:�6��,+ﮟʀ�Io��15@��1��ʄ��U^�cFK_tH�y��۩ZS����=���^^��bw�@�)TH�f[r��ϝ��*J���^�X�?_�+<(KK�/Pc"�`�[ku��7#�OY�)�T�U�Y22�\�On\cQ`��y��xҪ��X�5{7�o%�a;ږ�-w�ad<z�'I�N��$��<�}*�d�/�XG��PuI�5QF��7H�X'jO$�}NFe��z�U���!B�J�_
�O��������)E*U�[T�p��h[��s�R�c�?���>��U�D-m��H�%�(�ZWy��*[�d���OV��S֠M�KP�YbZk��^B���M�h�.�Nh�9�<]x��ms�z�Z͎:r�5@Y.����y�{ܪ[��tb<VCs��[��a�Ag>��Cr��0��C�H���Q��P�Ϲlm����V�u[�3a)�����4����Ǔ��V�R3�������S�f�4լ�(�;��*oU��� �k�9��]5�;��ɬ
ر\ѳQ��֖m��[��Q�̢+;��V��7���6�15i��/�ޘ�Y������g.���F��h��]:s���	3��O��TrJŴ/�q;�ގG��e��ps�dZ�7��G����M�����_��r��mb��n1sm<�έe�u�:<���B� ~u��|�kꜶ˴32�7u�6����X��b=\�� 6�2/[;RkQ��j�hVo1b�/���a�h�v��O��si7yNd��P�vL���ˉ)RĤ��qfc�IWw�n�s]��Ř�m���ٸ��wC2D�oׄ�+��S���H�u�J����-ت(���ԯ�qB�F��a��u̥(�m��n�oF��m�>�1]���J��S�2WwV;/0�tr���]��
՜F�J����A��m2���gM�֤���Q�{E�չ���T��-s]���E��y��2Q�m�w{ȠUK��wq�p}��x[�f�f]�Vp��b���g�n)��'�[szu5K7��-�P��e�ԏ���ί��չK=��Ko�{\�IR��Ɋ�5y{y*Ŗ,]�r:b�X�;a�n��o)�����s{Q��w1�c���$�`�����PӮ΁*B��{��u��kUʹ��jq�:{V+���w��`��f:�ۨ|�d�n��]]Ԡ�]������w�]�k�|�r{�Ѐ��ە+3a��;�nMcv��u6�JY�C-%�Y������KY�+�i�CC0�����k�p���O��*���V�FWm ��[k;nBi�u���r�t�=|�R�*���gV
m�8�M]��� k|���g@�{-d����-S)�N�km�s2^n#P�W�gk+>0�Hj�[�wLW/�Z�0�yj����ǐ9�n;��,{������<���	��v�oV6f�]%EX�[���f#��ߣuɹ�WoVIwQ�릷U�rZӸ6��S���E�bv��Q�E����R�]chw3s:��`Kz�ݲ��[3xT�D���2ˣ��с�'0N��9.l�2�8Mi�.:�F����&a�v�];Z��e�0�B�\�=a@�5��;shY�J����&#Ӝa;�riӒj�T���i,Nwp���r�o�؂!]������ͱ�k]^gJWCU���N��7��'e��ux�e-�ZB�g�b[ʹ�z�����
u�Ӻ������٭�H��폛S*-�b8�sj,�7#�z���hb\��[z��C8Aҡ�t�#M맗�y}���ɄC�� T�b�J��\�F�y\��Υ��yDU3�j$A(��M�bB	tb�O
��g-�i��/5V��:o�8�u8E�6�}nn�n;�f��F&��"��U��/�
��	Ř�qq�1��bs�gG�;��WJ�v��{�J*Z*j��Y�9�q�8UT�N�p��Y%�Ԛ�*J���e2�J�U8��T��r*Y-�[]�N��K��p�,�*��k�7:sr�(�K�ӧ.��NN.E�:VS�q�p��8�}����rڎ"[qq�̫�$uËK�z�:M.J\9����ss��뤓��r�D\U�+��n"[�E8O���:[�EÓ��+��q'75S���J�[rqsY\Lz�sV��9�9���L��r�U4�[��ճ��M�9+w�-VR�n�:����.��[��X�k��#�R�&ܲ��q�jeK:��U+t�WV�T�jI�W'%59�mE+"�;��ҥj�j�:O�YZ�_3��T��N#�9�ښ���9m�r�Jr���m�nG-ɭd����]� �Ac9�S���a���uAG�lG��Y����.�tެr&F<���oj�δ�^P؝�7�����	h9F��e6�,	�����C��3x0�7H�2˦_�	y�_<���<h_(5�,��,�]�&�W���}��8����c�t�V����[�D����|����iO��F�8z�8�(���DgzUW;�Xť:���W-��K�`�_b �acE09���L~0E������5&��g��[�jl����f�z?Y��W!Z�G�Q-��a��v!���1C��c��'��'�w=�%?JՉ�x�,�����"�\}sƼ�����hLMPg�8>zCzz���������5nV��<�k�%���O'@Y����*�6��*u�;�MP~��z{b�ꛚ���ﳫ�D��[�����ׇd*�jZ�ؼ%�Pe��L6��ŭyru<�q�.l�6B�[)M�
���[w���["�#+�e�*y���uJ׳��)z:l�,��F�4�2s��ӐG_4\^V5�>>��Eʩr1�l�a�fS�&s$��.�	�s��VG-K�P5��Saǻ~��Z��t�B��L�x��P.��7�fo�Ԟ@�Y@md`op͈�7W5V�Q����q���[o>��x�+�ت1������Bv��n�lv�>�9wWm(��g;'R*�)�[ ���_\��r�c1�kD��,o��|��8x!o@,-b+v,YU�e,�꼒�T{�®��5�������=�;y� &���0�������Hu�6����l-�x�j�߹ml�bԅd?}*����4i���4w��dQ��М6�v��E�͕fL:3:L`-9��jWU6SGE�<�N��>.�As��0�x]9�P���y/|Z�a�����9QR��)��j��Q�E��Hd�u�C[��4�;j�I��r"�1�o�=��N��6��_�2Y'�C0a�Z���DF�>��uk���A^%�aoCg���C�:�����c��6����~�&��Dޚ���s-d�=}�<��je��~t]�r�����ا�3��d������[��YQIRF��]d��&�eV��G���]�{�[�a�2w��xc����l�HH�����5R���	��[���y��h��1�oH�3�ׄ���b���Kϡ�^�"#c���(�ztM�&�C��BK�M�P�k���D��v[��p3��`BS(q�U�������|kf"y�U{b�j�u�7S:����鬔������Bǭ�)ܽ�B���+�)�<����`�Lb��˜�9¢=79i��y|zS����-��&R�V��Ьl++NE�Jn��DBĒ\�����AXYXź5	�-F�'�l� ����o����n�^sJ�p��.���5�e���5+&��R}ݚ��ȝ��b[��1��F-�6˹�>:��w����O_P}&�K3+0���������f�\%��F�ƶO��C�a������}�)~��^���!�]�%�=�A�Qi]�d�[ ��\󵽛��p����D����S9���� �ץ�5H�WxǹL�5�����tGs�7��i�C>ܺ��Ѓ�y���
4,-��_����`K���]��y�{��4��.˵v��e���Z�����׷zҚ��W�z����7f�����5�$27��^��ԅ�!>L4�&박Ss�t�mZ��+�ǌ_�����3�~�x;�V��ܺ.ܦ2Ǡ1�hOPz�J�^����S�yx�y_�I�c/��*Q��S�Ԯ�!��b�����BH��Y4z�����i�TS�E֦lO�3(_T���N�Zlbk�w郁NcYS�?Ap���(��������>���v���1B(�\�L>�j�LvO��W�cћ�?6A��#x�� �yN���x@��Q	��¦[gۊ�[3ɭ�>װ�V达��|q��tl �sr����MDv�y�w�	��,�P�_��-��+o��K�cn��ڻUi��oi�!.�����Dw-�����n�a^[���a�غ�����ۆ�Ҝ��v⒋��׾�N� �z-�����-žwB�����jʲ�ۓl@�g����l��/�|�@ʑ��}�w���m�8Wm��?�U��&fVl(��
͵�f��[`�����=^=�<{}�K[t�o�J�vRY�;ϹL�W���:y�����bx�%M����mZ���{�O%4gQ�3�v���R7��O������ q�h~j����lvKnMD�X2^�3)7f8���-�4y�a�@�&0�{�ҠP��#�:S��4SI�{!L��[j�+[�{.S�p�I`�Hs��=q�Z_'���>�ջ,C��ܑ��ۅ�8xZܶ_���fX]�R�vK�����iX ��kK�h��^����������·ʓ�y���g����t6�˰ƝV�.���`�Io���1Fo�O)����YeT��oF8uK���"��Z�*k�������>�Q"�mˆ�e���d����0��yӊ��\dī����օ�Z�_.jGgt*汆d��,�i����Q�f�[�jwy�8��#�@2V��eX�z�����~�2�s�7�x�����	�N��tRr���Sx�j����XR��{1��u
��v�*c����	J]��GRvy����"�A�Tu�%����G7�Ӭ�N�TJ)�R9�m�!8ٜ�m�Y�
�6v��9�􌥑o4܂���zY��vY6+m2�ކ�7�!��B�g�xr�Ӟ��IVcn������]z\�.l�j�5Jpӥ�;kM��2�>/3T���\�ƬR�ܓ��|.\��}fea��Y�Y�V0�͵m�P�l2�Xj2�
4�mFj��o7
�ul�ōT�rA��&�����}��`^�G���C�rj�@�^Ă!�q*p��>i�X&�&b���8Y��X�p���,�{�Ү�1��/�X��D��Qx2�?2�t�˪}��H�{���ѩjF�A?�ll>6�X7�����C��a���o8�8�a���т�ֱ~�p�fY�ж���Z���^���g�+ܶ��FC�0�x �������S���2����W�:a�7������^YX�3��tv@���m�wS���&�_vɇ��d �g{�::8m�|�(������E�o��M�u!j1��j��颲_�_~���z��x�D�;�=<Xe�m�g��,�����,��N暥�K_e�ъw^Ξa�q�wr���M?SS|�+U���c'"��a~|ƺNv�q�k��O���z�g�#��>��Ƽ���%����s�7��ˢ5�o^�ì	Ȫ��~��y
Q���wsN+�-��3���%RA�QNU����I�k5�E��u^2�TDda�{W�m^q�����֯�+-D{�!0i��lf�]gQ�5f��f����UBEFv�_m�Z���i�	Q��U]�w��'t��n�����ؓIYR����[��������B�U�']��k�ϯ����f�ͱ,�++1�)���3Sf)�ڳjͶ+l�0�%�o<�]J$Lln?�K�8��{�C��UR�2u�'L2WC@��ا'S˗F���@�nbm��ij����txPv��`Db�b����)�����&𖥑E��Y>���e�7����|�Wa���q��7�P�cוtME����hrfS�19S��#�ScY0�s�p'��GR��c��zY��R<��m�&�\]�[P�o!�U��Ρ$Ů� 픧e�������Qט�a��_*d�e'��S�M��x�����}��Pũ
3�3�O�-b�s��U+o6����04i�ͺrAg����{>G�v�L�������EɁ�
g#z�Z���%��k�ǒ��^C��4�W��LS�
*S#��y�����gO��:���ۮ#��;��8��lNA�A6-��p�4L�ѕ�=,Ҟa�#%���&svoד�W?x��g�X�`$0�u����ޮ-�'3��2$���6����ԋ��ݸ��MG��oI癈r�OkޖLݢ������Oɍ�\A-|��H�����Oz50`yk[*��!�ZJ�CgɐK�粐����	�tSսǙ��=�Ɨbݓ�+���}j�J�o{}"���H�͘�'�7M9'�Y�x����f�6��7*���ͩ�`u�&�|.5�ZJv��������yqЛ�����N��N3	f����3���y�x{��y����6�+�ORc̒[���]%�-?3֪�mn�A��3��.w��xc�ņ
�]��e�H�u����4�dĨki@I�i�������J����[
��5�B3�@��@��t3�i���A�A�L�Ȕ�;uF�Y��etX�����A��.ց�N�r�By� �8S� ��؞��m[�Ã���i����^��DH��.*&�#�N;��Ȟ7�S
��Z��<�9�ֆ��4��C!y*�>v���������L탏����������ꦖ�vAn��� ۢ�.d��h��sUp��@��p���a?�4s�N��^�Y�����8���W�T��[Ct1ح<��Ll�A�ॡ�k
w�Zl�-�3j��Ǵ�6 �B��j�L�JV�b!�Rd���%�h؊�pJ�M��2G�B;m�$.�nM�g)�i����hY+Nva���������^%�;P�].��HA�����s�a 2����8�m��j�RQ�/�<z��NɯV�=}�#c�&m��-�&\�1�h�=A��*�{"S�L��%V�K$��[[�:&MDR���M�2h86���+�bһ�"gb�6>0q���u0DgG%R�s9D�N����ܓsiN^�]y�g��X��*�I�ƴ!�K��l\�&�$t�u&.�S�,�"YZ���(����G	Qug���ŧ�J�9���������CmLl�m�Y��ot�+��9�'�P�&����D�	��@MŤ>�R�ʎ.�E�g�7��(F^��Z˵���+m�)���1��Ӓ��(�}#���.={�a�8�"L�������^�vF����!qH�:��>m���lgin�O�����l�^N/J]EV�]�/��T�md4����B�`{���0Yi����9ܘ�Z�@~}埄�Ͼqd�ʑ|�\�A���	��UX���['�jz|�)�� ����lv�=�ǍI?G���K�	�˃����o�k$4�D���<~j��et|k���-�{��6�\�6.�C��PMg;�.u�b��=�"�Cn)m�с��Oh�����8�P����Ʌ{��I[�N_st"d��VHW�f��->�TP�f�8v�4��v����}�!���A�v�]�m+SH�#�m8z���%� �9Wə�}��Д���'�λ��;�w{L�f����;�N#y���Ab��Lk�
< ��c�Z�B������Jd�jm5�V��xSL��XGo8mM�f�k۹��������t
�{*~"��
�.,���:�:ܗ�y/w��m�#4)Nj1�G�[�Ky���x�4jv�^u��a�ѝ��,��3V^J}RĹ,�4���[`��Y%qP�\m %.��x3/x{��\���U�������kmx���7�7<qRY�諚l��*H�a%}��<�$��~���K�NO�����B��)�]H�y�]]c�%i�)��o�Y22���
���ũ�1��.���wS �����H��k�(pŦ�H9q오�������c��X��K�zx��hs�ۢ�s��̞�5#��_�7Β�B{��ݜ��H~R��<)X�e�5�jm[���"���W�x�H��/�֯79=���/a����x����՛$
[�����)f���9��<컝k����R��k(l����48��dK�疃�4tyf_-b��u�a�5�����S˴�3�Cz�X<�=ڢ�#u裔8nv���i�A�7�5D�\�Fuj��^m�_�D��|�SW��{4�?�.�8�����n}�d��xC�P*�nMc\;���20�>�/��]�m��Ў2*��L4��nOV�|�AtN�o5Gr�79�ۚv��mM�B4�KG���v�`R<'�[o�}fQ��2(p&58�(���-,����Oc���;�o��!��i�G��G%u��C��	z��ӗ�B�j����KoE����z,�oy*.�W�~f��>K�<���8��fvBf�V�����B�$L�7�i�M*7۪ʭ���G������o����1�t�{j�5�٪j�����x{�ox <��Ĝ'�A��ى��{�x�0� i"��0�Y���5�n3�s�����J�Goe� Pׅn�
�F�~��+΄~U�%���:���V��P�X'�!xǨۅ��0��(
�:���֤�gI�ނ-�y���B��ޚ�<���'^_�tlL����J588�g��!_��K~Z�>e,9o�ߘGx�Pa��9LkTS�-����#�Ş������:F��v�W�V!F���	q��6�7K���Aغ*�v�y�9�8�%������\&�sd���7)Qn]G[�����U,|�c4�z��A�p\c��M�6��C��xQ&��5{6�!��SF6O�͟AׂeGn�pi
Q7�7b��t���Ҧ��Zˠ�͗9�"��U�����p�$-�CϝB,O�����7؂�1�4m�V~U��i�&���|">�����]�-�x�j��-���}w������W+4L���]�@�ea�H�@t� ��A���]��9�^)�\�S�j��ջQb���� � @�,.(��17=澞~���8�F���Ǔ8*[�VQ��n���
vRT3b��5�jVa�B�7`Z����Wv�����f\��=yϥ�<���9�fi��>�dD�n�c<8��T�`(_C��Sb�lA��a�m֋�b�_
8�!'ҁ��5�B��$*܈�YvE�{6��(5q1b��6r���7�1׫�&>�Z�E�H���T��"�]��dWAJ�Nv���j��+��1�Ҿ�t�s�r�{��ƶ���Ce�'�3Ck;�ŗlPy�{�$' ��C�9,���5��k@�&���Z�w@w� �X6��*����^eWX�1>$��=L�j(�i/�k,��\�p��h%c�t3�]3�sn�T�k:��\wV7��5�lSu6unhɮ�Q{�*�H�i�|~k^S��5֨��U�޲Р�)>�3��F%!ZJ�타Ⱦ�n��Pݎ��<=����Z��Յ[�g�,���3�?66 �G��
�lՠ:��S�+h��u�:S���G,�Y��(�L���[�<&��r��".Y�VL���;�c*�Ϧh;)
�2G��T�r�9�ł]M�T�i:�݇�<� Β�^Ɲ�Ϋ�ʼ5���u��:ce�1��dNt����12 ݩk��z]�|��ؼkh�!�*�؛1�!t�Y�`kk^�`�5��sM�̓y�*��G�Ɲn3o.^���7j>�Cz���ʵ/��ж�o��M���눖�ovک��f�V��3E�&0F�/sz�w[���EU����k��,`�#x6݂zveu��[�T,�����-V.�՜��(Kz�0_p"�U�Pp�,��oh� ��L�"��[K�R��Ll����������\�O2���c�\�ad�eu��m4��� ���|��F�l97-p*)\f�awܹ\����5����*Z|�[����z�%�en�թ�x��b��yC��9]]�WM�2uF2��)�#�����4r��޲�D:-�f���D��9[r�?�h�4��t���g���{���F��D��	�����ޅ��%cMs��:��]-�q�Yڰj�s���|q��c�۽��$�&��v��Z9c�dԣ��ΫQ���ĳη(�ھ5�%�*٤��m|dt�k�	�_wVw7w���b�9��ok��m�C�n�]���wR<����]1�@��k�6�D)7B*�K�&�W�i�r�����	WNN���c:��[�l`�Rò���L�oe��xr����.�n�u��̄���]�Z�R��N��� ��W��^��1��>�wt���cB�di�jpp�n��,�B��ݼрeA���-[!wD2��f�E��+t2�Cb�>��Y�������s^*�)^�'���{�w���yz�Xh�o1�r�;_��F��b��4N�g`U%Nӛ����[9Hz�}�$N+���$��[\32�wʯ껻����\�:\�w�4�7Nq�n[ݜSˌ�ӊՕ�i5Z�\q�sJ�[)MJ��G9�T��QL��:�-��qUkMIT����VܹikMZ�e%�g,��gW)b�NJ(�[5jڶ�LJ������';�wls�6ܶV�"�wc���J������IZ���Q˕TՕ�MYM�m�ܩA*ڊV�ەmZ�Q-����Y�Hԧ'-TU1YMZ�g�qW�6���cͳ���jյf�YB�Tb�9YU�K�9(�U6��������3)$�B�7��X�^�v������-�QϹ୒�v���Hyg�R5qWC$(�/2��h������j3�ڳ�<��vu����7ry�{����  x]�^6��ZW�/�d^��<���z��a`��=��L{�9����pVe�l�,�cA�]x����$q�(��N
nɀ���G=rh�5�,ҞaIt�q=��J�d�u���4�0���Al:	��%8���g�%��?�_X���-6��S�����߳�ȵ$�13�LN�(�Z`󌴧��M�������`�>iw8�A���j�4�fw�e�/;�k��R��8hb(��|{O���d���x_�y{�-�$�0�/������j�0��92w��U4Jɦ,jx�3�4��g����jKP1Ba��ͤ�9r�@������ȜY��FF�g^�7S'�e�g�����'��������`c4���g���huW���E�i��2j��D"�'ҙ���x�{��v��aY��l�H�4���.��I�&�=���� �7ҋ�_����g�� g�b�\�k�Zo��v��Cq��$��^�A��'=���	�V{����@wV4ﮙ�9�	ÐySƄC����ϼ����Ѧ̴Ke:��+��4r�+o���v	���엃T�e���Av��d�z�������R�66�>�f{���]�� �g��l���x�J��(��ﲽz/���[�y-g���o����@�<m�����g���f\�.��h��}U_��xxz�f؞�Z-m�n<�^��&�����}ؠ�ϲ�Sʒ�M�'�tt4:��/z"�WZWW��p1�}���C�܀��s�J���Q,���7����b�w4,��
���T��{��J���:�T�|��CE�mb:$��fSª��e�C'Ԫl4��n��ۤ&��[�%�O[���+�l�	�>��4�=!�U�{�0�R[�Um#f��s尢"�o[6F�uPq��T��KmQ�]��OM�쀚/�H}�(��4���t����ſ	 ^��_���QFB��Ci:��}	�\c��RK��(��vm�t7�qS�lޱ���hr��&�E�����i���K��$v�.�h�:A{Z[��hwt3W=ì�
�G<؍���q�T��
SV@�O>��6Ӣxk2�0FO;�]���ؠ��=	�j��%7�Oҷˎ�$~���ܵ���/�2�G#�_��ҟ0ڦpKo
�:}�h�DU�}��{ȥb�Jb��0x�z�|�2�e�F�`�;�I�=�}��B�H|�3^��"�W4�[��Kx���}�N���I�W�oWJ��nd��˄?�e���9z�u(�ӷ�s���uX�f�r��^+Ӆ���G �?��j߲+�N�?vU�{�"�k���Ұ����;U��X����D�w���u�f}&�e�����{h��7V���f��s2=;&���� ����"�����v,��-���+�C�`&�&��y���� ��~�/N�T�C��.4S�&ջ�	�P�ָ���,쿄U����n�dA����ɓ�1���'|�k�mE�v�]�1����y�I�LO>#�2/��������-��m�R,g�.���' \�Z\@�<K��X��g�f��ȅDp�L}�fڅ��l�aB��`[U4�9\�3�I�%�0�v��"�/n*B�hա0E�#���{����X,���P��H��[�D�[N���;�Q�/��q�}��G4[EF�pRr�d�l�ɀ�˩�n�݉\p&r���׵d��d�pT.����;mf��ˈ;x��N�n�$��N�(��n7�G���V<��'{[^��-���(Lc��tr2Iz�4��^<ѐ��8�=��>,�d����[�����ō,}d9T��7�Q��fH���t1rq�yXοd�inL9���x�4�Dd�B�@ۗ��A�Z��NkB��~w�D^�J�2p�)ޓ�#�՛��һ�,K�26j#l�u�~.�ͧ���D�q9�IS�nx���.�VI��9~�����\�C��襄���f�l���Ep�KouB�B8n���N�Y2��s�(�S��:��2"� ް�g)o$������n�,[�� ���c=�H���S|�&��n�j��u,MB.��G����ҽt<�ԗ�a/r�G���=�W�DZ��axh.���~�R)�~nSA5ˣ���+ɸ��h)ɛ����b+�I�7���="��/��UJ�N�h]�*��-�hOV�|��֯�~��7*�d�@[�ls�	�[����<%�҃o�ۆ��r�O�T��'���>�L@酐�n7��j֊�� �V���xM�r�D8;D���Q�Z
�k#ؐ�|��e�~hܜU��c^!��g�r��;َa��3E�y�˾�xE��|z�Y�Re%��iͪ�����)�Y�o����$!�ّ��j�'4���Dl��>4<�����jbju:�i5zJ�br;�'%0x{d��fD�^��[=��+��/�ITS�vG0�Τ���NgH���t�4�>k��>����'^�Ŷb��m+�{<�2������.Bk�g��Uec�婓Z�	ܛ��7���莎�O�~���n����3�*��aKT�{;2��9�Y-3��N,��WfC�UA7E�N��s��P���k5]v���8�K��y˺��w��u����Cs�=�s�� N�x��œ�������gYE�����������&�2*J��P��\&�r�5�i� Z�%meea�ܔ*�g)�㥫"+3!�s�� {����8Jx�KZ�z��B��0��֮bv��ԻضG�_`	G�Ɯʗw)������a�}#MR-mX�]�I��-����9���K��$-���Ρ'�yŦ�c��j�YCq�@�7,y���d�ks2��y(�"q]�ǫW�6���1� ��d$k�n�g�[q�����o��+�u�ټ�L!�; ���9��t�&yeϥB6���L�LvA�<�����+
��l.��J�q�Npw��7L�S���;&MJb�<�e�tO6��RZ�<���:�,�Ó�l�l+����ok1�+qj�����,ڮaan9}j\mA����%�#��nxA��c������P�D�f
su��4)C�L*"��yv�p`�̳��jɇ����Q��/����渹x���⸂X缨H���ٵO�ڥ�,x���hh��K�W7���ƕ�P�{��UR���1�� ]�q��u5ށ:�~��mK��υe_�bP��L�Nr�j&/\WƷ�q�gǡ&��ys�C���!��Љ�I�M������d,��udz��j��~��[��z�]�|3�V�Ib8��'R[lRX�k*�m���@�0o6��OwX���'5Չ���ۜ�d՝j�\�u�L�0uͣ�1;�=�	���o��|��eٝ��[���H���]��`�����gG!�+�ɋ�{�a�����v(�����rO<�^
������8'�y
�{�z��ļ�T��9Ɠ�0�X��T����j�{�?>r�>��:�kծ���)��'ih����67}��"*X ���j�UM<r��z�\�Ɔ� ��7Aud ���"~���Rp�+�+4���#��ԝ���9N�F�H|�}c-S#E,MD҆C'ܪZl�-�3j��֙%�4�:��8�l;ϲc��u��jk�elU�>��I�k�d�c�~�����WMU�Y.�(�8�]�]�������n�M��v\."���=J�n�}x�(2����8��*�oز����j��;3��.���<���r���Qhv�pYkϭ�h�M�R��1���UIm�zJ�g�����Zԁ�Z�����C�Y��f?}�S���c}�=���\Z,DTVc
vN���X�EŖSk���Yϣ'ܡY��88�]�'����#̆
m#�S����t�N��Θ��ȧ"
�ǚ�����ѵ�/X����uV���(j�8��6����J��Q��,�N�8Q�/�ݣt-|�W.�x=pV��lb2��2�Af��'���d%[��5ǵ�Η:7��.�\|F����3o-rb��� G�y��Q�q7��|�~g�� j���DޏG������n�R�Oa;�֪%�3# �u�v�����_CL�4��ۜ8�64��um8�^��eXe55z�UAd�Tsr��0ZV�K�рͽ>Cs�i��e�kU��l��Ťݕ�1�	f�>lH����(�niO��mS8'xTݘ�M���ݢe��Pa��X��qH�Ao��]��s���_�f�&�|r,)��F����*�5-Z���\Ϣ�,(}�����69�R4���и���͑mG������<wV�Zy%_ޡ��>��^n�dMm���	c??Z�-�\aQC6��9�v.mv.���FA�zx�[��3��>%�!)�����t98-���������7Vc=��{�s&��`�[]V��`U��	�ޒ"yBa��k��1��R��i�qO�Qc�r�_��&�������7�&F3*=׃"q�P;J��9C'�	If/E\�e��P�qE�Er_8G+p�n��V�jR��ס�^\���/� �˚�s��M5�J���W,��x�u�g�����x�����z5�#`!o�>٥�w�l���a<�N8YZ�p�]X�.]m���u�w�����1�8/Y��y�Nͥc4�a���Y�j�1x����2�!s;{;AڿUKu<��ho��W%�5��j��Xx��٭3-�s�Vn����H�������Si~�-���1`ʎk�(���7U�mʩ�]�RP�.[�U���5�*]��d���yo���hh��/����\doS�`p��#N�(�+_�O� �B��V0�&����c�u���`��H��T\vOh��٘��}�!S2U;;i�j�p���)�4%@�Y#�U�#Ð��x�������XWٽ�y;�:���]W��;�����2Fjw�ܮu��}��z['�vX�!��Ak���4�=�T�����6KA~����dȞy��Bۋ�y5	�_OG1�����cQ�f0]�t=�,hh�Dט�&׭�z�ˈ���T"���U�vWz�`%Ja��gO�о��m�Īj���{��PE?ǌ|ytL6��4�p8'l�0�6.7cJ|��C���ܫ��sQ�.��;��Iq�q���妄m*�碞�:< V��#�mG	�*�F'Y��CZ;*����t�^�^�V=�ܡ�ʢ]��/�Ҽ���`�t��l&>3�^�{���������}C#�e�<,�;`��x��$�yp9���3��%�Eo�G����{T2����$i'�%��<c��2m�-P�A�n��N;N��2B+��}g ��s�}/h+b7�����V��7������jm�B��x�vW�a�߾f��1.v�;���H{l9���F�H�1��qz�w��`����!џ6�':��א�]-�n�pQ��D�{�3������V�ѱ뷒!�x������+��/���}��L�j�=[ն�T�|�����I���V��4���gm[ʪ^�97K�P�m�
8�;ٳ�"R�2��-ȧ&;b���%���Cx0�T	�",��Tu�����R�+I�j���ԩ�<�˫����>�aRW��u���[~F��5xb��y��e�� j����z����t;8�*��îl��E�PI:M,yGj��k�Q�Ze��ˆ��r1��fΡ:�_U�]:�"c����,�eZ���'b:tW�6�T�%~�i��Y-�ڲr��&C;�=��l�M6~��?�g��q��u{� ��0��.rL��<�&�s�G�%����A=hY�kt*�fQSYB��w���`��}f���2���n�t3J�<�ҝJWO�q���m�R3��^���B�&.�����sI~>�d7�ٍ1��!�}[��[I̙y<�h|�Pm��{�H1(4Vqr�eۛ��K,�ۺq��e6�-�X�ÚP�q�G�u����Řo�&�3V����o��Ƀ�6�>A��)�}i�x(��ݍ�y���Ӻ��ј�R��+G+�0��,�3e��Fndܻ
MܧY$�}��E�;��ѷ��|8�,��a>[L����k����wâZ�#я틑<ʹ�'3#'*n�s���hÎZg�׭>�k�r���D�Ӎ�0���CLS澐��%�3(�m����3͘r���&:S{��A*K�X��t�����cA}��2��1m\�E\�c�.���#��0����P�58s�᧞���y�Q�ޮ+=SƇ�ςw����e�5ȷX��S�S�djvy��ZGE1�����v�c�O���ɀSb98����zs呏p��1R��[ϮhD{a�H�Q��Md��N��@̅7�%;� �������:�8Q�Ї&��?{��3�zQ*�Z�������5�@�X�O�5lk_J����>�S`]��1��3�"Ѩ�2���z���Y�}Ս;�D���Rp�>�Q����+�5]Ǧj���)���M�S�C���
O�	�W"qѷ�$bʈy�<�`
(�8)eC�Ўi�9��%�b�0�S=��ޚ���nuĨb�p�1�ͷ�AVl]�%m�:�� �$@@x
�\a��>}U乍����v�ݔ����q|�v:m�����u�C��Cm�x$9B ݂"�cI�;��3>y��W+�R�㦝cHY��;6�,�*� �n�t��J��u���y�!�9�A��9���BwV��-XC0�a�׋�8��.��]BEE��Ȗ�~�.�&�r���Qi�׉\l����g^8�D���n�$:�/�
�]���P}�%�;��$�J��V���`�M,A��vxnwپ�!5�h�W�{�L���ȄB�i#I�k�f_�6�j��Zq��V��,�J
|r�/:vT��(]c��.���Yٶ�|�Nr���|��V^��ӹ�ثR2� 0�^Y�əN�u�8N�NH��~sލQ$��WfA�J�b���:��*�%pW�����)o[�����ŭ�3ZZjf��C��f�MF�<�Ng^,eM3����mx�5��gK{��{$��*��&֛�$޽F�۾�W�y���Yr,�]J#՚���*��p���&[�I�blLN]���������	�"�c5*��iTً��Z}�:�p�=x���Qx�zE@[Wvަ��[ՊPԃ[vv-t�LsK�H�[ud���[�[13x�N۲�FWVRW%��|��`�Ԋ�����y�KB�+ؒ�u�s%���E�F�.�GV��\���t�|p���	�J{ |B*���]���b|�U�=E��uN�;:��^9E���;9�wӯ{C�7��@x��f�H��^���i��2���gS�h4y�s��F��;Dέ��B�� �ƻ�( B��(>��ݧ���X���5����˝{9�w�������3��e�㇫�as�����6R̢�R�U��<�xKJ�n�uہn@p��y�+l�N���ke(�
m[X�@�Ւ���\�HۻW��Q֋-�<�����Y[
΀���d�ؔ�b�]�yc���d%|s�wvh��Y/�*B���/���\�+@��9� ���\����H�	�|�5VqeK���7����>��r�6�.Y��']��`�N��a�H:��4�[Crn����S�V�އ�,'�����m�!�N�75�S-CW�2{�Ǩj��}`q)b��v��w�c�%�:����.mG0t�x��IV����2�D	��wG�a��sn�f��]�	�P��̺��̻ø:*��
;1�Âʌޒ�/M����3\��S���a�����l��|���Hmf7i�7Ku,�l��6+�'c2]m,�Y� P�o���7� ��m"H�,�a�MዮN�&`v�������w���/������nW'���(�,��B�42Q��ڞ�w	���4yY%:���	�8u�21,�Y��&�Ε,��V����Ԣ�t�Bl�j���[ݽ����v&n�h�*ɝJ=�|��a�B�躍�	�븣ڌR�����y5RL�	�+t#�O�]]�:����+O���˚납����G5�\����{Om������:���@ :v��|�:���}���u�z�m�g�ӆ��s�QB�z��uV�.-��ۋmE(J�5j
j;�r�{��u+H9�5|ܵm�y�ʂ�Hw�l:��ug!F�a�$5[+H(�Sem�f���'9�VJ��6����rgW-Efշ�����7&�C���bC̓��Z��9��P�U���u���[ej���ܶ���r��mՒ5�3ec�s���n[ulܶ)X�����3�=�ô��<����e2nٯJZ��Jv��f�Λ�Y�_B���̰�b�d񱻊$�cZDj^���ٌJ��ˎ��a�(D�y���l5ڽ���Ȣ��{Ǘzo��K�g� ������!టfST�.q�!t�n�r�<m�=�_x��F����}x�x�[���[G0Gd��ګ{i�\)\@(�n��=�'�����b5ZM[mx�~��X�OmI�J�D?}�@N�����}���X�����Ƽ��vk/�K#
7�y;Μ�O�uGC����v��_�����F�÷܆�BzhB&V���b���Nޑ]�ň*9:w�|�^Gk�]��@�wh�l������F�-st�p��7y�F)`�DKi�T�������n��囓�Վ��V!Ƚ,�W:֨{m�@���w}t,2*C�+���(L1�bE�j�Goأ���>cT�O�Y�ʦT4�{<�֮��F�,ZȆ!�̝��:����Y�a�a��?t�|��}��B�Cb'M�����{��lO�!Ô-��%�~s�`T�^�;c��T:��>	���fE�d�a�Y��5 ���s�h`�B�O_���Ykh�T���t0�Y��k�ŕU��"� ������76�"cӒi����𬖆��&��6\W�{{]�5�kZR�xz�޷W�6�u�L���Q"����K�h��0��y�H���.�w-�{lIxb�y�M�ļX�olk
�Z���Wv���
�M�����H�6�[�mu���_*��Fm�1c��6Mi��K3u��[(0O���
�*�ʇ(���8�d���7ms�i=ԌU���՘^��q��w2��z��Ҙms�k��{�UK�-�I�*�� ¾��j2���4�0Q�ii���j<��&�#��I�,^h�iS��e�.��ɱ���s��.3v������I�s��9�0uCT��HWU �y{�`�/��j41j�K&��U�G(�ʌ���Uc+fɸ���E�
��3-�q+����RF��>,K[@�tIǝ��Ι5/.2n�GUč�\k��;���.Sxl[,{sVHR�׼�M	�Pa��c�b��O��rԏj���� Z��d˄�Z�='<@�B��YX�Z���z���]3�0�)��Y����uF�c��g����Y�΀�PA�⨵��*-DR}��*bɐ���[u�!�䈎hC2�N�ΦGKR���`�P!
���'ת-�����.��{��1��
9`�|�It/,�?H�ש[x�zY%�X�c^l�np辉yNT��z�[��d�x=Y�M���(3|�e!J9��3yyYwuS������q���m.��XK�tt1���T�2-ҝ�oG�wG�*n�FN�(E�)���r���v����"�u�l�۴��� �Qm�gQ)�P�M�x��V��L�S~�r����g���,!��
zܛȟ|<ߍ����t��~�%����̤���$B�/B^y�{q|���E`�*�ă�@����,��7���p�+{�ƒxӾ֬�ӂ:�7��u�P�|�hD;<��e�k������.����#�}yN�S7)��phcu�i��EsׁQ��*D-"q���%�O�eO��|e]u�~B�B�zC����〵�����A�zIa��SI�&�<��<׫}�;������ڕ�ʕ�"�;��.F����n�W���Nx��� �b�JW)�M	���:��t�K�n轞t���������>���Ql��k��y��Ő@Q�.�m)ɞ���'57K:7.^������SQ����=�fbi��C�7���c<�A0�f��W�N�Q�ҁ2��(@_w� ڝ#�}��ɏƲ�>�]K��x��:�k:ڱ�7V�}��;��r�QE��VP���c
j�q�SG�8����W�~�.q*ߦ�N>6�y�Q�����n�n��cPvh�6�=,�O�rEbS��jۆ���Q9=�Ye6�Ec_:��@�b)ރ�-f��i��^n�/;���jh�]{��|a�ҡ�ŹLCC_'fv��i6Eg?h�eJy(�KPh�y��Wo.%sǽ(-8�8n�kk���������nq��m	�//X��a cِ��z㲜��j���%��[�ڝ����������s|%�3��,�o�Y5��M�3)?`*|�+�^=�@����N���
�i��ͫ�+��@F;&u�m�K���d��ܡAD����y;3Z�}עmS�`^3/c�Z������cq���S"~� >��-�<��y �5)�}%�̘�w|�8�\+k���i)X�(�xז����D�<�������?�~��Ⱦ�n(TOY�,p��c)mU�5�ÄZ�a~H�dp�a+a�Z�}vxZ�@Lâ���7�����X�yQ�ս���q�xɇ��Az�σ��-�EA�<C�[<40ZWl6R���F�Ś�Bf,�_�)����ޮ'U��O���t�3"Ķ��}3�0��b�|��������R�*�Q|D�7��1N�Q�i ��8�&u��<Ϗ>�RX�=I&���F���[S�����F�ކx�6E�p��Ձ�lڌKu���ڸ�8�_3V#sgo�_�
�;W����eV��P�����#� 6 J�.(	�����\@��Q?߈��-����wK�s�>���d�`!g���1J��f�t>1��e����M�i��Y74�b��9ѮǎZֵ�/�1�@G�W�]\)P�Y���#3F�X���fțG/Ou�b��m��z1b�
eu����T~o->;�wS)�L^���y�]�.ߊo�2��H�&��j��������Sl�S�toa�,���7��}Q}���.���=ժ������)UBEi��a�t�J�8��c�Rᡶ��c���ρ�l7�%�/�z�J�ݭɾڍ�0֙ɚb��T���)��jBm�U-6sk!�Z�˹�i�l-��H�~�a�c�N*mc���É�����y��aM�$����e�f�پ*�şz�dt;FϾ�v8����j3�ׅ+KLJ�=jω�\<����S�;����z�h�]1rl�wIUT��D�ؓK��_T���c/�:K}q���ʆk�izC�:�C�Ud�{"�ݬ���ݫ�8�dٳ3S����)��T"����Ά�d6��r����S�r���l��/�"��R�����ڟ��(VtSBv�<u�rAt;�83YPDSs:��V�D�k~#�YM����'(E*�=��	u��;^�E�s�~wx:Ƌk�a=�R��������؆|"zZ<��k{a�e��B���6����s�0Z|��]����퇰̚�n$M�1T�2�7^5����n(3zl���b��A86�;�0q=
�.��[t�	l�I���/����c`��p���`Mu>�ĝj��'�Ⱥea9F�׀�Pd��+9L��xp��_^���9K��6UѶ3�ps�z����`6�i`+��#�~ ƕ,`@��B�3R�;5�mR�A5Vӂ�; 8̼��O���PFθa�C�`��F:��i�8�dy��݆��e���E�n:�死$��ΰ��'�����pOAq��#/����4��3ױ#;��槪$}Y=��A���q2�t����G�����^���CB��2���P�үwDV�L�`�2����r�v�/�+��#�6�=x�S�Vs���+��_.���׹�v&vL�Z^6߻K���W�^º�ǐv���y�$D�(L2Y�Ab1+2�}����K��{��Uy��˾��'�@}�M")��mO��&�m-Q>�N8�O�Y^�sM�(���(�ܻ˨��M
wP�q�I�FA���5�;��׿�U��S����m�aY�@3Kah�\5� w*�l��w�S���l��!�<:��Y�4�H�襒�SOU�5�Ԏ�W���$L�5o]Z:�RuρtRs^Y"咊�U�Q� �5㐪|2=I6�
�m`:1�)0D�����͋�΄&�"��
�o\ՔA_��䃪���4���4��1��q�]��uNo���VJ�SC ��Jr���K5��5��K�n�w+a���L�yYt���4̓��&��f���Yn�\!��`�92w�p��qK�|p*ǣ��.~�ܖT���J���%��j�{^+kQ�v=�A�1��Bi�/�y���ۭ$n��Z�#b��0Ԝ5f�Cn�<(������fy*��-�ʠSA4:i2V0�v����K�ۦ�A�l��gØhv����"6�L	n��[���^�1�n��gm1T�ݏ�������I2�F��`���K9(�E�F��w���WT 肦�h�������Mg�"<�����<��q+��#�`:��'���*�r���*��ƅ�T�]�iC2��!>ִXb��,���[����#�;�29�X�b�%�a��ČvqH9�%ȵV��#ag�B�euckM�3�S�_ʿyx��8�+y"~8�<R�^N�����Z��͸���5&��`c-޽�y�T��P�/^�|驄^�R�8�a�ƶ��J8�C���C	M䑔z�ذ�ޛ'l�{��`��Жl;;����QX�N����bj�g�9�zi8�����32S43xH�(��]�Mp&9�%_�b\�v"&)�?\ǎ�{$6�J�[�Ꝝ�"�8���'�!����vZ�:���_�p@_^�g�{�u0�%�ȸ��Ӻ�*�;}�7-	�A̾ƚ֌�vm���'2]�s��/DE䚴�(U���W���#}j��m�!��O=��_I/�,L뼷��������P����/���/~����*�Ct�J��n���.��S�7��.jo2j7{)��v02�dK]x.��y��o�<�>�~T�3��Jg�b���Әx�qN���j��oZg�W���A��QE�����aMC�C�ȿ������Dk��z���}1^�Du�=ψǧ2��֗B����Zic�=cн�
���&U��-Y�$1�-�e���ʘ�� �e��_pBZ�/o��-�Kps2��>D��V���a%�.�&U�H�� T��#Ĵ�cwu9��.C.��C@�C4��T���"��ą�Uk-s�ЕV{��6�v8�
me�+�=}6&���K�a�q��1��3��A��i��3�sCm�d��]�������'C�6H*N8�	AL6�	���]��d7��Y�%-hA�G^���o�UΗ|�CP*T8�R�8W?��44,s ��8ArX�Y2�n����8�Ӛ��v��CO6�R�}U7d�
�,�>��u�_)��sT?>`�O�C�8GǕ'��}�S��--x��mK�".��;��$S�������hV���]��'2�|�Et��i7�	W�[���Ɔx �AVU�GI҆��)��w�C�Y�ʭ�1�n�!��.��� eel���l�QL�tݾ��؏Z��$f�:�Ѿo���st�"b��`��|�ש����E2��M��uX�*K�P��tU6�{��~&'-�3Zd����t�
�XQLqHp]0��}q,��"+����8�5<�N�rNڱç�0ؚ�l;����X΄g�:W��Lxy�?k�)�a���6ڜKv���)�гv����L�
��`G�fxO<�r��8{�����_���F�� .� >�򘹦�cKtsk��>��r�bl��K[G��Sa���(�Ü*Y�$c������U���;4n&.sv��,*�tׯ�sv @�<2$�O�h��6K�R�:��lo&J�e+����p��3��f��&=93Ck�+�4!����R�f���4ͫ�r-nQ�9U\és�Vmv��'B�2(��)�m3�pVY5��zUcX%K'���u���F���q^�����H��@��mY�M�����5_��Q*>�ϾJ�kd���Be��#B��.4л�%�tUeB��msȹS�{�v��sc:����d���+{a�f*'�&_�~ϒu�C#vt��b�I�.�tuw��.������ʠ=��qU�ݕܖ�PT2�Z�7�I�z��5s��RߵX�kz&��N�EHC<S�cF�9��ӑ�p�F���iby>��v�j�xV���SƲ��g�Ǐ|�s�����k-���嚙-�Ὂ$dJ����B��i�ށ��`��t4�t{ USV�6+[g����H}1��4��ሤ���ܠ�P�+EBv<�ih�f��M�T�v�U�5K;{dM!Һܲ��Nk"YH�T���bt4�:�3'~���n�Z} >�n:Iiݮ���#J�������{N:�� Ğ�Q)?��S�k-��[��Տ����u�t��)ϻr�)7�y��'=?&4� |�ʀ�r��P�lݚ����b��0��,OR���̗��_l�wM4}����h.�
 q��4�k2�y�6[C��&��fQ/�t���P_R���-t��f��9�� ���q��S�hs������{��Ew,-z7�MĦ��֨*bgX"��1;�(B�OF"�C	؇l�xf�e���D�Ne�pJV�T4�G端���~�͇mT7h;E��n�pZ��9��E"�z&]m0N	q՘��˦����>���^�`>�4��׏�终v�f�i*l�e�cO�[Hw� �(
���;��/���`������US���T�b.3��|�ݦ���)u�pˣN�(v����:]�g��4�ӵ�^6�a��ij4ݖ�]i�ҧZ[�[���=啭mkl]ݝ�4���c[�b�POLQfYC�N<q�֋��o�;hX��eu���j>b�BE��xmN�����:���,rFI�;��G�~-Dm�@(2��t��.�k;����eLY�Ts���	�V
2���Y�����=������ƣs��wG���*�`�W�.l�̫JԨ�����ݒ��XS�J��hL�:Z�gi�:���d��>��s�i�����+k��ހ�ʢL9x�p�D����+�!a�3�Zó��m���͌]�{��L9l�#��$�^[ЫTZ���g�̾ر
뜣�5�{b�͑R(]�́#�b]K_&�oU�*�4�ۚ7Nq
���Q�2�b$c����T�$0X�p�+U��N�\�#t��/R�V�6�'�������+��C4+�`Zʵ�맹��]��[w��WZ����P�c���AMp �y�,Jc�Ȫ�*�l�9��	K��s$7ʟ)B[�9���s@Wh[�w�4\kGiteG����iS_-����h����X-�4���ek�Íݒs2�Q�ƨv�Z)ʘA�O���sj�(��gM����+].�tr�5�zyiಅ!@���i�Jt���6*�N�t��z��,�v�[ͫ��1;��ބ=���G��纹�T�c���.��r�gc�mЩ|'ϻwX퐤���<���V�-��Vq3��ݘ�&h�T��0����� ���b�{��n�*�R�+�V���WÎ����¨��Tb�kq�ݓ�^,��Y����iPY�j^Km>�����N|(q'�t��v^5���{y��V>�ݛE�6�8��U�%���4w\��Ybܹ �*�dd��5y��Ioք&���^����b��w2��guJťi�*WR�p#��+Ŧ��uH�%C�ZA�.,�4�{��ʬ<<���L--Q2�63T��KŲ��Lb���9��J%ې�Y�Nǩh����q�}��oo�����J�:kҎ�G����eȮ���N׹�j3��<�Ձ�ü�ʳzM�n�p�s��KR�eca��P�A�EٽL޹������t���ϰ��De9Vviw�uӬ)���Mh�p��Y�t�J�x��'kA��9G���\�;Ʀ��fr0�]�e�z���]ţ�ǡa}V�D��dmі�k�{�,է��vW��ώoy���rhx����79f����%ݦV�^*���Q�]{��y�;��t�m�D�mfo8L]iK�WEf��\ކ��N�z����K�ȓ�am�;��v�;ܫ�/qT�Ŷ��T�u��:S���T���M:���-�ݻ����q�����(���6u����e
�7^�u�[9*����c���:��s��f�����l�uumW\�ܶ��Vڶ+aՎ�L囓�u'Sucr�ݎ�u�g-�7Vܳ���g'����Cr9��Y�g��,��u͵nX9�6�x���S93VՕ�^-��<[gVM[wl�V��mJ����3|�ỳUf�z���\bYusŶ�|mݎ�6.�[�[��gv���1�m�<n��u59ly�93��w;�ۖP�U�@���؂�}rfz�[u�T��`��6��8gV�:�+�@S;<������ʾ�mMn�ѓ+������,�N
~< �ߑv�1�n��o�/�5�a�Yl��W'^9G���>��+��m�����.�n\4^�;�6�&��|ǐ�H�#$S,�=���'�;�Q���3�'g*�.��CSf��Ԯe����U�S9���Ц�v�v	�!EM����Ss��%�1�ћM��]Y�d�QH�הyc�
��oߓ�1V�*����hI/}��Q��e���N��:h�f��e�~*,�,�^J���&;�r	��1@�&�aWvn�y���$G��8Gf��v�� ��Jxqp��OI�ߒ�K�Ŵ:�l�ґt�ykB���lA���	x\�%�mE�9��˽U#��)���=�6�����r�����J��bۦ�h�bI����z P�ܧ��w��A5_|���s��M$=uH���U6�t=�hz9��:�sǟ���7��#1������Z6<4:�����4�d��g��z85�,���,��Q:;	�}��琒�>+���N�U�z鮬���J�55�<��N�MW'���c2�l��.������ӵo�Q͝���)��4�e����S*r�r�5�_S�\�A�[��.�Я��#aLhN��<	�9�oz�V�B����^[}:�k,�S��SXF-3�vA���ik������\�l�F���8hcu��g�S�}�탣�0� m��V�e���g�p+�;Z�B�$���:���j��597�;�[�{���A�.(���ћ�o��-T^�Y��NK�,(���� �xX��f�8v}�{3u����;`cf�s���fJ�[�oǸ���n��CTK}@&&����G��X��vf8���}�K�����òG5�+OQ�3&�<�_�ǜ�<��"�rRxi��z��Y�9P5��m������:�\�/D�A��k��p�<��ጻ��G�"�DY�s�30j�{��[+uw�ɶ��A��j)>�+(V�6�[q\�<���σط��Brk�f�eV&<�^�dg<�ʝd���}��M<���>{\��{�H)*����0��O|=z�g�*������P�5�Ma���(�-�2j[}�	?G�l^?<�1�n/F��/�b����^���F����O�"}e��K�������7{�J/e����˧r�]�� 3s2�M�N��a�k��e	��������R��=���ح���c#�w�������W�cUkO�QDQ��{A��}4��˃����)�%���v8��A�3WbH�Jm�-����'�|��&sT�S5ȒմzX���־����>��rx�����O�׺�a�bb��9q�I,6��ʄ^�P�>Pgo�1i��{qU�N#;��fW���xW<��^4d�e���ra�<ْ�c\6��o��Z��Q.^�=�fV:���оM"�_0�f�s�Ԁ/<�k�V��o��?==BN��&ds�A������ŧ���>�4*���;7������\r涞j�7��E��Y����Y�'������F�[צc���GOQoW���(��еU��Tt�H�4�T��7�9h����@0��a��P��:X`���t��+,��\h��䬣�ݘ=�gb:%]p����uL5��g��'~S�d%���g�����?�>���7��V�J�K�\K�g+�ɮ�L�!�zqj)��T�:��Y��D{a�ȉ�8\T�G#UmY�\�di�N���F�&nO�f�G"�S
�.���EڢC�-��
�;����� �ˋ�}ĪGl���vQ�����ݽT��9nנ� ډ�y{�U���T��.�\��(�����=���:��[���V�?���,�e���$���V���⠧5�(����Gv���P˩�`�%�K�N*U�S\�˒��mQO9�ۊMZy��ڭ�'BW4�������6Y�5���H�$���8��a{3�b�/0��|y���^��<��D��藹��Bi�ګdpo+�-�:m�RjU"m�v((Y�Y�����S�kv�L���*KL14(O"��H5,��i����J���������g`�uP����w�������.U�R���v�BU�y�)�+$�Kd�=4X%b@r;�f,C�w]�Gm"�Ț�%�.U��2�G�z�v�U�T��l>uA0��6y�^#0��}�MsO� ���F9���]�'xG�W)�3m)���=����)�y���<3��H0�a3܅��Mf��`��t�{�!��E�y�*)��"��j:/yB���;s�u�(v�dL�I�+n�\վ^hw����^wy8����Nޞ�b�W\�;��J��At[G��P\\�Z�b5]aեI1�k�#w��%٘�q�<(S_%.)AQ�ؠ����(Lcڗone�ι�jt���P]���v3��x�A�(KA��23f�f��w�Hۓ/��	�	H��edk����G��e�6%�P�#x�x�CcK]� gQyQ����i��k>2�U�����qQ40�3;��@�gEnr�?]5��!5jo�g�*u���ڸ��l�� *2�f@�kB�sS��+8�̻�Ѿ&��Es�K�u��:P@��Sgx�O-��,�q>˚]v��q��E}k2>U�q���ה� ^dG�:�����M'X>��ۅ_�s��]ꅮ4�:�'Xe��p�9�eUuT�w���_���J%���9��&F7���'z)�L�<�L4y�܋��p.��]�>\T[G���4M�>�Fd`��֓��=��!�o�n�^l%�XJ)8r��GPyN�.�_I�|��,��{��'b\\x����m�^�]y�=���*�Vw@�+����=s᝝��qz�r�fp��/�����r���15O�����/��ku�S^�R��O5Ί��O\o��#UPD��it;�k�vL0�g�$�	��#0!�ʣ���~�MW�������)���������^{� h����W2:���
�Q�\C5\	r��L'�;9���*�~ųL�Swu
b�z��A�6�LRsϋ���dP��QVk�ۛd��Y{����"�Yh�i8-�2s#�C5��hcZ�K��R�쨴���^�YV�Z���}�]e���6���@t��6���������u�=��9-O�VlFjQ����z/�iP%��0
!���E��bj���ߗ��FM���	8�^/u�[U6��`A�æ��#��Y�\Uy2m-��(�+�����[1��NS�:�d\�c�"e:֘W[���P'[n�.�Ι�,V�*����^\�
��c���AikU�+\�urۍ��K����ʚkM/�	WBk���h�,����y:�N^�"�=n��anm��e����q�z�x�&���$��#_lew,�|�ч�?_}6�n�|�.!W{WK��k	�AuB�.~
����ri3k�$a9~`k�G0�B��R�΋�9p�v�MH]#1��8p�6�F���U��lsr{[���O�1�_���p'Wo�ޒ�ϊS���[\�yq��U��/K��1輏_W~&u8�	�kM�3<�
��{L0`�+AF�2�������#l�L��Y̺�M�ߖ|�i)�,ɦ����6�.�	��#�c>��
���n�/<��0M�a������ס���"���\c]��/���|��b�	�����wa��X?˛�๪/�G��Ohl�yB}0�v{�x�����m�p��Q��xVj��7���-� %uN�[_W?�~q��ߘ���.V!f�-��Q�2�X��t<Ԧ�ؔ�V�A�N�B�n+b�����5mAs�����,����:q\߼P�m��ѧgE���,���go�ÝQ,x�^���sX��󧮼t� �@�;a�zi�ڗj�{�M��^�eS�FFi�n����u&DN�͵»�C��U��=(�<�*	�\��NN�آ��5k?�����;$�o�n��?�u6µt,5�邃H��W-8�(4���s�Nٗ�䰹�1�8��cw��2@�>�� N��4��:]
��-5i��YB���qHC����z*L�3���0̙�����1c����I����L�-nfQ~ħȔ��MhA�)��FM+izC��U�(��נ1��KH|�T,Y������y�{�r[qW��z9G���~C�)�_���υ#�5�,O<���_�xgѣ�*��(��[胧������a��R����)��R�K%0�#l�a��'��uE���ra��T����D�=�����Uٿ|z�v�[tv�e��
a�Wƌ8�f�s
�]<a}���3i�`[�7��S�U.�Ih##����֩����=�}����C���P^�j;�e������Xp�v��Wu�`����F���-ӻ[?���9��2���z^B�lf�X%�� <�-G5ŌV�E*Y�%\����͍��P v��i5G����w��t��[u��j���E(�5��sk�x�W�ɡ�M|��R�N���ybd��m����X�^���Z#�ϲ�/A�])}*PMn�~F��fw�2�v	kORp�r۹\��Ɍ�h��Yw�f���M�m����vt=6Q���FW��{!�J����r�y��5Yyfj���ź�~�)�5=D�������gǡ=RZ��k���@���_zٞU�i��xG�R;���ܬaQ�Ut�o>��e�"��;Q"�lS(Ks�*w|�!��;�[1��E�`�Rv �WT�Tu]�ܻ�IM�"��w[5���V.���`�9M4'�����"[x�-�pԞu;��K��RA���v�����xp+�ʦ��5�y	B�"�&�ګ���u�1(��Sڦ�˫�\Frb�6�4%��h-�a�&hmbS#E{�4!Ԡ&� ��X�,�l�+��!⹚%܃�J����lQ4(C������;r��ɯp�u'�@㬷M��*�O!�s]Λv�R:���q�M]
�bڈy����n�!Y�)r���VKtgR��D�;I����6Z0��,���J�e��t�mWX�ɁB�\Pwƍ7.�S2�ٹ:	Bm��S�[6b��Z�=B�;U�{/)�
�U)��*��Pq��&r�qm3戶�3���/yeZ��=3��)�	���@�����(���oꈮ:-�Y�b�.�C�C�bz�=Ӑ����e�W3�pnq7<��N]����Y�{�zOc�Y�f��ڵ��n�q3�_^E�KQc��n��,���q�an��b�q5�o��z�M��x`������CV�sK�P�3n��I����<{&"�T�6�W�D��}J�\Kȉ��Of �]�D����߭��=\�C�O(лTm$9����O����޺�22-Wy)q,�YOf��}�;6vD���E�T�:�ݸ@���K����~�a3��&^��~�3���s4�F9(�w�1���s]֩㉵��>f�UV�"�.ƌ0nc" k@��[
�pF��$Q&ߢ�WK��V+�R0��t0	*�ks�q�8϶��Y�&+��5-Z�p�w3�,�� ���z`eVWa�Ќl�^٭��#Pbd`\o�=�yt52w�t�`ᬒ+-6�+�5������$ )0���+�D��Evl��A�{7�S�X/�(�0.QNX�e�{��x,ʡ��j�ЏF	��¥�����(&<>�?q����#�Ba���j<^Q�Cq�tY2�g��՛��07�]]tԱ�~��^�c��MzL�:wTFd4e=ET�٬{�[�4���8��\��>�D�3�m��I�2�n�x�!�m�B��nG�3��q�e6\�����Y��D�����^�*�yf�M�%�5᝝�Ĝ�o���|�o��|�%�~�F�.�-����֨�����,"-}S��̭��}Kы�Vݹ�ֱԯ������60��oLخA'X��Ҟu���Qv�dX�n�}��_iq��E�}ۼ�e?�_vag�<	W�ڢ�E0C�<܇��Fj��3j-ˈ��~�Y�}pf�=17��?��i�]�5z�\��D���"�!��uF����z�)~�h�E#X����2S'�Pd��n�4�����^M��M	��K[�h�S��"�)8�8�����`��~���.&r��Y\�zs@*���]N�x����=��j}��h�5'��v[�\e��Nt�J��a��H_f����^��<��#�<���TO�U��?L�`���s��tl���K^�>q�{m'8k�6�5��н��Q��F9$��0���`��*�|��`������Jo2�+S}��{���`���nj�sW/��]_<;V	�6I��������`�e��ۣ���nu夺J��l�0��ւ��Ϟ�D��Kv9�}�F�w�&m�Z��^m��x��� ��tLV�|�e��q�q�jq��P�+L��
����F��N�K�W>�o�;��,r|_�V��D��#	�Hu�k#�g���s؃�C�1t��� 4``1N:�a�5�$lc�Z˙�}�;H3��ݛ�S4�A�Gtbd�9�#��W�Y�޶d�{}��XmC|S�7ljJ_e䚰�2��`3��κr=6T²v��U��2�ʻ:u�x�l!�]A�P˝k�f7.��xc%��<VI=w������QC
��Y�z��r����{�x���MV�^_�d�;�5��l1>�qN�n���_.L���Ӈ�w.+.ӻP	�؈�8�k�]=�����zp�º�m��Z�zr��6�Z��Ε���gI�U�/6S<뉇��ٜ�Lgl�(pf
���`�17ƳhG�J52���ͪ�J^`Oo��P
�+7�ë���gp�˴x�Si��s�L�R�^.!�Qf���=ҙ��2�C6�>��尒�#jP�]B��GծM
��\�[�+���\��v��#�}����o����ҽ�U���hUkF}R���o*Kz��,\S;���W��&�x���D�kj�[���g�����f'Y�ݜC��n�	��U龪������|��|�Z���*X�ג���Rlr_q1\���%�+��%v$jV2����NV'd�FQw�m�kֺ#4�.߶�2n����K*
�|�ѴݒЦ�����چ�Lh�&g(nɾ����r�6{��#���i6��YP�gSƁ���7g�3x�V(�(��i|5l�"�dޜ��M3k���w1)l��;����T�g�wK�k;�td�{soo�萮�	CC�:�Ҥ��,{sG��o�o�L��W9���;�KN5L^�)ඕu�F=U������
+*lM�7������л��R�Wk��ܸ���Et�>Hp��*�^�v���F���3��U����;rǸx�y]�f�-�v�7�7r:]"�}����4k=})|��tՅ���pw�uڬ�)��vQՌ��H{R���r����fv����y�H����h6�<�A��ʷ���m�F�ιͅ�6�gg����%�6M!ӘDj�pD0�[x����1�����L��.�*�8ټ���EZo�n���e�U�1��oY�h�E��@���d�ݹG-Ttf����J�l���j��e��sV[��
�JvCx��b���l�(b��}�'/q(�:}�m���wtC�����C5��ЇVd�Sh�������D��*�I�,˻�}���V��$�v��DV��1�D:&�9y��ٷ1�E�'m_`
A�7��I�{v�mYMͭ�m�;�鮆���]���N�z�\�����0�~xL�e3����ܫ��XR�����S@DQ�o�{�P� �T��,a1��w#{#�}x/+��먇H�,�B�]���s�0\Z�fj�D)�xW$�^ԭ��w�MM�͘��&���%oRU;Lȩnp��>wC��tU���s��M�6�񫙠�ӓbшV����92S��r9�98�h䫧B�]j�/�5عƭɄ��̭�ͷ�m���V��wLrٝCn��ܰP]�r��rٹrڵ6PSj5lՇ�g!��۫r�nY��QJ6V������X�g"���F�ܫf���M�ՇQ��.��r)��,r6����X)���nY�z�r�m�F���-�%3r7#nCz�:T3��B��j�>nY[+j��՘���X�q�ʈ |( C������ͶW��z��v�Z���@M���;0U�h�cu��Z�­�um����t��p� ������<(:�����4$���R(���(��I�������*��͗mc۳����~�h)]�v�R�-��:���{0���Ox=�f,:3�0N�Y��NϞ��CQ�c��CF�]Ս74�=�}D&�{�[��q��#�T�0�ڢ��>��c]u��)�E���̄�K��QN1��v�l�ʪ�M�0�)�b�h+b��]^������I]S�T���=+��F!(Dn������6�5B�8�2��=6_�d���0�®f�mQz7j�;]
��7��!�0zQ�x&g�������.���s���O(�z��VU�Z'+mW���G(�<B�qȎ�a^͇l�h��y��E��k�Q�*�`�o���C�C>w�`V�n�9窘^٤��Vj岷�+$ל�vX�sG ��p��/��n�.k*��ϑS�:�Em�8�uǐ0:�I�iW]6TtU��i�޺3����ɟܘ��0�Y�~>�̕<���U�����7AEJ�8;����B�ߣh��MXaa�nx�_��S�D���J�a|�<��)g�L��9�+8�v�|���� �!����q6ړ�]���Yц�'C���nWS۽6�T�s����|�7+\��2f�)�kΩ?�����<f���{����0�&jDc���òd�c{�;�O�W:ĕ�2�D�,���Z�g/5� ��g��ߩ��m��Sͤ�*��,Ҟ`WG1��s
N�Ϭ[!I痼���#q5&�=���@5F�út�&`�6*=���6.��R����j;�e���Q�S�O]�Y]�gU����z����̐JyA��TS)��-�,{�%�+8mѮ�-�z�-��u��2"���_��=�S]��u�D-7����џ�^dV%ye��O��խ_d2b���݆���t3��ͭ�}M0u��I�_3���Xg��{�7����x�4]c�� :�&b�~�0,�����%2�p�^����W��3���iBc�v/���_,�Ml�{]��̕/[�S�{�Pe� Ԍ�`ܢZy�9���	���ƪ�V·m�N'�m��Y��	N��c5龿��3������0"�Uc�z^4�xڸƗ��r�+�Di�ʍ��֙b��Cq��'�4h�jP�a��, E��3���6��w�AS�cȬ똇�zw�f�����P�L�󂶲kū�Ucx#��uAg��y��$��t��Av�h�K(�̡��t(	jJ�S��y�5tp�'��d�V��|7�#�z��l OADXJnəd����=4	�t%��uw0"Y�S��K8�T,����;՛]:�WZ%�pt�*�:�S����s�#�{�n�js��F�dP��%ymynh�%i�1-��f� n�na9P��QDfUfI���(ɤ���W�U1Ns˦�k֮�7#U�D�|&��:��O���#憜A�B9ׇ9Ǩ=GE��J<�L!�l��^܎��`k���3�[��N>w�ݼ��.�︩M?��	�&���-A댢�Ү/��R~k��@+���cx����v�����0pW�;N0>U�wtp:#�[�P�\����LP�⫓�Q���,IP�K��5�V5SѤ�'��}=�i���in�����m�ndd���"r�*q�]�3�Zjmd��A�!�q��)��}��;C��?&4�w@���T"�?^�m�2��W�����e�n������|�p7-J|���%��!��wlyضƕˬ\������7h��i8��K3`ӿ ��_y��#�U�0�ɚ�5-Z���\Ȉf�M��cs�`��ݻ]xr�5hb.��z=�o=<�p&2��=:]�##��O^"�CW��������q�ׁ��j$���r�Nͩ[�U&ݧ�n�r���d�3{nst�tP#n���5���Ks1�g]H9��� ��s+��:�)6��Ȗ���V��:'J�: M�3N��tD2��Z��"�q�_�x��"��ۈ��0:�������`�������'�:������A{��c'=C��4���f8�k�ZA��-7}
l�oe_p�^���ҩ�Q-1&r������4K��EϴC]\͊��#���C�2L��u�n�;�L*`s����Y��M|��4�A��Y�s�+����Ɵ$�{
���9���δ�b�����a���,�%Q"�mˆ�ON��d��.n�1�R�!Z#��m�������nJmz�����z5Q=4y�]-"�H�u��F%Qbs!NAq,�Z��I�^탻�!tźo'�w�wmC`�&�h+�'ɊN��tRs~Zh[m��U���.�:���u#\q�\U�"'Ry&�ƨ#'����mF����xR�ߊ�O�t��8l������f��\O3m'�6mE���������g\���#��f���v�䨵��TZ̾�P��i���":�r�N�Za���V�Gw�\��:F�m�l�\Ze��E�ޜ�����y�[���z<��go;���A?�s������M��Ipp5����.��w�_w��Z~X�`{�z��iޡX`�܊I#�P���S�Wy�p�KX%�XW���7g��ݥ�<Wet]Q�y.�G��~�$���S�N�����1����ֽ�[R�i��,x��\��.oT�w�͠u�Nn�i�7�z?������uya ��0?��ߨ^ӷ{Ӵ�`8h�����ۙ"����Y�M�tu�|_��roH�l8�-�d�P�A�j�Լ��{�=�:7��yB}呡њY5:�tKv9�}�#�FS����y�AWz�U� &��>���-^`p�����}Ӧ�X��㖹�m�#!�|��^C8r���X��k��l�
X=�D0���F@<��S@n�;���������m�݌c-�H���%���g��u�W�]k	B6V!C]�T(��A0u0�a��&�� ��׹>�����8�4I���M�9�{ۮ�� ^,��&]�4��SP1��ť��ɉ�,�O����|�=�c+g�F��WT�9ctK/Jj�SN)��Ţ(�bQu��1`Jۗ�˕~��w���W�-�(7�p����o�k�ep�������-�קh+�3R�2�
��'ˡ�T�ا&E�=���7al;8U�]��tn��ϵ]"�Dmu
�}Y�X���,z2PeO`���+(Q�.� �Y��^#�j����܎�Ӻȑ��Ðֿ@�J�|��P
ɧ��BE�:�фp3gd=�_i��`�=>�5�c��C!+��S�}@�(�Z�"�'LY�SW36)�=��\������R�9��.�f����2�G�{���-��9͌:�9�*`���5$�&`�mq�����O\�̴��av�ը�Yq�D�� �Ko������E俾˾��94�����V닽�V�v�z|�bZ|�g��R�(d���W�7��-���g
"�}C�=��%��z�\�j��9g	i���sE�&��[�0r˧K���JD�c8-Q�z��-��2x�� `+9�G�<ʺ鲣��t� �����am8x�^v��$lҀ׎�<��v���&8Ԧ�6��-�kƌ��
�K:}Lx��YG:�'��v�uClV֥��j`E�y��ɤU�FY�<ÁFK#�'�O�9�pS)'I�^,O�\g�#8� ��Y�����_�h�BR����|U(q�����w>5P��ND���M��[1�Q���P�<e�����3�:��3�ب�Reu����T1��2뻧	�ϑDd~����˯o:�$:s�x_��W�����
~:�"�٨��G�n����U��8]��E	�kzF���Ԗ�b���@f����מQ��������=���GY�!�&�1B�v��Kie��v�}��O�UI��KC��h�46<� p������n�ݘ��8�of��&z���=55%'�wB�K�H�c!~�vk5��Ax�Q�����Z��ͧ�3�Q&���ϛ�h�s5��Zwn[u9��v�#�j�|��c@x�H]�;��@�pj�X�����vjݾo��6���߆}9+\T�JO���j�A��~D��\��ДPa�C��+���y���k�{��28���!����g�1BS�c�3f���0�����QP�m"�'	�ћ���[�1յ�������tȽ��J)��'��@c�y��"��۹)����)�Md�F�7�jk���֘��c�EU�˹�6�&�x�!���C>��NܣҎ��&Iݽ�]/W*�`�)��O;M��q�Ob����r���W�(�+Lӽ����9pPcz�^W7�JsP�]gt���Xa3)�s�U2.qt�mWX*22㺘�|f d�=��֮�K�����ڨb�X�� [��\������W���+��i�!Hx`���u��F�I����<���y��vB�����.ʒ���/�z��c�,y�+p,}�i��}p�<B�}d'�l<�0+'���3���c\`��ȡ֞G��}�-8���:���Q//:�Gw=f���A1�)��v^����&���!�0S�EDBn�LCn�E��	�pF���ȩ8����kq�ڇU��{y!�Ǉ���^^�V��m��O��L�
�p=�8o�u�W70�d ��lS�fkQ�2�T��(eq����Rʁ��Ɇ��)y�g-`�`<��5ƀ̌ʇ^N�u#5F4�N�g�ts��K
���^��56H����~�T�+�@�-��+�3�< ��	���҅��\�*�uE�E�]��.���T��E��e䔖���^�w��o	r;Ha�{��o;�tֹ��d���w ���f�Q%Ay�(��ӽ����V6����ao��~�8��#n�V�Y�󝉆�r�d�m	t��5�0�i@� ��w�H�����hc"��8��K�^S4�C�5��v.=�U��K�#�?�g}a2u�`�d�{�@b'=3��3{�H��7���SY�-lƪB����&o\=�O�~�ZbL��U�f<��qa��Oh�̙��N�v������9��[4��u�ض
{���بCmU.��qKKE����~�?zV|�+�ɛ�;z�o0�&'��7<���mz�W4�k��4Zzwx��&��9�0yCV:��DO2��&U�I#rж˘Ά^�X��S�W	���ʢcr��U�1ˈj,1;�fmZ��*ÍZ���4�_L�m Z�
�v�����<��(�+L#��Eϒ��A��)5��D,��'��d��uWפ��*�ι��"�����P/�%m'U�!�f���j��1օ��hk����J��6��O�(1���Ga�J����o�mS:F��}=��z����'�NZ3;����;t����t�H��/k�$Ρ[@ꢚ}3ryG��h���o��>e;�P���hdpe ��	��*R��2��ߒ�NOe�[-����,�K���1oM�I�ʯ3���,���k��R����A����õ�^��F�1�*�y�F򣍩���|3�u�i�p��[�Md����Ұ�Y���cļq���ܹ��:�2/��L��&�>���af闸�li��׵яtD��*;��q/>2������,hl��~���4�mo�v��q=M�	Ev����k����Z�B����,0���ɉ85���{��vG��m@�k@n="ķ�i��m1�O*�����9MO�����&���θ���>����p4s>�Y�8dg.�15���!#x{��^7��:^'+��V��c��*:����2:��d�#o�*}b��N����;Wx�w��Xܹ�ZA-aq��T�@�m3�/�b_y��uA�D��5�5�q�U1E��k#UM�:ꬨ*j�X,�a������fmţ��L�6�Ä#o3 �乇��s
�P�U���L�+x3��N_Ӧ]+ۘ���T��K8�oj9|�Ow�[<{]�'V]lJ�V�,�;0����2��~[�_~U�i,C7�rHZ-!v^�N�6�xݙ���R}����|����8{�o8����r�Č�yM�]n��8x{���e��;��XzZ᷈u��r�>�W OTzjkkR[^:��Po<7�V�H�ˈ3�l�)�z^�l�z����©�;a����
�ۥ.�vz0�v�&�3�c�ou�9<N�7E[bk��m�!!�=d>��K���dKeʍ���h˪�!�fqH�훉U���2�Hl���"[QM$c��<�6�֎��JnD�u���+6�%l�9�{�ۙg�WwqZ������/Y�ײ�V�{@2ظ0:˴�K�����[{��-����$OV�ō� _V n��b�'A�!e3��7�捥Q����p�w�]�_�w%]�E0�����\8�� D\��n�X����s�=��U�'�5�� �,
��_��S�jπ~-/g4�g�Yz���0�>���F�Kpfv��y1�*�]Թ�I�b�����v���oJ^U��x���ِU�j���^���%�j�c{p��sjZ�q6r2v�8:yI�۰G%`b����jw2��e=�x�G� 9��*�C��5�^^K�<��*��rF���[��yv�9�+4>����M�����i#��_��u.���oFqHvb����c�e��:ۇ*�0�l����-���Ԫ��[���^���&��</o��W.	�0;�i=�K�^������&�utW֎-�Vs
,q��^��/��S���j�r�j8��҉ru�a�c{7	�T���\�n��=;������F���\2�J˝b����2qO:�>���&Z�4CJě��)C�s��`�P�	fuC{��t��Vf��2�*Q�L��z�<�k,���~T�Ɵ���ko����;���d�(��;&���(`Q�,�9ZUi��:*�R9�%ԡ��)+*b,��OUռ^��䆞��8�c2�:�n�H!��q*u�t1dn�r�ԣ��-�un�Y��J��Iԁ��y��{��y�q*�٣x�quڧ��̮�a�9]�{-:�n�(P�qo0z)R��A3�i��j"z$Tk�V�Z1���𙟊}G�2�a9�M�u�5P>���DS��s*5I�0R�)�OkIQ�[�u/�^_jD��d{��+
�蝽Ŧ��k�k��)Y�F|��Cwc�5M�eu�W��'"We�]q��1�[�Yq*WZ�a�uK6;�'pǒV��X�N�P1��U]�O�t35���wXl���*�/e��x��>�/Rd��@i��[Բ�'6r�g1U���K���-޼�x����ٮ�}��黷���4�M����*kkgQه]o�r�Jf���y���eNX��	�[&dH�Ȩ+��΍���ܸ��62b�^:���,��(t�f�
��f��Jv=�j`#aO]�7,}8��z�ܭI�&��s65��ˤr�֡��i�n�Ӓ)�����KWm��"�n�eءR�&ښ�ƍ�m��,,�]�q�����Jf �W<�^�67OT���k��)���|Y�
�T��l��><�r�<�^wd�����YqUK'6�Y�iN�LS;�EP�"�ͩw�����l��(�U���(��[��r�i;�x�	Ve���0��שGO
��Ѡ���z��+����I�r�� �|-�^��3,6)�q�@R������	}Xj���"��A�MW�f3c{�]�EC7{JƱ-W��u�v5�'pS|��|o"��ي�-XhVd���-*E������{L�A�wt�,�9�z.�:��)��o.�D�����4�l����Z�v���5zz6C+6��O)wn��γr��c`��5��ю��;Z:� �go2��v�����ڑk��f��pG��A����X�q�$�18�}�}着�������LH�[5aM����՚���V�|Ö�ݷ/p��+
ͫ5V*����jf��L�+(*��jj5jjj�-�\����>u������(5���'%mM��Veem��WQJ�j)X�(��rڌ��-�6�͎El�����7#)�P{���39S+5AZ��Kj7�9e��r�jVi2Y��V�ڶVVSV|[�Vd��*���:_{Ԝ������W(wVu�?vP�w͙h��wp{X	�s[����F��׼���r�0�����`����/*&�����O57a�� ��-!����5eF��/��n���4�L	�����k�5����E�+�'�Xl0�iS�V�/o�\T�
��6��oT���#��Kx�4�=o>�y�?im;�싆�߯U�st�R��F�� ^��øv���cQh��)R��O��'멎��'��li6�/�&�x��"&Ѭ=>�O�)�x'�r0.l�T�MY��f�I��o+6����h~7L�dPv��#J�D�]^�Nl�N���9&CE]��0������L�~���iԁ�إ�2CrO�:�Ժ��匵���G�}�	3ڗ�J*9�^��n2B�y�n#M�wʧ�}MtO�F0�i�#��#�^�^N�|�	W�I�륓ʮmQ745U�{]"/����+-=Y��2O��5�����F5�j����5o�YsA�h�)�ڛe.���U���2��s36<{>��$�A��}�&��+�7?)ng*<�D�]s�]���,,lw��[�X��5���iۂ`$��wo��RP�!j��r0��F��nVŹ��;g{�7CuZ���1�kU�F&�l�9���<��U���R��_������Ǚ-*>K�p+�3V���*R�iVK4��]'1�h�<7&^��k��ٜ�� <��+�g�ŶD�o�|Y�z�6Ч����^�#�o \��.M~�̭�]34�0����:݅���o]��\�F�s�R����s����3�b��s�n��N�O��a�$2�0�d��`��%X<.�j���֭�\�F��|y�QZ�Wr�Q��-�96����Ù:*�_����8�݇u�cUP�ue����'S��xH�n�k��㏨�Z�5
�8%���6^Ϡ3rcϺ����_�j��|s�C��Fq��Ҥ�mg��^�Ƃ�0!Y�b�b�n�(�-f�Q�e�^E���Ӓn��g�*#l�Xu=�\`)�A�0p���/��8�k+�1#.@�l��C0�p����`��I��%ֻb��������5^�<�5)1#�7��kĿ�G#8��(	�.�!����u��Sgs�u��i�ɨd]�;��U�	'?���V/z��vQ�ذxޏW������1�53�c�fؽ�v����y����W0�E�W{�vt����M��`7H� ۃ����Kt�9��܅ʬ_����]��c��։�$mt���٠r�R(u6*x��l5"/V�Y��v�8�i�%�$룈;����M��%!�UMJ�*���«��X�������l�	�/j�N��M*΅��E�:UE�,۽ƽ�����F��wޭv��D5\1���-R˕�:��r���P$�8�"k�
�nOH����F�ȼm��M5��7�minK�/	`{Oݷ\/xE��3�G�M�\��l����S�C��0B��U�̯�H�c��Ee��N��]'�螲�l@I��N?���6�H��`o���͝w"�C�m$n]I��WD����34D�f����hsx�J���&��p��9>e�!�N�u�ٱ��l����ʙ�^�5�j��9η���m��s����u�7SctX��Z
�Ԧ ��ƚ���V�[Φ���� ����ȫ���<�<قʯnS�ZA0��\�^C��N[4�L�0
'k�õ/lp%f���#��67��,�-�'k�*�x�O�`�"vI���)y*b�/j|��:mފD�r����)G�\�m��&����>�O���5��ސy�ќ�N���ym���3S/�z�`�7&��=��W�{�x�q]%�	�m�I�X!=����F��}�a�{ڡ�8m�6#"� Y�>�]tgܶ����xɞq��k �������-�������������x�����1�c�q�o_f:��>TZ8�_�y�qn��U
��t����J�#7��r�nYIz's�уfE�k{�TFO�5���l�ӈ�Z��
�v8�k�W�<m�w<"mU^�K��p�;;yE`]�lz�j���2���RN��M����.C��*��f��=M5;w�-��'!��]�|��Ӳ�\�]��y��*�F$U����j���79ͮ��8`���@�;�N��CT�P8��¼��n�^22�4�d�)�E�����TC8��e�T���/pM0NX�6�R�����3_���@��"a�vcř���ϩ��~�3��J0D:c�VR�����sR����+[�w�R��w,M<k���S�%ϫ�RZw�;ȳ���m�`���s�|���%Mu�,_=#�%ԮM<�1bU����"�7��y.�뺾i++2�T�h����I��m�N�8��|C�o搸�h�����~%l�9� ��mxKd������v7_Q<�:�}=��a�!�
=�]�@�䯍$o��-���F�ڕzЋ�TĎ�ͳ�x��kp�)�$b�Y��z�k�E�'�Eu-V
'�M�.ܹ�6��񭎭���51�48l� 7oO�>�G$�}ƨqI�i��-R���{�޾-^�磤��K�kn�}�|b�8 3h��u���Z˳Yc�sXVf�,�8�=%�0�Ϸ�GQ�-š�$%�4�Y��m5f�	�ƻ�E�ɵ��#_�{��z��Ơ4!~��Ȯ����~�?]s���������,���Ÿ��[������|^C���U��3��FNM�]q� ]qT�/����*�g^���!?><��*�����/�.�=BbU>H�m�|��0����j�g��r��V?D�-�W�}!�|k��6+Gxξ���z/p1�bk�m?@�YkV워<O�j!^k@�,��Xc5��͵�J9�E,�A.�NW�����=���wݛ��خ��4��͌���-{�&�Y���O���
�{�";��fɕo�1�]j��i��L�t�׮���!��lW.�J�חXJ~��W=rO��5��*�����f��3s�*�z[ij���v�jN�7K'�\ͫ&h,��k��ǌ%�R�,�ж�d�͓�r#�اϛ<lt%�R�Z��3K<Vd1��9uvw'Y�-�vp�a�8@m{4�"]XC�i}K���yX*��Sw���n��t�ז�	��2�o2y��LO�d3�,��P�{�EO~��Y˦������>���E#�JU��a�V�fa��pޟ\�L^�q�-Z
�"�2�B[���N�n�crN�����n�e�D>��[͑U=A
�'G�Ǭ���ĽZ�TWu�ݞV ^��-���+S�ﺱ�7c�ٚz��6��4\���Ɂ�;�|ueYֹɪG)����F7���� �7�74e�>��/ޭL���;pP�`;=�3dj9�[�5���_-�)6��N�>-^ �K�N���WҦ��%(�h{�h���;9Im����$0�E��W1i�4��Wf|�������x��ҡ�wP�C�&gnSK�:����ӭu���˺� �B��i᥼>�5��z`u�ܬ�s�'����ۍG9�}u��5�9W�ж��N`vKP|#=�3< ?";r`,3�`V���b�oh-�$ Ԫ�eـ.i���4NTq;8�Hܗs��L:�bC��<f��E摝���q��o�~���>�|/ʳA�u=�!�#�|���6n�8���9gN��<n7�F�:]�AD^x�,��٣ܪ.�wV8kz�0�'95@m�k�GA̾�"w(��n�{8�2h�"�Su��F+w����;Xb6���]Z2ۤ����O��ˤ�eM΅�|�V�悮p���UӸ�NĻ�U���D�ބ��,x�UyrR+8�9��v��=��BL@��ɡm���z���h��*�����C�MnSmpݵ���<:ɰ�5�D>(Ȟg>���=]Ϸ�{^*����yv����d-�W�0�:�1���gt\t~y,+��E��VDp�=��kbt�!j;���z6X;�&/�+_\ˠ�/N`6�n�9���#YB�V�W��zn�X���gU��$.t;wx����I��ͫZ�D�ݥ���SkSz�;pښ���۲wR�^J"�{eբ?�}�����Į��V������so�l�VLuT�d6e��F3��4Do�/'�͸��$�oK��(�lݶ��ˈ}�u�Ga������t�����n�#��=����ҧ�� Q��
��㌗�4���)�c��7%ua�@��aX��wC�����oF�#�5�
[�j8���-ܼڙȌ�+}���Cg�{���v�ŗ}X����z�mTGK���$���g���{Ty�8m�p���R�����S�$�����p5�^�:����w�A� ��3��g�0$�|�G{ߟw�n�>ޛ:��挔"���7��N6�O6p��=��s0ka��<iQw���
cݻ�[�ϣ-H���`�7vL�7���c.�䤌PSjغx3!����v ����mi��x��Ԉ��/��V��SևD�#'ǔہ�or��%yբa�M\�Q�y���v�ݾ�W{�Ԕj��&��\{x�kn�K3�sS�ž��n� ̱s׆���G[�*���W�Le���;8~%f+���2���z5�pKm�k#�W�H�i���)�ӎ�v<ǫ�M�!a�������n�I�O�D�����k�� bj|�j�������Kbl1N�v�s7Dv廾v��|�|��S-j�}��<j��N��*��ZحM��Wq��p�w��i&o����$z�)]^Yu�U�a�Z/t���u�~B�A�VkT8/a&��m�Y�r6zy���p0�6�H�W���/ٖ̀��TR�My[ø=�LŷE��XC��ƮH˘u��>�o`KaQ�~�(A*b9��vq���:�;��Y�u�)νt1y)�K�����679^A�{!��3�2�t^&}�t\h��ϫz�ߥ�	��uծ����U_�=��[��5yTz
��M�����^�ޘ��I��P�0�C�^!�jW*��_�[χy�$�,�p�jn�}�ρ��Ù����j='{e�oynw5��GA�H��Qi�Ki��f�;�>c�p���W
�]}f%n���4vr� �F�4`��e���LF��s���:N�Q���a�W�\fTy�}2V�v\��w�Rkvܨ����+��ڴy��bahz�m"�#�����������1���36����gZ�����-TQ{��bN����n��7� W+�������iy�D3�!�t��9u��Y/Ү�el�8�ӑ�"b�h�n�wn�����$$��V�B�m���3�nm����v�r�/TV�ט�x����]�&��7J��s����U�����C��i���f0��M�����1�́��Me�ۻ��.���F�-8���u#`_C��(�WK�����~�3K�9�bZ+*���;@�&�[C��ޛ��D�w�M������  4-��&�vv║�����|��t,��-��w�Z�,W�Ղ��-�u��n.2��u9�痭3XݯB��!�V��q�L��T��p$�)q�A�D�^� jd�L��!��0�\�+��A�zZu.�x<��9?�,���]�w���ԥW���Szm�y\��r�_�����x>���0��4��J�L�:�������n��]h�M��A���- ��*G%Ыo-;���܆_Y{�Lq����7F]�GP�
ӣ��B�]�X�XY��G��v����ə1��F[�Ɲ#[����C{�S
�WX+	
`[�R�.�)��h�4h�ÈS-P,�!N�)x0WA��j3�fA5NV*���z��fvV7��ղY��b�å��V����Փ
��V��LO��"�e�F��4��0eҕx&�ay�&�̋E�;bř�č��p�;��m;�N�}7����5¡�b�h�c�=�+0�2/M�[���:0>K%]nڇgI۷���I�����-9�k˽�o��"!�c���q*���b�˖ye7�sI�`���H�`Ɋ�=���x�V���{}�m���+���})b����&����\]�W�/�pu)8�5��8�cMVҷR�\�%�<'!�a��&Yi+xأTv᎖B6�G}�`�ee���2j֓�(�,F�c��л{N(2U��%7�;$��^����)*yκ��1���z|����e��'3F�U�W�k��b���]f'B�W,��JZo]cݶ�R�U��n�̘��UK�M�Ba8Mn����E��#�e��뻶7�(���2�B��Q͡B�m� W8.�6Luv �#�ӕ�o�זn�Bw��=��n�G���ge�N�f�!�>�g,,[W�1�:�5AWG�_g%lv]� �t� �ǂ��Uu������m{����V-�$�
A'w����gf��.�j*D�:e��x�8�˘��F���N;pT:*7��kTm^)��^윥2	'zWY�bM����{�.
ߣ�`�L��qJ3�z�&�8mE�빎�b�j�s�Y:��q<Hz��:x)[l����޼@yQbgY�X�����v�P4*����Y�l;	�
mo ��S桭�ᛶ�ZF����jm%M�L�)i�|%�7�J�!�c��e��t3��l��������vi�B��l�c���i��4�oi��<v��yC�W�֧�>���z�n{ԧ���'�*�^�ӥ��V��u7o�-a�Zu��L�fJ����57}��u�ha�]&j���k�91l�ҟ�K`-]|l�L�|)��Ҳe�����Z6��4_Ҟ�+P7�U�q���0,Ѣ�a4�Ke�2f2�Y0� �r�6��_jv&��v��خ�VK���eç9��PTF��܎��e8ʭٮi���tM�wW@�3��iΙ9,�����4S�T�v#�c��>��Û9�] r
N�g,�	:ˬ;Q]���&��(PoLke`�洉�\$�����&���hi\�WWF2�j�H���i
$�vl%>����=����˰�Y<È���VRk�KY�(���x�8�R18�o�Ѭ�T>����N���+QY�b�V�Z�V���}m��ն�M��'!U���_K7R�S55em���[S%���Jţ+�9l)��J��SQ�x�9mZ�*�����n��J��+V��VɊ���$��R�R����-����,��qej���6�N[��EP��ܔVo��\bFVڱEj��[QZ�j}9�lVڱ&�����+c�8��Vڪ�Z�Ԧ�ص53�9�̕a*���p��z�f�I'�#�.���*~�Vp����
r�s%�n���E]ۥ�t�R��;b�-O���f�>Χb��+��ͱ45ow1QK�JݝGGo]����5x�Q���g����풕�a�7V�g��5.�}q�y*XLƵ6�D�9;�={Tr���@�/Ir��w�����Q�y��n�i�����Uf�*l\���}��o:D��:��|K������W�J����&�m��&�:^ks ��Rb��N�f�%j�s^ۉ����Z����L��?i��R��֨��g�E�Cjhb���2ʏ>�{W'䧢ە�~?���������Q���&F��}� q��B7�Xd^6�|:Ca5��d�t&��L���vvSXq�ٍ��D1Sn�Y�Uǫ���I��)I�x[L�`s"vL�����걳�+n[�[?��!��
�c�Q���+LzP�fUs��כ��r��N�����ښŞ
 �<�5S5�]�����Q���BD��_L�>��֜��x���է�������2B�u9�� ��Y���h����1I����C(���߱R�Ǔ5��t�d�D3g����QcU	��]7�Wa�@He�"m�4���Wjy��e����H���q���v˄�0���4v���iŘH:��p���Y{F]�ˎɂ��ț��z�[�v�7��;���wVo�d��X0vJ�=��j_y�l�wy/�yd��P[M�#\Dyj��[͎��|
&�&2��>���ދ���=ʲ�&򊋌̧R[L�ϡ![x�mi��h8�V��TE�.��Ɏ���L简'����yK.��^D��R2��p�M�x,澺ɮȬ���`��"wOu�H��y�VYWVTv�(���0��\X�y��u�kE�g�z���Y�o�t.%�=�7Js��!0���6&3�l6k�\��O��H�$��lZ�v(�4Wq�uo���|�d�ڴ��z�C���[Ztٮys����j�5�f��/�У�~p��[��������~�fN�6ϻ�͂[C�7�s��p������ْ+�v�6ټ6�;Yִ�(��Tz�}��"���%N�6ʂBŗ�F}���7�TsU��(�.��eW;{tS�j�od��~7��+�o�=|*N�93E�\���U�>Mw�ާ$��wQG�a��Eم[-��ǣ��}v\����b�8�M��$hi�ru�����V,!�nf.�����9��rw1}�m������{�X��x��W%!�ˣ�->�ӵ�#�K@s|0�#��&���0���LS���8^613��z�t
�S�u����P6dκ�T3�H���T��;���^�6~���С��ʑ�Z���$�Ѻ�>L���g���5�r�s�܇(/��+\�)���`e��P�$����Oq�R�veq�MV�G-�vC���:顏*�=1�عxʴ�4q�Մ	��2�Ix�d��]�1S��SjI���3,5l�S�ED��g�X%L�p�|cf:hh���f���9c�[Bԥ^���U�8�o֪�d�DM�Oe��N�E���i�p�����^~�=л/�R&��ڹ��[w��y�"���ә!����2�n%��ܝ���{ɫ�2^i�xJĬ�Ⱥ��їx�=V[-��A�橇\�mڒH�˵f�U�4��'���lB��j����7�A<+o`��wU6�ފ��^���fI6@��.�o]���u�=L�>kk88*[]3U�ݳ�&��E�p�<[ۙ�Ez|z�^� �xXw�z�y��F�uǵ���Ξ\q;ے��'���� �yg򷻪�<���4f�s�ۯ岍X�����L��~ܪ6��o�jѾ	3&OZ��^vjGwVI�� ��g`�a�9<�� ȍY�qL�-�^�OR�;1�_y7���ue��W5�I����6��[ݔ�=\w5[����`�teΕ��+��V����꿊sݞ����f2���A�ڑ͸!�z;X��SZ�ޓ!�d��#ǲۏ5��d>�<S��yt+��t��٫�0r�Vf�"寧Vǚ���5s@�*m��I�n��Anw���׬��f*�j.���+��Ӗ�[y�����/�b�v����fu����u��r�F��t~�������Z�d�)��VI�x�� Z��H��-p1S6�*��7!C�ήG7� �?��l�u����q�ux^f�Cp���\�.��/>����,�w�Bc��^��/>̹̂�Kf�P�9��q�M�����/w�m�7� �巖����"0�\>>�)Z�U��o����PX�or������	௸<�*��8gkGl��������%d#3:T��vTu^!.31nEs1�X�+24*��Ih��)S��6ą�P����'��^�Pfm�u���u8��ж�()�+x��Us6��2Ʊo��s*0>��9>���CMC*9^�M�i�J�^`��q& ����.����d��-jW&j7�~��a�~�e�`�E�z�e�.���G�X�ؓ�׌��\�~s��xﾥ5lԪ����Ɓ�<��eq���՚a�#z���y�5��5lE���E����}P��n� WPe���΄W$�&h�7L���ۮ-[F����L<�+�m��s��U����ZF�SȇT�&3^E���:#�e%ZhL������:�ܱ>+hk�ٯV�tc;�b�b�v��o`����m+&w_:oy,�1�k�4�7ˋV�����?��+ќU����u3���!���YƫRf��N�^{��hh�/GJ�;h:���-�wLb.gqi^���Nd�]̌1��o]M:� c0�܊��rW���1|��_�B���\�����c�!�c����E�T��#Os:�C��O��E�"l�m���#F�Nv���S���u�Q3r��j�	��(Эa��6���W���L�Wؗ�>sm<�,T{^��B��:�6��-,��7�I�~�Nf��#ts����#�R�^J�qj۰�;�Ƞ��!桖���s<�����Ҁ/2b}�ŤE�<�$�PU6��z�F�⺶�m�ٓ%L=��s>�È�Nc� b�P�J9l�|�H�N��PxV��u;i���e��J�y\�&��*�CQ��;�48��4���^�����&r�gD��o��T���5|m&\�o5�+�m�t�����������ӄ
�ίv*�^U���n/���G �MR��5pL���Ӓ6��/ZJ�xK,w�Me[H2$x�Ԇ�b��Ļ��9��'Z.b�{��7�s%Ǽ^ViWf�iF���Q-I����q�/�;p�;D�v=V�AR.V�4{o���W�.=���� ��yFxO��_����s5��k���<��]Z�v�lKL+��T=��^�O���=��:4�ٍ�נ��=�_���櫩�)�x�Ù�)�ڞ���(��}�f��2�)��03:�Ϝ���vo 5]̻hp�y�^�fۻw�I�F�	t��Y��ͨj=���:�[����d��T�uθ��֥=xL�\�V�i�f�C���d����o���ښX�#���5����zy����V\<�0�����=�25��U�]��Sl��7Fm�t�b42S�q�m����O|4����#M�'U�/Ң69Q��+b�Xf���u���\)�w}ņ{{7�^�$bΟfqy�5�z�����~�O(��'�c3_c=��]>ޜ��ݍ���FfO�%+�V# on,�͜p.2�
�TmTTD�ל+N����f�/N5�:���*��we�4�Ԓ>E�sӼ�����������i��TL7��E�g톰���EW]^-��S:�Gv�c%]G�3�6�Ͻ��G�C�������L�{��˜M �&c�*'z�1{��7Q��+J�ww���"��jn�ҙ�D댖h2]{����`K�Ru0vY�y�F\�s����J�\̙2q���[tdjf�\�2��y�%.�����+�Y�b�%��|�<�Z
�"RuG)�i#�f��F�]���ݳ.��k2��qx��S[D���.���C�L�5�a�.��SC�����[�4s:Ym�1�]�#�(bR��suMM*h,i�Zs ���-�^2�#�3������Y���A�s���7嵒*��}v�r|hT->5��SS��p�����5v�v�Kh��ZA� ^�RsO���1�zj)����6�{l�xA��S��[Q�t��f[7�<i��ё����'[�4�maȪ���OZ�;�f�wY1�z�\�Nيyw�'��KX��w���i�wp(#S�t�ߜXU��w^S-&a?���,�p�S\z�It�x�<wm_��>E�ζjg�q���[�Q`)T��בS& z�}���Cyj�(��zg'y\ ��)�Ӷ�z".�s�r��bժ}����{��x�4x�n�3�b2��x���ݧ�5-���5��8�fDfE��ql�v���x9,���M|s@'2��; `���M�̆���v��h�v:�������"�Σ9�ʫ�$��J6s°]:N�ms�qg�U�,�i��ڽ��Ð8)�}u��8�'o��6�
,��nQ;�h�q{�4ӵ9�qTc�ɇݧ�{���^crpN*�WB���΋>��+5J���t��x�kM�	}��}Tؾ�^n�#F[���i,rf{zL�G6c^��&�O*u��l� 5wH�"�,�@�x��ѯNrû�^�-7S����6�����{ ?�����^�(t����c}�׳�3wl��ٵ�&7���J�� �w����v�"��;�4,~��7M8;%:���%�p׻�mx��JP���*�F���d�g��)]Y����dv@T�AM�iE�|��fe�&z-C�fMv&�ѣ��5��M��Vժ����fCa���m{8WZ�d�m�Md���l���}��<����Ug���*�}�ّF�<�Q�)��,�Ճ�e�c;3��92��T�>��~�揽��%Ά���g��^�a���ܻۖ5C61�<�u��
��N����c�]����Hfq��d��}ɠs]̦���c
�OmH��a<��/5�&g�&�I�.�a[�л�6��U����%�Ǫ+�c-�.X�u\��Q���Y�}'TIej��+�R�M;�|��W���\�j�Kd�jS��H�
��ykz��A�Ӕ�xi�{�"�d���o�(���%��j����]~����`5r�qO��NY�
��jhr�C��`�9�	��m��;�����{cz��+�����s�Ꞹ�ݜ�'���	涀/<�-6�i��7*���'h��|���7K��^��mqJgs��Ӽd9���p˺c�ݤ/F�����r;"��尛�a��;���9*4�Z흎�ʺ��J�k/U�sH��G�{BQg3�6��e�l�*n0T68��8�mw6CɆ����b�bF䷛��e��7�J�LNo��]�W)0x���X�v��U%��h��0!�-�U��.�EaΠ�I8��H��T]N��N����u�jsI)j�]�l!(�3���'T5<����ܲ-ld�Ohj�M�*üg�ꭗ��r�e�ڰ=�5�&|�@�[�{@�,� `�͆h�m�m1mèNǶTu�̱��$�b ܾ�f��IC&����-Q�*��;����J���Lt8wA|�\�a\�.��[V�V4����#YxU��mJ,���^U�a���`9��_+g\pv��7��%�/ �҄�U�ѹ,qj��-�`���Ay����2�_V�N�_M��>�zL��c�¹o�t��v���fIP��l���a5�0X�X�o�fcv^ͬ�FZ�w��~�A��&���#݇k�h��pIIG:��ol����E�%.)�Lߟ�e���շ֟!���e-�ʇ� �ͺ�ԭ�������)��9'1 ��[PX�׆�u��9��D"/�R�m���j5C�7�)�U|��rkY;1e�$vkNڍ>CBJ!ע�b=��'�t��N���$�L<��GwuX,�+gN�˾�˰Е�����!.x��Xn����AU`n�gb�Փ%������}RV*��PA��o���_X��1�w݅�x�0�X$�.��fj��W�M_#A;�Cu�Y;l
�)�]��=�//��U]�݈��^P勺-�d�=(��#����5;i)�]��ƻ	�5�,,��0��n�o\r�[[V��r+��a��nS¥�z�� �c����w[�+emvͬx��ո��Ĳ��$�9�����Į�]�(�qtz���q8�-	z1q��Vc�2�d| �=���}��Ż	�@�j ��wA��ו�:���������Ӡq#��n��b��[�٫��uVl������x>�l٫ύ9���o�X}3z�m�\[�'w>H����k�7t]E�i �L<
:Ő���$�.�Z8�	��y��i[b�nL}�n%ݫR,oچ�놮���w�u��#qb�]d7[YZu�3�YfWayN��u�+J�f����;�|�r)����$�s��Sf<�� �\@8��M�w(���a	]�2�Y�un4mË��S�[��^�t,C%g����<�fh�yv9�3$��J����.Nܗ�:�z�c��L� �ɧʰ��wu&m�L�x�؂��	�	9��}υ���"p�.x����"�1��_F&�/9s\�\�H�2��aؕO-22�\61��n�dy��qG�XD�l�k1u��#��n� Y�:H*p+���:m!ٯ6� <���n	��	�EAN�!.�Pm��i���wQڶ{&&$��b���˒����u�c{�7*,ގ�ǸG.���6ae�3��o2���^&gRI]��w	��.Ҷ���_[a���-s�F�vWSWk]���S�������؍��@9���Wo�Cv���<:���SZ�xo�;kIY%��i*nk��_��X����oz��iȘ�ܲ���ގ.�!5�&��jC%p윌�f�+��D��P @udG��w$BW4����3�.�c�[��6������tֳ��C�;sg�N��[�1���:bqI��}>~��V�MYMMJ�|�+ݹ7�92�aճ�O�9VΗ)U�QEej�#Q�9J���i��B�Vj�՚��jR�����I�b�kW r)��$��U�Seeb��Ԧ�eR�)UG�8���x�mU�{��V��[QFQJʓj�QEe)�%�%�ډ眚�Ur�[K+��Z����YT�����V�YZ�Ԫ
��ݷ5����ԑJ<�Z����mYZ���s���emJ�Z��x��VV%Z���Uj�Z�Ք�U���^��|���Qȕ{Ϧ+�QӋ�Mp�+w�
�e�]N��=9Z�s�j�x�b|���Ƕ��dw1�ix�73�����V5^��UW�#��h���9%8�Ec��X�9�(�Hx�Z��Țͳ�0�9\�&K�9~Io��+8r�� �����짫����=3l�����x@�j]\�<I�f��d��~�r֕X�.63�7�itt���;~}�����W�׹��t.4]"��۩&dk�ǌ�b�v_��H�b�����W�r�q����}*��~,��.���Ʀ��{kk���]׹������l#���g�{h�����N���g�;���;�kع�in�{��M���l�������1T6յ
x^<��j��4��zA�w	�ZB��.�z������v�g�³��+;��į��lP�«W@m$��K@��� �-��������U9��>0�ڞ"�ȁ�=B��^���^�������n�-i|�6,�'\��_�ӂ_i�z�xwln���Zz�|��:v��'M�λ�;M�rsj�4EI������e�/b�3�K�O�2���NǼ�ެ�;�n��&�����"�5/s!�la�.�R.�Y����<5?����<�/��~�����a�<8dD�*1��az�-�&AȬ�]M��ʡ*-�&nfڑ��:�L�ly�Ǟ�x����Ž~���7q��ft�6xƛ��;�F�(���vFX�Q��!��f���R���U\�V��S9"�2�'	�'�9T��T1Q:�$L�պ�������M��~Ρ�r�FgG���6�iʼJ��=�u>�aө��aF�^襽�W�i���"2@��in�;λ8���-��Umע�=�֝���V��w�����U>l�ɲ@VȲ+x��rF�ўS�pe�7;�x�?P�}�0�yf_�z�	h;�����#��;^jBz���q\��{�����ǧ�� k�����4�H��L�ka�2���d����������:��{��暽b/�;�uqD����� �3��ao{K:9{zfw�E`�A��on��+�e2O=i�vpevj�i_HZ.����+������&�^�M����,��5k˖��N복*���ݡ[�6����F�Z�Ѓwu���/���s{��ܬ��	c�L��_k��U��kٜ��WS�Q*I6{2���=}����t��	��'�J�䓫��9��Xd.kn�ހ�0ff���T����=��:i��	�O]�wW��ն
-t�^���W�s��je޳%�2�^$T^עy�#��[��V��mY`6�c�SO�G8L���$�}�ʌ�ᆃ��m,6��̈
�ؾ��qm7v�v����*���DJ�b5X��2�x.����"��ZdE��X��oe�S�V`�nA�O^�IU��ƹ�ΊM&�9S�v��=�j�tTbc�S����$Q澳XոD�nc�����Z�K5i�R6[�a%��ӂ�KJ�=��p�������zm?~3ևD�R�\�yu�T���!��3h�C9�叮�ъ�w�Yl�js��*E�텚9
��Y�Y���@�8\e\��W�v�=�u�m���~�G�dکXp>�&Q�`h]ԼUHe��6�O�.��u��mVI�)Pz�!�훴��}S��LdN7�V����D�lS�h\c��w�R��K��t&Չ�t�(�#�z��9��W)��s%���ⶩ�Z;�d:�]�W|�S9X���H��f*�lQZ�f>`P� c�f>�T��ͧ���|��;e�Y�C�aU�b1�&Rɽi�F�S^0YC/	Òm���ٷfu��.�W�E&�W�F=�S ��%���uo�i�T�<m�B���KS4܉�7.4^{��d$���r:x5�����\�6/�v��r�\t�R��R�W)O�k�/���;���*h^c�A�I˲�&h��h�~���>�;��{jkW>���YaFE��Ѐ֔Q����%3?K�7���k�?�#��1�S;�w�J��q�D������Aѓ3.�q�%�_��Ӹ��ٶ�`��ϣ��ʁ��v��t��XA��g#��Яl.l�A��ƃ��0����ax��v"�`��30[�GtM9�'[{RBK 
FTJ�z�l6s�ɸ�Ѻ��y�����=����r��*Bu���+�l�s�^��>*�̲�{,��K�F��|NQ��A:����l���0�1E����Ks��{w3��r#��ñ���\4<$��'l���ȵy�;�Q���*a�ƨ/wn�EǻsP��]����/��UJJ���߽����e��x�=O_@��TYxL����'����z����P�׃7�k��rY��x?�kT{�+�J�8�T
`,Zc6Wt5?X�ϒԪ@�TD���ʎ!���14��Ji8�b�\C_A�Ru��];����R���^��:^ݖOU%�M�V�q/��RΝ�	,���"�;�&D]�8�3�!�.3$-���q<y��GN^sS�$�fN׎*�^U V<
�u,��a6ɯ�vW����A��T���xK,w��\�4���2$�ˤ��}n���C=�n/�e>�Ϭ����������se{�_��.���Ӕ���u�z�y��beze�i�T(�w3G��H텽M�-]�
)��4�18�2��˕�n|��;;D:��.2.6+t&��/��Rp��ӣ1���B�#+t�<z�ƆζaC,�
[z\�>�M�萤��5k&3��p��'��Y'Z���z�����2�qk_E�w�w��Bs5�<�%{2CR���X>2�������e����au�:-@��]��o�بl��z��ڈL�7�ň����N_!��gn��޿�- ׯ�����0T�D�	�m���}Kv���jm���y�?�C�+���=w.<&|���G�|�e����姵_v����|�zJ�2;ڠ���tm�4��V6WOk̇��&Fr�L��m�9���ņkb�'/R�ƆaŌO"�P��w�׻� ��6*�t'�/uٹy�ݻ�O/r��:H���x�R��j��y�7�9�r�3�+�3e)"����@7_�'M9�M�|��a�'��u�Q�]�#�#FL5֛�c|�S�$o<���n�4�CY�� 1U/f�6�n�ڤ�>㮸΋������
Hr��P1��Su^���� ?r���]^^Y���H%j{�gM��bn��3��@#�cԷ�-6�*����Uu^����,���hP�g��2�-~��Ob�M�,��Zi�s���r]��&�+��kg- �!��e�O�˵hL�:KH�]@̮���ɓ�Ho7��O�����[r����������m��G�g��!ugJD�Fŧ���F�tՒM�X����a�0{,y�qJ�ְP8�/�jt7�Dq87'�f�p7�����Sa�0�vgwx��޾p'�wm�q�!��$B["Ȼ�-�q�tb��ˎ���;�ɠb~�����ٯ��
��0b%Υ�YnR;\AsE�5m5��=��ݑ��iq��r��rG#j�.v��8j�π��?�/͗<�:�0_�l�M��{U9�}w���up+�$�ܶ�g�o����t�6�Tԣ����S���uK�0��n��B�~�������Mل7-����}�M�k9^
��0��w�%VT�wW��sDLS��o̍���݄6�7L�5_���b�<ؔ���Bql�]-�t(Y�����dL���K�3�f`^Ps"�3��g�������m[�L0 H���i���='�A������/!�k���ȼz�+b]�2Z�t��s���h����D�i9���x�M#�:Ά{�g�ݯ�����������,9˟S��;�ڸd�q�̜t�RӬ�qm����;�^#����*���L��psd���fLyl �@�iπ�r��>_.ްnE$�>r��tv��/Ea�-쾮�!�%��Sx�HlꕭM̰K\��3��w���j�I��[��e�a�y�3~&h��-p1S6�uce���ߧr[5��Y��z!�`=�!)�^6�'�ևA(愮r�]o�p������+r>�3I�xHs����>�O�&�MSd{|z��+���֊͚�� �ݻ�w|�8��{7���C�fz95ǩyW�q���h���c�)�z��OF�3��E���2yf�{{��~$Zw�~��	�Բ��gK�]T�f@����F���`�[�9+�Y�<�8�K=�r�e��*m=-\��82O�����X�h��l7*4v+�b섕�u��b'8�K�V��ه���_[� !�dB
)�zq7H�� q\�֣N�NqW�����U������̼��6gL:�M1z�6=���Z�)���m[��~������Y�:뻳��s9���M�C�v�댁�W�v67�y+��5��Fe�F��5��ܥ|���{ϰE[6N�g�fkx����_�=^h�����n��u��:�1L�NVY��.gD��Mc�$;�3$����pЧ[�D�H4s�����+*u�lB�����+�SB澭�[�UJ5�8MM,��5ˍ�~�2F?<�r��95�w�τYn^U���N���o�k}9��������fqղo_����3��-�wH�Ega�C,�7Rl�o�w7�z��`N���~8�H(䨓�!ֻ_akR+�J�sA\5�U��+Gx�T3��`����8�#��P��!*R˩ݓ�5�p�y����v���#�q/�n���%�U��̘�$<���xm�V����Ϙ�u욌k�n���3u58s��A�8���4���5�`�ǠJi5������4ޏ�~�&_{�h�*g�S�/������/&1a�׾�޳�G*��9@����mK��L�@k�j����ۉ��v
6�{;'voꢎqm0k.�7$�e�*�ǁV�w�'�U��n�tg��"��xtv�p[Ts�y�2�F�:�5�K(f��M�-�?8�6bn�Lnx~�v䕞a�U0\7X�6f�f�J�H��`�����	��x]9|Ydc.4xd~-��b�+vb~���Z�ZA��!���5׋	��2,�M��1�ꐑJX8��vf��l�k:�s'u�N��:;�K���S���O�T�K=LY�>�vs\��� S{��G�]t	���.6^NiV�������`�M�l~a�0�ڍ�1��-�#L������Q�=+K�l���o�&NgKǱ͒���w�.�2��q4��gj�u�췽���`
ԫb�C���Zh��ڌp�֫��޸܆��ݭt�V \{,��"�� ��[3Ըh���9�$��s%f^��Z�s�ݙ��|{Ҹ]	�����o** ®U�K񱧱e�<��m��z|U��j{��wQ[�.�E�}n�[@j�󍭑H�CO@bf���n͞�V��!jU���ct�mĆ��6@g@�耔P��W#>�:�^/\�4���G����*�ʧ�ȇ{&L_S5��d?xt6u��ؽv\�AO5�M�ʌ����~�׳zV
�iB=���/(s������������ǀ��m����m�^�G���lfj�?�8�O'Y��.���ߞ�1�Kl:9̀�006LX[Fuׁ���&�m��p��&l"��,���"�����ٺ&lp� ���ف�6�D�D��tXXL@6XC[m�� � ��0l�h��m�LXXM��@f�h� ���0m� �E�\v���&�&h�h�h�h��-���M�u�]�D�E������#6�cD�GVsa��<�����}��f`��`�`�d��������z������s}�����o��O������7��I����y�O�����=>�����w����/���o�M��~�����x��~������Tٶ���3���Y��������la����;VxL��7���m�ſ������6ͷ���_ݳg�����˦�Ϯ~��oY��?N�Ѿ|3���>���j�o�ᙆ۹ŋc
`+ ��,&fŀH�mm` l�؛km��F@,��VFMf��m��fc͘����-~}�<m��f�����6a�����(l�t�gݷ�u�?_���ݛ>��O��_\������[����/��l�s<s?G��wپ?�v�{�����~�M�Ǔ�l�u�m���7ݾ�{|M�ٶ��l�~͟���gۯ�ǭٛol���(�a�ޙl���Ks?���Ys,���9�{a��>N�v��6͵�����o�ٶ�3�S<�o�����z϶K=������Y�m��m��?g�?�fQ�f��Cf���`��+b�³l)�(�+6±����`�[f�m�V��6f��V`SSf`V��P�Y�M�SFaLaFm���ն�jc�̭�b�`�l+ḷcm�36�fS`��(�

cb��5m��f�+ff�(S
m�6��V�Vڳ)���Ƭj6�j�Y�f��Pj��+a[mM�m�m��g��>��͜ο.�s+o��?u���s=7���~����m��g���ɽ~06ͷ��,���~��m����~,��?��ѽ���,���N�#�gY�����������Ӝ�������d�Md�`�t
m~�Ad����v@�����%x�7�RJH�H���ET�)R��)@JPQT$��RUB�+v:�R�U	�IQT�b��T��P�F����[b�PRZ�ؒ;�"�ِ�֒�"�J�J�)V�IDFl���!-��P�T*�kU�Uon����ptً����Q�ZaT�&,�kM5�bDC5�T�QAT��JhԤ�� U)B��ք�(46c�a������FZ��l���j)*��*�p v�J����YITm�i��5MX4S�Pm�M+EA4BT��a�n 7���5���XFڥF��SKe��dŦ�h�,j���JkD� ] N�5���CJ�3R�m��CH��ʄ���c-��;XkF ���`��i,ؠѦ�Vi*Y�m�ڴ*�*��p�!t
,DjL��Z�e�j �mH�e 0 la��)n Z � (�` 6` $ l ـ �h*l��aD����8 	� �� ,��  k@ ! � c 5� �E%�RE�� �:�f��� `�3 [`E� H  �J =� @   5O�%*J�f��h���a%)S)4 h�i��� �&MLL`���~%*�=@      RD�h �44jiȘ��&�6���z��JP       o�ϗ>�e��۪�Wƫiڶy��ʴՖ�!" ٳ�kyI�:?�%�L���H$Ay&O�HDA�oӇ��������m������4�_[V�M�}Z����ֵ_���^ٵ�\����:N�<��n12)�x�_��-	!ihe��eF����w�~vλ�=ֽ�mqK��A|~�c����	DH��O��a�����3Q�����c�t�ɨS�JY&��ʒ2L�U�Zr�]��/���t���T^�[6:K0��&�edJ�AN�9��.ۚ��E��c-�U�҉�)[���"co0V�^EY��Qdj�u��J�a7hێ�
�y��i�SH���u�$�A1nf"2K��q���	Md��k����p��jB�:��^��4�����&�5���Ӵ�K���R���}3�z�aG���Փ!�k(�nҊ}�d[JjU�ܶ/D��ʓP����Y�6���Qk来[����ZM-.6�RKFIa���3F��,Y�T�U��C����Yz����.D Ӣ�>����K������.]�v�7���c��ިd��L7G]����^�1\�5�53r��s"!PF���4���-U�M^�a���6��y���"�wJ����M1i�-Vԩk/%�&D�~s4 ���֌��\��w��8�����
�ˉH����X�#)i�6�[�W��H""�����u�Bf�%���r=_I{	8hJz���/n��j(t�=�o&1��U�+G)F�����n��aZ��6ͫ�����;�`I�w�6�A��6�Pʌ��qF���O)�!�{�bZ�����x�R����q s/(�n���^૒e8�����J%�\T)�)��/"���y�M�Uz&їh����-��3pӀ�bԄ�˩����Xq�F�P1�F�ѫpҴ�hڶ��v1z�a�mS�»I��u�y����J�Tp�� b����X�X�Xw.��͌��{P^Һr�`�D�#L2V�N��h�u���f��Ɯ�IB���"X6�s2��X�9�̴�u�C�%�[����ӻ4u����w`�伣���$����b�&�7W�U��Bl����,��ǩۆ�Y�RϜ�ј�L�؊��E��ł���M�ܺcr	$j��í�Oq�Ԗr�0��f��5�E޻VV��
iS��7np�m��骷�7t�+kb	*��zE�wjKߓ��IF3A,'6f"kKb#��Q;����0�̫��mZ�%)viV휱�pkU�LM�22潋/u��}�)<�����*����,�{J�h��cv�RZ&L�ڲ��(�X E��fF�9Y��괁n�`���cJ�+5���.�w"Uv����,�-�d;Vt��f��/�v�V��N��^djLN�)�YJ���]�F�k�r��d�7�(2��j_f-�*�4t���4"�Wڊ��x2�ܵiZ(=��U5t��)]�*���KM`��k�n"��RbU��q� �O]���6�7r�3b�W&�Jq+H�:/�u�`.]EYZ�¿�IQZ�m���O�]��$%]�͵O�[{�\�Ш��ڤ�����l�(�$U�ÁP�:��K/fEĸ�H�hf'�,Az�ˠ��VT�S�Ph<�7(�+^`�t�In�,�!fQ�Cʛ��R�hQ��66��$�v�DG%ShԬ��Jk4�0�5#UdT�&�Ӷ[�$0����i��)�L�2��Ÿ4m��5c�v��hD[����-��ӁN�(���2�,-3�![��J�f֤hc�yv7�g;\����#�&2�)
a2���e���x�ǫǚjaQ�����"w``JƘ��T���N	2L�̐۩Щh�ɓ�	-���iMB�_���S�4
see&��T��׮+��ŵ�t���K P�XIǄi͕md�jSi�@2햒b����i9иe���X2�kc�GX�p�]b7�%MT@�7ZА�w�`	e��UG	VJ-]�\�2�ɔ�n����bʷL�Ŷ�c̷j<�
�P�E��� ��*xM,���mI����fY���j��4��R��nM��0�(��Q)����S�Oַeӭ�	z�%���),[��n�8����T���q"mu�@^���ԙ �M�W��&Q*:26�MD����4/V7H�zHN�ͬ��)�K���iU��7[t�����2eLR��oI[���&�A�ȷlD�AB�.+5=0:cI�z�N��G���T�^�K���,�r��U�Q���ւl���W�q֣����M�nX��.�A�RIe�4�#i0��v�*���԰�\֨�V tq�܉mf���Ea6xeYD݌�Xu��<Ō�u��(����q`���!e��|�H��Z��.Y$�r=���1�J;wK���@$ҁ�
��f��Km��d�����oq�t�d806ν�Ӡ�:l�k�klR ������&�D8.�yrAo]km
Dʘ.��d��$d��7i^<�w��;�T���K�c*���5����%T�\���O6[��-ڎ,d�1b��Y�%�#���L�j�B�㐭���Ɨ�X��u�Vԧ���B�)Bp	A�f�[!)mf�Ve����%��[jm�3w��
ƪ�!KW�X��$�u��o�2\��BI�}�����r��o��t�Z��ц��ۆR̲���Tc	��l���D<��|fG�P�qAV��e��V��Tu��--tif�cl�D 	�у�-$j@���VÃF+�Z��d��B�N堨�u��Z� Z���/ZD���	+��Ro����2e�n�!��_W7v�y��2c�B�5�=����d�eTV.� Om���	�bЂ.R���˒�ړ�s_��+U��fh!1u�^�S��P��PJNs�/��KIO0֌�R��Q;K.�#�E4MG�ǁ ���v�-Xd)V���v��p)����%V+n��9�1�kH+���*�)a��Zē4�r+	�i�bLv�h01�{R�Yˁ��>)�u'���l�	h��"�u���!�� �҃15{���U�O4���DawD\ͺ�n��!a�5p��i����MXa�������G�.&��5g3#�kZ�Y��:��M���i*�A�q��\���c�f���̋e75�^i�Mǻ3{���D�R�\�3Q`�-`Zi��C5K��'�Ct��8�#u���z�=���pã��X�l�6B�ҡb�yD��`0&J�`^c���6��O)T�v�!lU��D=8j��oP��Ǳ�y���@}b(d�:N��َ[�00rJ0Lwr�e���.��Q�kv��n�Z�`�4찴�
�������YP�ı��mn��\�?(�]��f�QɅŬ�751rZz%[X�h�,e�) �L`n��t�2����{�X؆��P���,`�Mt�夶�EeH/�2���R���r�NA�/3fZ����Qœh�m:�e+;A�5*	e�⽭�4�F���j����լ,0��2��]֫E��ެS6�:�&��2#s��n*�L]�RT��$���f��,��ol�i�FRuR��㷢�m��YiQ��`�C&�y�S�4�J.=�e]�SF��OŔ�T�A!P���X]�p*z��f=X�pz�ݑVd �Xn�jۡ�H�����g`����L���C��C�ֱ2�E��WK(.Kp �]֗Qռ3X��Z`��]Cjk���b��ɖ���{�4ۧʉ���bӢ gF��m�r�5i�(�vI��N��u6�̠�cg��&�nـ^�B���M����t����z%l��73J��QM�Y�I�qMw�(�Z�^�2'��8�3��U���Tnn-�h���6�Ke�yhޝ:��$��m��zvY��m�2�⤪�7J� ���������7���hВ��*+�63t*��������R
J���`Q�K�(R����uT+�ۛ�&n��_֥11>��*�^��k�}�4Y�a�v�{3�Ip�Z�S�"���jmզ����v��}5�(-t_i����|�AKy\�t:������	ǜ��(򕆻1�ׯ���D�zw'�T�o��� dn61�o^1˅��(Ovϟ ӷ�OkF��[��"�a˫-�*1��F��z�LL����{djQ���Zε�%��V�1q�S$J�Ԗ���(^��K@�F��w;/�V���)�q�Jv����K���4�v�8;v�n���U�'h���%X#����3%+,��7���0f�M�Ӭ��;ln�Cy�������*`.��)e7m�g7H��0\Ē���k�Ω�𹺵��� ���'�V��;VՁ�������ɝ�v����h'b��ϊ�A ;d���˒	��R���^����W^Q�k�/v���b(�a��Z��Z��\n,C��.���I���)��x/�%�޸�>z�'T�D�Gd��瘕e�Z(T�Í���Nd�XJ�S����wcHC�&o�vlARآ�>������c�KiN�u�\��Q�TJ�N��S�R��Ms�;�CUdu��[�C�<U�vs(�k���I�wz�9z����[���F����S�v4I
z cy]i�(e�����]��i:��aͷҝ�Ty�m�j�<�y�8ݐ��ږ�-t��m-1���î<�v���d��5y�&�
�z��|�6�Qc.���ehV_^V��|����Ҵ#�\����{̶Ky�ƍ�S_N�ޝ�ht�)vf�u=���*C/# ��f�L�B��N�����oX��4��e�>�4�hv��i����,�{��u��fR�)�sxkHS��}����vͰa�b>q�\��t��rEh`��>��\4�$Ţ]�?1�>wz�e�u��(QŴ�LcON�a�+�iJV-]��.t4;9ge�mZrbx{,e�t�N�Q-R�]-���6[��ɱ> �fw�*����79ڭ�M��_�`�j<;�p\����w�i
�^�Smڧ�N8p.f�����bwka7�|�c�M�b��ϫT�H�&�ݓX��ɺ ��xq�,g>; ,��QH��3+��w�=����*gu�Фk^�@�����C.�K��Jyغ���[��a���0ᩝ9���n�S�VkUaP�l���]�]�������<��f�u�o�t�C.�h���㳒�́"v� 0�E�F���ӏC��Y�16q!���*�\O��|�X��͵:����7�oEFJA�B֕�yx�e��:>TPE�h]+��m�l��L�]��Q=[k��$�e(w���"�q����
R��b�r��і�Ruj�kѹw��[��M��FR38Y���܇r�̧��@�����X]y�*+ptǦl�ͣ8�k��;z�q�V@�� oyTN-x�u�NR�v7���-�ieMOs�鶰�ZN��p�GX&!�A:ᝓ��s�P�N��ys���g����S�)���u�i)f���2:V�ZD�޶�AP+%v��nn����4�t6��(�ީ[�P�;b:M��[�����+HE����2��׀��2a���F�GP;�٭[�,\��CvjN�)��}X�T�3�XZ�ͣ}D�x��̻�s.���Y�[*^u�m
����X5��z1K��5����d���l%��J���A���M����v��Ư+/m`[+���.�5�P|�j�ç�����\R��`�z��[}W�/����Z@��f`�F��@�X%�ֺ�j�e�$�'e[g�^�;���e���v!h�80����&�#)�#N<Q4�X�-��n�c���p*�cr���]f��Lؼ��s0�у"xA�M�h��*��sT�
ٙ�U
Nn�0qǴӥoMn�c-5\�sC���f�H>�afu��D:��?f�5O�����Jօ�S����\�YZr?��j�Vi �� ����"��FX-f8�ND����K#M�#B 
�0�S�ɇ���j� C#��n�*��,m���t뼋@Р%uib-KL�j	���wq��o
�Av`N��&���k�a�)�es��ښ�q�t�oP+4�zޡxh�ΰ�]D�C�I��ė� y�띰+�˼c����<WbY��T���8�!Ij�6�k"�g�
�lP*U��7M���p}Y���*�X����[:j⚳P�,��RnR�4,��9>�A���*Y���U��y�.�ߏM�u2���m7�X���ՒC�P��ou.�t�}�l��Sbv��O�ՙZЮ7����{XOM3�2�upb�i���b�����@ �AsDپi��PI���,�����¼�=��ː%mdvd�h�\n��yZ��Ai����;�u����Q�8Oo�ذ1O��ɔF�q��@�&�P@�Y1Omɣ��7�6��0��G�[��)�ugS�i��0�[wQjd��)��.�K�Z�Ne���YgjAr���}�,�yi�y�5*�^@|�
��0Ӌ�i<R�;o%���O���Ư�)L�9Ք)�/3w ���ͥ��Ŀ��V f��*�%��q�z��eYg��ӻ]����R�v��m��֓y���0�wxqAaL�ڃµ�����|�	&��-�x�[�,s�LoW/���᫝Y�<v.
4��5췗��Y�c��'Q(�w��V3�S��,��+nc����I]夭�zy�r�Qe�{\�F��iC"#�4�s���V�\t�W)Տie��[�ݥ'n�j��þ9��x*9[Eo�E�i�΁����#���X1�s��]u�]ا>�	G���P�͵G����;+U�PrC6�ܴ�w`J��w�,���n-�kP�99���;e29^�\vp浬�}���v�T���T�0��SU����ޙ�%˹gP�-,���^.�3z�6�,�S�k��O�;11���mYj�b��6�}�鼉<��s��pT���lC9�W��zU�V.���w7Svm�6�R��]oT͠�W55۝cuŊ#t�!�Rn� �i��rv�!8�K�G�,�g�%+E1ҙ�r�3��=��7�+;�Y��؏�זs혝q��a�Yժ⍌����왙Тk5�V(`�xq���om֠���Cs`K;��Ժ�a�\�JǷ]�{�yV�Ϋ��]�_O��u���t�m�#�lMD&�X2���ws8����0��a���2�`oc����T���7n�[:�'}��șF�YK��mg��L�h��\�p�T�������K6	)w��Gr�Ӭ�/�iu�E��G/+֝BEKf�ٷ�ëF��
����}�f]&��ojj��m�p�n��Z�A�%I� nQ����wr�Gu Z�*V(q�C�o�%ɑ�m�/�����������y@m_6o��yӨ���|�TX��v�{��8�S�KiM���R�ڋ�6EP����[�ٸ7M\��Jr�n*�ژ��z�������I�R�^d�%����X�9�kMUc�p&�W5���cOw,����0-���Vd���uw����DM�'&_mB�қ�g
���� ���i�d����n}������蓳�b��՘�"�X��Yb��a��k"�Ӧ��i��q��Mܮ�S;X�ېh�W�\Ś�k%p�����̹�p+���\��&���FIf����Ԧh�mMNS����sA�A
�n��(cgd͹O��oq;��w�G���R;%�٘�[�E���f�; )�[V̎�-�G~�wtd����4�"���0;�"Xw�YP'10�m�m��m��m��m���p[�yZ�Td$�e7Oyyy4�:rf���h�1f�
B�n�WD�]ܺ�O���MI������Z��r�Mu�v���Do�)�_"A ݞ/$��Rmy�l�c���O����?� rҤ#�D?Y�,�o7l	�gq?�n-̪�bB6�%z��"�5��F�j�*�vVtH���ێ�Te�i�%(Խ���Qu�q1۳N�#��6y�;�bȒ�Gn1ҟn�|�vh���7i=TM�(�3X!5}�}:!F�r���]��t4��Ҝ��ߖS�`���6�����T�=Zqq�Ic;� ƌ8�����&�m72)�n��6�kЂs�@b����]��ht:�o��W[���pU�</��]�컝x��[1]^)q�<o�Qi�F�vl��Z���������Z%���Wi�Gx`2�>Al���;���X�MV`�{��^�QK5�W*q�)�;�z	@���$c��wp� �=X;�ҍ�ë���K��ga�~�Q7��&�8��<�_
Wzp�w�Gjo���b�Z+T�Y#2֐�F	��!L�F�Z�f����}r���)
ĳ9n�/#��o�;n|���@,Y�t�� �D n�#���n��f�Ҳ�H&�{�^�*ޜm�ٮ������X�]05�L��}U����`{זf;��K:�X��ܶȽj����_#�9���k5!�qK���r��d��Kh�_,���#1�����m^@732�M65�i�wkw��@DoUΫ��O;��ւ<]i�T�%���L�B;B��7-m��%n�E������~V���Iڗ�VTV�Z�_Jf�v��Oi��-b��y���=Qb��.-MІ�]Jj\b�����`���v�Wn�U)=�u{,Ki+~�CفGV"-��f
��H]��7�Pt�ʇ�X�L!�X�+�c��]a��#b]��nO�3�RU��++k�7��zr�JM���xв.�3hW3��P���mS<�8��YQ�<"�G$fl�{)Z�銙��Iq�$�fY֐�j��Sk�'Y�����3���UqІ'�Q
P��x�#"j.#�Z9I�<�	��w-Dvf��nr˽|��)D6'I��>/c���GJ�n�u��8|Uf��u�)DCI�-X'v�������\��7�G6�t/k�]*����W��u��K�?CK &e�mERne���ܻ��tJ�=)�o�/��]�U/����t�zv��Cs�^�V����˹�4�W3Ǡ�駶V��T�AAޗYQ�ʝ�s���v!��5q�4����\�ʸ7�f�}�w#���T��z�י��SNV
paгh�,���4o��@2���wBU8qU�\���׷pӭ``W��rf9�{onN�#G!�QJN�q����6ՀE�3obC�k���jb��`��sf��3p�/ �6_Aյ6:W�j�)��f=��]��[�����]wtO%,� 4f�,���׎�sZh��}���[/�n|�;Lk��D���1-X��}y*�r���S��ʭ�@��4`�;�^mMZu�S�͂�����9)E�D�higoj:3���3�s�iD��-d��`U(�l��34V,��>���ga���؟F�;�#~����2���{v�;�o5���L\�`�Ls�]��+7N
�)�I�,N�FcӘ�D����t�>,�o3�F��'{-�����قC@�X�q-�r��@w!�Bx2���fGܼ���b����{(��ֹv�K��|����[�ηrV����%t��F��L���CoxP �H&a�r㙶���-��NQ]�ֵ��ٶ�N�iK�y/����m.:��JG�"y��T��bK&��X�b��(fA�N*���rX[���
����"��FBe ����[����퀦S��N�m���./�6sx�9�-/�U�w�����t����v;i�+�� ݠu�H�G@�����X���:3Y[8�k�]<�й@/i^����U�w�n�A]��AC)<�^�b�}�����-�	V���������w�Qλ���2���k�Q�4�ltvwem&2�N��K���U�-�!�cޙ;uŗ9��I�9��kˋO���������]{�b�7��;���=��m�č!Jn��x(���(s��Hit��ijz�������,����.2��|_^+j�����
�:�����珂��ӝ�c=��MnZ2�O��y��������xP�f�����p6�pY�9��q�'ay�EI�i�(�ΰ鉼q��Qo�v�Qƭ��S{�:F���	���D�[i��
��e�u��ٽ+i��gV�{/H�S =��A��W;�a�
���p��6v�=z�AS�6�hH��y��VN�9�[����ʎs�΍�����]���Z%b8�tzq����j�I��)��$��:­g,ѹ|Q�%[Ļ��U{��t�2�:��bs�q[H+ߘ"6�i�,��L���f�pT�v
�jb�HT�a�9r�wÔ��"���
�.��u���oIT�J;�f��nA�h,�݈�0*��.	�'o�y�>j {t'��ؔ+Up��&bu��r9�1>X��L��pn��Y7z�e�q���Tچ��!/�4E���r]�E��`�`ٽ�-v�t�<Ϸ���T���)^��2Pr����ߖ�ҳ���zujO;N�R0�li���ݬɢW5 #s��6��Kڀ�ݷ�J߃ef�{H��q}���/]2�Xr�յ@�DR�왂�Ҟ�)J���BCu�C��p�*q�;�9�	TA�n������"{��]�z�I���")�/�]f���ik�t=Y�)��$��2���BF��eŉ��ʦf+N�g
rxNx6Rϳ���WVU��c�����;�cQ�6ν����o;��$ocn���M�ub�q��ad�<��i��6"�ܩ.��K����Og9z���*�>��7djS���
����Vtv�)���U�9j=w4A�q���ᠫ� �X�R����TWbe�@�[�G-��u6��&���n�_�C���mV.b먼=���*Vv�,I�PWqu�<�8��VQ�&^(rOY��G"[�܏bخl�u�5��Yl��=�tm�tf�P�����v�f�� ��y�,-��;�ם���r�q֔Vw뛗9<޺t~������U�i��}�� �*�7���cOu��hrŕ��5�|��q��a���j��9Cx	�wQ֫c�h��J�]-��d7��T{^�k��� �}����S�2��B���]�z��X�Ev�����[��HC��nV$�v.�ɬ*3���L!T�T�Rh]��G��HT4���EŔ�(dł�k�И%�JHh�v�C���D��o����Ǯ=�����J:$��,�qj7��P̧�_^�fB]�����+Q��ޗz,8]�듙![���o� ���G�v�D=ph���q+����s�bb�8�zR���1�T[8�^�TS�I�ZX�uDR[O��.M�ɧ�j�ٻ\KYqs+P�6B�݅�y{:��xt���0��y�ƞfV�ҝ5�%C����K7j�����l���9�/dX��x�a[�u�R��X�YSE����%�U5AEM�ߋ�����P�#�1,��#)�'+njxj��S�$dʾ�7#Iϭ`�4����"<����]F��79Mش@^��5��U��W|�v!Q�A�Mm�Y�n7Y12���V(�r��e*�^2�`2�a�A��UyJ�m��2�hE�8��u���ڜ"�9WN�ܧ���9]}Y7iȝ���@���
�_r;/��vԛ�wPm:Sz�����-'��h䖓Y*S�6
4x�7��6*<����1�R�z�yV=�	
j�3]fR��.tkD�&�l���$`^*; ��e�S����l[Y�G��_|>���)����m��ʿ�wM�???+�!"ɿ泝h����NyMC����Zhؚ*ʗ��Ќ�ӻ�t�r�ጬq�wVG�z֜��w��+��M/T���W����[y��]73x[QjB���Cڏ��_f��f�Ԑ"S�C�U�5���F���=��M�Bv���Ԣ�qs;��v�s�R��E�yLU����Id6:�\�-Ia��{h�Dh�J<]�,s�
�������A��������Y][n6C?�g��PsB��&b�駓	멡\!�=�P����f�҃@�E�H�{N�r.̘)V1Xv#є�iU���]� ���
Uy�gR��"@�2��Mڱ��Y˻i��*)ʧ\�d�ò�9�b�9�Yg��|'�������o҂޹����N���ڹY7����櫤Ntn~+�ލ���\��5s�x����^yܫ�宻����r�5r���e�X�.ƹ�sr�Z"|u�oY4sh�"�^0^�x��ch6-Ø(��rs�ʊ9r���3��.�_q�.�]/|�O.�j�.�'1ˇNQ	\�!i1�ԙ6#�WJ�܊M�qEE��ξ~f��o���s`ꝴ��wXQB-[.��u�.S�V$�wُ5ϫ��R_����D��H+*D��2P�!BVF���K�GB���z�o��G-&�Cb&�au�bԘІ�o,�$o<���]'�8'uT/�$f!�
"u��n@��w7O_`ȥԂ`BCC7�*pÇ6�8R _E2�d��n�f�����KZ����Y��wzn��n��$��D�<t���`lO!9P����n<����Lz���t�ݡ�-�Az*�<ح ?]���az]a��wV�&�yٛe��u
�ꤏ�T����:�+��~�#9�V,i۞uR[p+���<��2-iõVuh�S�K'_8�ޘ��,�6{U�/"���(��|�i`��5w�|�I�?ni��U�ʜv�r��t�qN���EWu!�B :�g�ܣ�:˵ύ�٫q�I�xP�`��/�/�aPF���24��a�$�=,���Xt��&5[XE��'Dm~���26c]��+G�;�!�E�i�о��F��N�M���ᖉ��DA�x�rjF�j����\qd�G�m�nWe��?n�����Y���҆��v劕����)��bz<e,jK8` �@_,TY�/o@p4�h�h+�w��+�d��'��Nw@`�H�R��DQa�����y�l���0�֙�k@��wA#�
�Y/�rU9�{����?A����|\���jp	�kIZZ�Z[�ق+��1V�������}��3��D� �Gng�����pwҬ܅e0�!B��ZT��!ִ�5
7 �����Ϫ����ݘ���w��֤�h^���MA�Ċ6"۹�T��[�Q��m>K(ŉb�I�z���ٶ;��k���R8�x=�#�l��d��0Ti����E��w�����|ք�$aC���!i�4��gh8�%�@�g{;.Ј��z�ڄ�@6���N(��b��'��eL�in��=��[A��y��������f������=�26W<��
Ԙ��ba�K�/�9hi��LV�"�yvZ����CN���9��+
��.��ʷ+U��\��
ң�#k����TYg���'O��q=v��X)���.�=�z#h��~�.$�!z�I�Y�L�����l�ճ�X(�!���I��խX��Zв�!��6�]����7a&��m�<�b��j��S$���iR��&�H��mb�f�Luv�@�x���&�Z�W���Xw�u^�j���۽����;"��<�gX�u�c�ήD���s�t:��@R�U��-?iT�M���g��S�W�n���0XR�}.H�L���L��Y�D�>��W�n�mk�y�ɔK
6j
�ǥ���Jف�t&Rx^ov����/��z���Q� ���;2��Ѭ���8���#�".F�ƒx��ƙ��li3S�rQ�|����t��L:<>u�4&q��a�P`J�mȣ�
}-��g�p�dD�3����$^-$�gNZ�����WHqNcy4�*t����PP#Jx�5��檺�/�Mo�R\���:b�2�X����@(���i��ʭ
kJT�#b������b�:gnZ����(΅L�������F����~�I���	���q�.�$�g*���wy[���1�
2��p(έ����&�z�3f,���.c�m6Ggf�B���������x+��Ό0#h�Tt� [*^�u]xh�di�آ+:�<м؃����!�Wo�e���KI:�����@�C�'�`�V�|�1N�BP�O���Y��o���fBO�����$Y���r�v�n�i����"I�8Qw#���P�f���*c�"p�wv��6��Og@��0�0�"hF�,�B�I6lJ�so�Cf�d�'�G�$�����dTl��ɮ{5���Pipi���a����R40,��Nkj"�#^U�f�_ڸ�kX��X�����Q����J�V�q6�^N#��dɁ�K��&6'���d��p�:[��	�v��ҡ��!}�� �oT�ch��.�<�z��C"W����lt�5�YJ9Ε	�����Ӄ��V�	�
m���l���i�$"���#I3���אMb�[�l������.�h)p&МW����Ι(��ְ�Mmk}�I��KV9Q�qdQ�kN�"�Π�\ы�W�w��T����ZBb��p�6��_h7�;��{����O��"���K��1�ڜB��NbB�8ZC��|Fg���/ �J�-$��V)a�">��q3T�#��/5Q.�*�f"Yđ���.k*=;R�b�Z�w!v�<����/#wzC�>z�T�I9�)1�a��	�;Un�3�P�Ŗ�4� ���@t1��w���Y���+�/w�7�	�����D���O`����<M���`L�{E�4��{j�B$)�Y�F�c������.N�h-׬�<�a�%:_,�[�Rr��w`�o�T-�m�V���ʱ^Ƽ%
Pp����hcH�_w}����f��8GMu	��o�n@��ҏ�g�+j$[.r���gN����r�;"-jCx�["���:����.>< �wdc�{�}�S��Nf�-Vx�4SL?�kJn4�9	ȵ�9�ݻ��O\kI<F�FN&P��d�i����.l:�1��\ؙ=���O!�
�ݐ� bc|l?-�A�ͿjW�����MNt��<+ƳL����So���ܼ0BoNU�u�g�0��"'\�(��o�f����N!�*�p��-��b���ƫ.��ķ������T.(B���
�MʽTC7��l�m�|V���g<3a˸G%}%�z�"\�TNV��Rd�j�>�G��gnfQ>i��i��c��4�ְT�lPf��Z�0�=E���w��������tһ�p��56f$�03kꊲ�	=�[�F��6~ľ�@��r�f.�/�\uۗ��
c'����Z�t��R�-�_����Ɯ�}�%��M9�͹�ӛ_WUq=�<�\�A��_:N k6~�C��&�ז�4�a:���a}�OC�Y���׷y��K�I8�=�r��r��1�c��lhn�VP���d��_2�>�z"��y��\L7je`�m'�o����B|,�n��\�ov�f��%�7J� ً������R{i�V>}q���w=�r�����jŋ��Ǐ��IR�(,�;Ң�3���;�]��]��q3���,Ŝ.��f��%�ݎ���	�n$S���~�+#��|��M@�{6��o�%��<W�k�3A��͆��qs,x����Q�ۑ�R�ʸ>��ڤ��]��r�9�6f�+	��3��Hp��A(��R��/o��3+�TeU�BNe�
��5�̋�\�u�+p������"Vև��k{����;L�x������kϖ����T)�rx��zwfpg�f%Ay��WC����9�ڵ��w��tT���_whr.l|槈W`Nl���)�b�����iԫ#CΏw)�/���'W[(4
=I)�����ԛ��%<	�,K��P'g�*���!ʙW�:��mf-Cqbq� F�IGԍo�Gpǁc2r�ԍʁ�K��U��6\V>Խ������ur��*y��h^����������ra���'j{+)�'�f�T��(}3�Ke8���8���μ桧�*���](���u����������ׁN��/�A�*���f���p��<y��:Zw0��dgA�S��CײB�9��/Vٗ������$7�/`�*�y|�a;2.{*T���g+)�-n�ێk��#�� "��+����w�`�5>ÒFle���$[�J�����%+̒�8�g=�k�q��AX�B�'s�6m�5w�ʣ���{;�$Ҫ�e�*�HjEY�K��Go�z�WN�3i��UtJ̙l�ûV�ު[>��g�%�.�Eh���VoE�P&g]ǽ Q�Y�{��P�9�U�d�M�h�33�i)�-PM�ǹf�L�8�y�p[�]���
U�e�H��ɀ$s��/,sJ�M�sEÝ�3�uvAB�W|/e\b��.:=6��5�P�}�s^��5��~��:�9&���*�օXũ �uo켏>Ʀ�6�i����f���6�S��f�t�_.ȵ�.�X]���]���73.��>��K�u�չ���_�<��tw1�ecp�*W�+��u,����m��l�	�Cd
���˻:�^��q���J4!�
�m�]\tf��H@��Df+��u��x���6�7����ͮ�eо��O�^N��L�w '5uu˲��h?N�w��t���YL�(�m�]�l)���f�;��z�F�V&L��*��{T�pۡ��r�u�2�t���q]�q��-�Y{ǻ+ۣ�uck�P7�pޅ-A�ԑ���r��`��;��,�F�v}��kq�v_26�����Z��;�'n �X���-���ƻ��!��}F��Ka��e΋��B��M��}�֡u���N��1�%�qy��n��xK�}��Ti�Mx��W����N;��1��Zd��4**�£�����Ӧ�ͭ��I�M�j9�lr%��Y���R*�E��j��9�}z���K歭��>J����@�y��2��AyJЗ�Y·]��H�֖l�ͻr�N�y�]ѸM�ok�'X�8��4�߀�¢� �ԉ�[���v��rDJ뺹����sr��Ӻ7:Q�h�q�Y���2�r��Y1s��̻���L"��JOy�HO:�mt$�Θ��.�w�]ݤ���;��������+����	��Iss9nZ�:��ӓ�������"�2o:�]�s�0\���뚎h�A�o;����w:�A&�+��ut�������g� t*�b��V-��ե��7�&/��/[{/ﾣ�4����NF�m�W�/:׍o;���Z��}��m}����_*�㶯�y����j�m~���������|,�>𹏀���@���G��o���ߍ]�j�_m�������2 'ﴁ����@�R�U�:�w�~k��
����Z�}w��o��/�[~5y�_�oƢ�?}U��_m���v4��#Z@���O�Gc>�.��V�}��j�o�uo��U���[�_Mo�מ}*����Qo�ο?<�^6�V7+|����<~���>���+���G�wv�kW�߶���E��}���k����Z�j�[���ϝW�m�����m�m����{||y����������j/[oڿ�Z�_�z�m\���������}��/������ <~���H��j}�=>����5�_��K_+y��j�j5������������^|�}*�6�^�j�|<G���#�����}����J�w�y[y����Y�">����LgYJ��b�����6�|�s�>�
�ij�mq[9�mņZ�ud�#��N�<�>���9�xz���P��"�"iŜ�xB́��g��,4k��Hn+��bJ��j���=%�{K_?��s�`��|�%n#���f�����&�_Lꛒ�W5�KF"\�[�NB���Y9�������)t���*n*��(<�7{�	>�l�,ۣ7��rz�a:$.Wn��{Y�{|����wV�'���=��}��������w"3D⤕�_cs9+�
����'pS��N�j�
����蜞n�{2>;�a���$����="��c5���cs��]tO�o�D���pŗ�mFt:_�9��ͻ"�t�bm�}��;��P����=���v/���x���H��g��ف�)W�}x���ɸ3k��sg^E��I��+*��h�tڻy*#un����R��U��.�b��]Bz�3}W��3�(��K���1��^���XWs�c(N��Gt;���~�V舘�������Qe����rkS�z�e�gyuJ��ݕ�R��30G�t���V=��JT�Y����T:�[�,3!]X�z�g����Q��IӛO{�Vml�q/s]U˳"�sʼ�3=2�K��t���+������̿{r��@�l�>�|����}KO���y�L;���'���z-�,�_��_K^�Y�R}����j�M�:����''��OS@��u�q�c����Z�y%3�jEwa�̔���Er��Z|{Z����Kȧ7�&ˎ�W���5���Gr{A�m�=��&F{�%�t�`���.���7r~�k�;������r� ��������{뫧��t�k5��{[��G��ωJ}����u=�3i������݇�ؾ��&��,�D5��Ud޼W�],�cxc��0�b�U��7_�����<nL{����p;�Z.����x�ؙ�b0\ܨ�Y��\�0��Y1n�;����Ǩf*��(T�,�;ݫ�5�8��*غ��ϵ�������]������0�d�n鵕8oh4끛�i����p�J��o��� �*\�RS0�Q��&�^[���&+��a�oV��n�F��O��,�t�EM���s;h�p޽�u7+���O
^珱8sKN�)�<+�K�^�L/޽}�MMQ��rx��sq�m-����|=C:f����S>�ȹ�.MH?7�{�Ч"V�[�V�c��RӦa5}����ͺր����kY�/c����؛�&u��ݯ^�����#� �@�Š�o���6{eθl<z��`����ٻ�7w:ENӚ+�d�p5�O�5��i�l��%�zw������7W[��oj{qs�A�\w��|8����$b�`m	��K���`���a`�qy+uέ�#/`�sk���/ލ�<K��1��]�r9�xft	u}{�y�:�xw~%���<���8��+�����U=�ϧb�w��*A=Cڶj�b�mB��Y��L�����1�Tf^�%])���8��� =ܼ�)�x�J/9�7�d��E��^�~�zcQ9\��=)^�6�u=Hܞ���c��7� ���?w�@k|Vi�s�;�w`��}g?Y���M����ݍqL͛�z�	�å��[�)1�hlǽ�jhW����j�z�:h���odwö��n9�Gӓ���s �<�PeP������[S��G��W���S�Ŋ�&��o�9Ռn��ts��7��oZ���ߪ*Y���փΑ�ۆq�j,=ͧ:��g�b֪�ԓ_��Q�?�;��̫n\08O���,�����)z�]eK	���=�����8�&x���3>u�_P�=��^��;Ϡ��Og�Zj��v�GƄ�Ӳ��+�]����e��L1]Ȭ���:%Ź�c�?W�B������1#<Z���sj����.�;���pd���~V���kcz�g\�h�y@Ʊ�S�sp��Hk�Ҏ��.���������@�z�*Ygmז�g�\)Ɨr��Tr�����/ S�ϔ��,t+jT)�5xYn�F�Y��	�T��g�^`��Zq�S2�'L�Ѐ��z�������,ʋ�>�3W���n��_�N;
o.^�`�6���ܤ���y�Zng��M��<) ٴ=�'zת5��W��{ؼц��6�?&����p�Y���诵���b����̫P���I��gOv�+��QC�Z���y�e={V�5v���A�c����r���w��&x��+=�pC��hG:bݞ�uٙ�F^S���X����$Ô�]��;��C��]��<\��*�dm��Z��l��ҋ=&/��e�u�q��U��E��h�~$'��	J����<���ft�&�a뻩	;qN�-
;s��zT�Ql����ż�]��:MA��w%�Yr&	z4�S�F�Y�����r/�=~��%UꏥoT�Ϗ'���}J��y�^n3�n��C1I�*a��<�a���o=��5�eyrXY`Wk�kҷÚ ���{B���cϱ�d�:�C������~�ދ�,�l�/G�״8r���S�'���m���W������7�~���繈v�*=F��w��U�.�{����Gg���s��^�]M�?+{@M��x��{������(���8������ozkB��5��Q�?eB+�:tוֹ� ����DN�p72� c~��a�<	��w3+�6�n�87���X�t��L�Ru��m1�W�y���ks���(a9�������u�X���| �������ֶzn���r���x�(��9��S�K��Q�\r��Jhva{�$E�_xՓI���N��G<rz�5_����9���n�._t�8�H�^T������}8/1�/')�� 	j�N�lI�P��g�'U>�|���SU�Ǯ�FYŜvN��c���:��)5]���+�#,k��ɞ��
�O9[��|_X�0`��sf����Vw��ț����\���ZJ�t�3�� *b�o�h>)�@<T�W�)F�3��y��MD�(F_�Q�����2����^o{|�u<qv�A�t��\�a�z8f��3p�5�LPi�S�k�^���T#���gEݬԥ�Q�&�\p�^����Wuu��*�y6%;F�ޕ����LgX�P&rd��]*H����Ԧ�̌"��h��Y|!���m�
�{Ӕ�����אo"&\�1����rNP��t��v��6ȣL�n��9�^B��x>ɒ1[Z�A�\�
5�nw7���Ŕ���c:��J��Nɴ��ƪ	׹W���� &��X��"WdN���9��:��I�e^���k^TmU��Z����^�:ܽ�*�3`��P�vS�J��'≴a+R���v;2��_`}Aܹf��;���F�'ָ�a֡3����\j=�^��![Vl��Q��^v�emh�u-!�w�T/R�*���L��6PX��N��TP������1}^,�fn�4�U��{ǡ���@�˱7,�}hʁ��P�khV8�W|�fvv@Ἑ΅_2"������*�çms��ԅ�{�6[nhB�э�����ٙ���C%.}�{�&��4o�U��O�u�I:^}�^���K3�����ى�
�`sA*6/��v�
NOlC����FrmS;��c=;"���ӽcPJ�v��7����GV7����^��Ґ������2�M ̮X�����hZ7�w��mL���3��=��c��+�]��NSz�x��_W2]�s��[�10���J8��p�˽��Y�f��J�v�1e���L�v��0۫4�p�8����2�	\b�t�'\ޤ�ď.Cw�ʑ�s/CG�wg������������"��8�.�����=n\ܛ��D��QE�L���7t����4�Ǎ�Қ�u��œI!�˼�� �z����9��"�P�M<��$̄�5�+�̅�P$d��L�&,�0k��#��$�κ�<ሼs{�dRW���D��ФP�A$�81��Ʉ�t$E� ��#�?���Ҫ��e����WsPN���=*��a�,�}҆9�ಲ'��W�}T2�q�p �kj6�c�P�V�+�����G�Bq$�����[��/w�x�V/H�����7��/���8��o*�z�U�y�rm.�{��P�5���_<�<��������sx����N'��w�7\
p�|�n��g1�y�{d@Flx��,���<#�9E�Q㽕*�W��#�1��V�L�7������+u�{�7u 2����w��lI��[·[�C��m-\ǽ=��}N��&���.�b.9��`[{�ws�����2XJжS�����6��N���n����#��̞h-�`3�t��Aӛ��v29��r�P[�p����m�TF����|�U�]�UǄLǽ��s]�l-��HP��5VZ���r�:�Sb�]�����RΔ�oO'y$�=�xOTqj��ux!�U��Nt�������h=��tX�;��;f�9+��(����8�4����)\�x���w_z���T��a���ޏ�R,)wA������k����b�FOf�n��o���jR�p�r�|�*�)��+�9�����Q�y�+t�p�'�k{�3m{���V>��}�e���6�R�>ř���eI���-vwY��t����� ���j��C���h��<���#��8ƳD��ԍ���l�G�@��Ζ�r�sf�#�����}�W�P���|qc��<����]XI�Yʄ����7p5����X���$\WΨ�D�g���˶��HT����ңN�7���-���W�{l���L�\x��[�|�ձԏ8�Q*�T�.z1t�?
�4Mm{Ƅ�<���n秌��۾//ɗ�O|�Ꞥ̃KU~�D�CGs:�j5���3���+��s���cqٕ�H�=���{�e!���~Sd��Hɖ�3:M�C��W�{�����Cg��x�ܮ����{��4�C3j���r̵��Z}���]�Q�f�}��ܶ���U��t�	���
=[���0�����&���u˪qy�����u׭���p�/��yS�t��*б�w13���W@��Ы�Ƶ{=�ź���w�P^a����� �1��w��{J��v�ս�"������¯�Sӆq|if���{	�}6�p�N~֡�q�ʇCZ���]�!�����*��Ú����o:�d�9���5��T�͙����so�	ڒ�N�+�qփ��9%�G������W��d��~��ΜR��~jJ�3 ���iȡ��)���O�t�<OS���Mm�v�;���x���y�l.�҅{93��-ΒP�{ܴvV.����|�k;i�����u,,�z���Q�s�_������������R��qE��.�~�2��*R�k,4�*��rO�d��v��r�����m��Q^��y�.#��W�w�R�f�m�M�퍓ϔ�삋ٿ���6�� Uk�{��6K����j�-Ъ��g����{ͣө��� �.ϑ��g�1F���vO>�_|��U��El���M�U�ƻj��%��N����>�ϳ^����B�q,>�޼]��2v�Ӹ��}�)�v��պKɯH+���?(U&ա�eq�tjM�f{%�#w��Ο�-���컿�����N8*ԕo�,�`��ON��j1��O	"�'Kz2��>��Ҽ9lt�z���P3s}����')�71����a�CWQ�f�O����7�������^��P�E<�g�sЛ��4�����b���)��S1��Ƽ���]�9�0cZ�#r����ݳY��twM��4�PS��V7�rk�+;7�}�P�/:�^v=i)��I���2��g�Z��Ed�H�kj�ؼ'�z�X����иsX�Ώ�
��I��K��{���	��&�/,�Ǥɹ�=a�~�Bh���\^71�si?wؼ����X�N�Ce4���'>(���seG6s<�V�j���,��u8y^V(z=���;��b	+�Gy��,��K�d�ƈY{���}��W�Js��?/Կ5xǧv*�sT��r���7_!����#���㏖O��x���J5m�WNy�w�
Ʃy��i;��"�{����ܡ�����'.z ��\!�w��6;q]���Kb>n���@����5lm�ܮ뭢�k��)
�D��zܼzb�<�U��g��|:�q�;6��e�I���e�we��s=�������m/?niP=��S�I�ؤ���x�zx�g*Vnmv�QteF_3��n�u'6ݘ�ootɊ��,����D�Y@d{"�xp�;��\��PN��d��Zck�-��h�n9�^E��l��;*� ���`)��Y_�z������eX���"m���i���"���
�����Ӌ(��@���9���~����:����<��ٮ��t62�&�Լ՜+�}����L�nhx�E�K}=��{}Z�l��b�����S� �w�ۓW=,��V�
��K��v�����y��Ywyo����c���}[���§N�V�lm�W-؊�'_�_��9k�6[֯wv��DM�Y�g���S��^�n9Jx2�qHK���j�p����NPO��]]�G��2*�M�n��m�ۅ�aΊŷ5��n94vK6���t����ͤ۟�����랼m��������W�`+!M��9O{t����r����}����sf�݉�$E�c,>tX������#�w�4�ʻke�oH3�������(E�.�j�^ܓ��}��e	��(:���]c��S��M�����t�y��2�]���ǒ��yL��y�E_�B3����R�C.��<d���д�����e9�hn9ٴ;��}�Q���AyV�ON{�����w���E؎�>cO�;�y�PX�{�����W3�B�ה�
��*��}��	��k���o�X���X�UZ3�J��i.&L��ym�����n2�G\�_Y:;�9� �=xv>�����m���j����+�<Lk�0x�>m.�痻��f���U��5�[fny��5�ȯĞ�1����|pzd�m�8\���l�e�WSzpyp�	����?M�X��^w�w�gzo13��������WP;6ddk��G��ا��o�i�܇h�7u.l�B>��;]�,���\��+�p�К,+��Gh�-o�Y�ȗ��IY�l���[��x��z~=qs6�+yw[+�=�*ڸW�~^+c^N�s(��ݾ2����[���=9��%^{|��$V��WA�JEn�0��ԃ�Oo;�����klM+�鮴��^;����&�­
�j�l���i���*�;=1<t�T0"5WT˽�q�è���4:S���W����®7k�sj�(�&]�V결��Y����"�4^���K�s�Ֆ���okI_a��S�x��ivv�J��Qr���Qط�t^�Cou���R���V����ЮWl)�{�n��4�_,������Q���C$:y��>S{8�|��Rݭݹ��WՓd"xjU!V���ᎊ�4��m1���)��ߦ�l��}��M��R�V0��2V�]:p�,Y�,�38����F`q<��}cl��`+�w٨�4U���b�Yy+�.56��bg-J��[��0n�Y3ҍ�4O!q*c|,�S�B�2*	�v"a\���k[��7vu��v��sh;1_A�B�tE�Ֆ�YU�5F�����HdX�TF��q���N7�,v7VL\.kt��l+�x/(���˺��'l�\RX�V�g�2����Q�y��;���bJG��3��{�n�]�:8�L;GU^%��mե|r�6�QO�d�Vm�L���!�甯��Y9�W�nT�"WA����[OeGi��&n�(��:�%�v�t��"(�[P�����#us_>�<7{���b�|qؾ�q��>�LhIub;�v�:w����P`n ���\���c�4��Qh#s�u�X�{�~�$�-��h۔q�\�L�xu�o����A��H �JQ�P����BK���tOZ�ID�������v�&�I#wrQa)0�w]��hC^.�.Wu���"�ỷ��ή����^���`�1$Ф�x�K��T�^uvy�u	r뎸�)�З;E#���#�:���u"L��/χ�ǟ������(�g�LR�l��P�y��������F��|q_�ﾪ���O��#[�Ҝ���צ�g�*Q�fg#�d�8��W�H�;�ڲ�}�RǕA�FTYI��ކ���j����4�BY�I93c��k�o��jJ{�VT#��ٝ��������{�3�O��B��c��^тۥ��}��Z�
oju��s039��9f7��yQ�N�}]��W����18�_OIc� �R�|-���|V�v�{�<�7!�Ȯ�װF�G=A�Qїu�WZ�+������6��Rx5�ڴ0�GخY;	�lg���W����{��ܶ�*�9B`8���W�RgJ\�0��X��e��6�UF��'"s�� (���
��=Jpb�1���١��-�q�M7��Fdi�57�8�-�t�>f3�����[OY��{Fh*��a��[j9?S��:z�O��4�+7&b��D1�G%{=Ƅ�Y�.Jj/��X�\��ٞ�l��=�W��й�x��Oy�i��}��$�}���5zb���_��l~��t]㐨]�Uj��=�j����'�+s��z��Ba�Ә�\p+�y���f��:W�+Ϩw�}�D���{[�����{���,o�.�Zh[�^oj0J�/�}��9�<S���k+#�D��}�(k���a<��/&�R��Ɖ���F�6���\`�UOX�w�N�՘f�"ě1~�����G���w��'�?n�=�8�o~�xkӚ�=���{yg�8�S�:t�����.����H�����s��hs�:�6�����S�7����Z���n{N��r������T.I�G����t9��:~]���=O����Ytu���n�^!\��U:��&�XA��p�tX�ɣ�8��`��q�j�ej��b����"��J�K���;���X��-��Tsq�m�XkG���Wv��)������\��6%ͰE�P��[.�U'�s�uZ64�=V��٢��5�_P�;��Jj46�,x�i��mS�3��ws�ܕ�����?���\�,;(k)T���`�ߎ"}^�S�p�L�|S򧨺�	g�Z���=<�����J*u���Q!':�z:Y�Let�In��wAcZr�ܼ[�����Y眻�x�9�������v,�'z'n� R��ޙ�n�s�vW;�������Ռ��-�٧����?�g�
�=זl����+;E��r�V!H����s �i���#� +�����2�t.�0���n�=��]ݢD�n髖�n7b�F�����xr��{+�Y����q���T���J�u!�f���737��+/��χ:ᤊ5}MlY@�{x�[�w3k�����G�]��At�T�Z�x� >�}[���[�������O҇WV(�Z��ܭ�^��~�{a�DKsö��y�]�Y諁A�\����0W��]Q`���p�=���׸Q���ߊ��s���&̮ӹ6�*��Q�Q�IV��'M��*yֱ�y�Mx�{A�x]j�^ru�n(��w�=��P5����������Bl֩���2�[q��#<���s��f���'�ƫ����Z��s����h՚>�/xb>�=N�ts]��.8=khʍ�����ɹ�0�G�UJ��sz{G�w��&�p���02p��ד���:����;3�L�N8�����2�oy���B�yt�]��gb��n+��u��;IO�:G�0��ב�� �B21e�Vo]�����;�hwԳ�t}B�)�~�I`ُ�!q[�`�+Scg^�4�V�T�;��(v��s����R�����J:��DZ��Y�A�7�쏎�
�>4���B��^�_ټ���n������l��� �h��2�:���n��`��ޕ�M'HE�{���ˍ��/9�IY�zZ�5��i,�[X46xh
�/9�͛𷵀�JX�XԌsU�=�L�Zx�ٕ���J�����q���Y8�l��/�(R�ѥ�6��a�|>|�݌�\�|�|}>���Q=п)u��/`���C��z�����<+W���Pޞ�>u����"u��>ɞsS�+�`���\9%���s٬cje{��x�l߁��Q�2�W9꾍���b��^�s�PSn��j�����c��G1�Z���y�8���+�}���8��'\�N��|�f;f�W<OR�=��{|��WPR�˨)��Z���nL־�̱���d[���y�3�s[�|��;�ϗw�Soi�7�:�U����ո�S�"8����� �q�,���sV�'|��w�G[�Ӭ-j����^I����|���ls����|;Xb�r���W��/u�?�<##x���ut���	����-�ˇ��f)^�(|�J9ƥF���X��ؕ;W/�t�3F&����ޘ�n��viB�Wi�-���˭[HZ]�u���9����;�l�s��c���w���KU��_:�����:]�e�o���`+|���vR,�/��U�{c�/9n!��Չ�o�w<X���]aL]e�Ws�����K�Ov�����>����=h�]�6����r�#����;�m�RD�[��]�M[���v.���.@��ܙ�Cv=!���|��Z�/���;��FU�/O�����Ĝ����)�rd��D{6���������S��!���Aф���`��%���eK��螐s�6��n���v����D���u���{�_hB��1�͉b3�E���{�3���S��VU�;�v�W<}�],��������s$���ysǧ����򥹹�:3��g��}狙�Ӯ���y���1���ڛ�芕.����l蟷3��A�Rƛ��X'c|���x�z�R�kŝ��V4�9��oDڷ�r��-�\�v��̕i[j٫��������y�wgwFYœ�;/�y���>86�M!f�Q����y�YS�Sf����|�U��].���%zZ����;�#�/1o?:nJ����m�,�<^Ss���<�n�<�.��r�n:���ܸ���,���1w�vlfiQ�P��_E�vL'����o!^�����n��-���v���OI[��!�xQ���28�_O��sR�L�<��g�nW�s�"[�]��0I5��c>��n*&}���3�[����Ew?K�*�>��[BX��a�L���͓/�!����2��Ԏ�#J&op	��H���Dk{U���R�3���Z�*���i<��|�3؆�C��$��h�Y���G,(%�(<��u/E���B*q��ֶ�;��We�X�J�{n
g^c��:y�E��h��˙v׮\R�g2�;����c���N�[�;�he��ՊV�����o!m������j���`bĥeuw���X}�׃5���$dt�%F�L3��Xk�C�4�pvm񭎅�0�4u*�&�H
t��%���}W�\z�4\T����4{��c/a���RV���E�&�hӾ�����隨�D�PK�e�tr���!{�̡y#��I�ވ�+�Ni��W;ױ\��- �n�\)��t�Y�]*���ΗHU�=�0�.M��dT�J��5e7wWf��ta|�B��2�*K�=��E�sw��Fd��i����BeAR&���1����J�č4����R�:�fP�@T�	�e�.j%��o1U�&\�Hl�J��vO�<���ǒ>�NH�'���Ys
�z��V�Y�¸���O�#Rk��=�J���W�]sATv���@�@Q}�oi)S���R�|��	'�`���]�p�V.�w�oE-�`���P�9�jP�+�Lu�C��������%�!���Ovh�n�lo@�̧��
K�d��f��e\���H����F��9ur�)����ጸ�k�)�E᥮��r<�}��G�X@5�����6F4����t����5�b�u��Y߁B�oZs^��i��$$G�:���v\W�:�}��bW(�1�eM�*�%�M�jM�t��A,��[8���;���g56�n�B��;��ʅb�:鷰l�(�q�\����"�(�<tA+�Q$ع�ۗ�\$�DGʸS��K޹$��%�q,Q;��h36	<[��B�r
(�.s�����-�ʮ�ݹr��|���"���&���AB�-�Ư.�A��������(��sm�scƹI���x;��f+.ฬ�%9��3��n�����ol�Ov�aG�}��Uq3w�����[�t]쌤�9B&ع���sٍ��g���=,orA�:�L;6��?fz{q�eA�V8*SSifՋ���i���{�V&�i�o�E�d�u2ܬ���1?`�:����6�x�t7��tC+y����/9�0��|��v�ED{>�0�1��sQ�)��U��w��'5V�>4^�M�����^�\f/R8��=쇛�1�|z��z�sS5�qA�����(���YY��5F2z�]��yŭeV��<F)��x���s�J�u�ػ�67�R������ց��2E��<gv��&4�Z3*�k ���ܖ+�Zټn�{SC��8s)vm�e��6v"�s|����Ybż>�ˁ:��d2s���Z���N�,^NH8��#�VC5�֫n�m�{�_v�\��U �gE��Wݳ˲�p��v3�@p<СwR�1q�:�E��CR�_?z�:������C<Ԗ��ޚ=<��#����"K�5�����x#�m@��tk��)�>�v���y׋ܤ|��8���}����_
u��f�����>~�۴�"b�V߳k�у<���}�r�^�}�y\��b�~}&�P��l��fmN)vvk�+b�^��Ī�d��Y��[m�!氹�)=�(<쾓�/-�\w�v(�E���ӻ^�}��}UI"ܞ����b �qS~s�6��D7ם��R�>1�6���e�q�I�E3
΄�Trt�>߱䠹}�=���M��u��qI�㋬�e׽1�tf�2��jo���xW�����5#���٦�rz_Es���ϼ�l8M��a�?�oo�%y��E�ٵ��ĺ00�q{�]܇8�ǒ�z2�}��"L��y}:k�yq���؍�pΐ���t�7����Ş�i�=y�جs�����_��K汝+3fSY����Cv�ڕ�rǺ}��{Z����1�~�e4��u�B�U�˺m�p��F5���y*=�c�m�u	����Y:owI��}-�֟��yC%��W�m,G����]Y����s*<��0�Y6��m_h�z�Rx�z�"��N=YO��P�M�Ő���Z��>P��+bE'F��?�`Une�!7p��I���8g�0�#2�]7����7���:RO����ћk�oM>N� ���{�t��4���c��:g�b{~�'�����˘�������PV`��"��=N��R��Vr����lV#y�2s�3׊î׸э��hC0�3\�d}X�^hj����v���л�T�!�CZE#nT�k�����\mS���6�,���i��k�U%�bt;�� Y���b���}�~���=��6�9ȇ���A�7��uV�FF߮y�L{~�x����x��oו�!�ze����Vm-Ur���7�L{Z�Or��R�֏uesgm�%�����{���f�)~�,J��id����������0��=�{+��O�#-�(�Nu�1�ίN�2��,���NF�{7��;�-9V;{<�V�M�HE�(��׉%�%�-��k�>>���ꌇ�6]v�[�'�[���w~-;��t7��������0�zh��u�K��1<Ls�bM	��;�jf�ʤ!���&j.A�e��p*udf�mI�k�Lx���-f뚘�ǩ�dlп�}_^$�N�~�E�-�p�8}n����x���^��~��sۑv3���Kr�m��:�D�@m��c��痨!,i�G��u���`��=3Z�.^ъ1QdC�+Ϣ��Ҧ��tڶ�k��:�NWOޕqᖄ?G�9�+��q���2OOV�}�R�^u��8���"����.����j��!4;�l�7t�V�
%F�,�*�	ޞ��Wp���2�m��H�$���W��a�)��{�0�.�ы9V�{��������]c�~�# ��8��M�R��^���|����8�=��Owe\/[XR�8bM�����fu�!�z"fo��U5\v7�P�l�Q�جtrR���\����y&��|������f�q�)�C7z��cc`]��nP&Ef���z�j��^�y�z��*r��f$���~`��u�W&�n��\Tߜ;�j7��}�*.j���8C�ʅ].���zb�٢5�豯w���<9c��oP�y9��F�v4�z��̀lt"�����ԩ��vi����b{�GkzmL�� ����X���9��������G�3�t١��:��#)}6v㼏�c�mfb������W�en��;+�=u{M�AۅV�
}�͜u��͹�M��rTνȸ���������C�M�/��Ϋ�,�o�f7�����;�d{4��)��r�y&�'�]Jt�����f�g�;�q����˞|�X2�k�d<��3s���瘼�������y~ڸ"�iE��n��~�~��I^��o�9���o8��jD���svê���FC1㽨� 5���Aޚ�����1�+y"�8�u�p�=+�-�d���y0Fl��$f��{ǧ��I��\?Q�B�;�{-Kq%HU�0�Z��^#-y��*�IFb��ͽ�˺�-���4��c�Ի'=��:îꮎ��j��R��(��F�vuB��Ic�q�ﾪI�9�c���C��j��C����[���t�~x��3�0�>�Gہ�Ϻ9ms��^L���&��+p{�S����7.����_�O1�~ٮf8�u��2b��������6�oN�]�μ��ćxڧ�ߏ˫B9�ngp���F^�|���;\�:�Z�W,�9�����f�k����ܳu nF�"�L�o�n�鮏��E�܋�s����f+���T���.��M!��5=&�WK�(r+�W3���e�����K:���YB�a7�'Wp�j���'ʉP�h^C�c�<wJ�9��NX��X%-�W��n�T�W諭������o��f�9�Q�좌���ʱ=�<5v�%�[��&X�������N��S˺ܯgi�W8lw��\Ì��^|WLChu�^k�*�>~=����eܚ��U�YM��V�T���n,���7�u���m#V"�Z}]�m��Oݐ��6f oYQz=j����u�	���W��+%y��Y��^�7�{��`��ݳ�`N+��=�3t��	�_w1x^��r�k�@�зN뵉���yG6q�Ϻ0���v,����{6a~&�?/�r@k�93f�p�4��rX�5��r^
hR"�&�����2H��.�V�u�pH���w+ksw�u?�m����f^S�E*0��y7��0�좭˥���:.�5t��m�fN��p��i�/s�۷��25���B��ڏQ�+p��9,��`�q�w[�_Z{�7M���[@��E�c�l��|�ܩ�D�.5w>����찎���I��g+����/ Y�I|���Y��{��Nn��\f����>wKz%�I@a�!3j�lkl+�%ൡl[�o]���4${�a��k/v�/�N3�bgCJ�d���]�z����ouGs����iq��ff����f�Qm��v:���:���;&�
e-3).ֻ���pV�/���e.��I�c閞3	cxv�����,��ۭ� �k�ۙ��֝�q��
[5;�c'-q�w��*�;Y}uѱ���Gw��k��*�KLҌ��Ԗ�f�=k�h�^n�t4*]��2I̧8/��0匴��T��**Y����*#���jڵ�1��.-�kb|Ebu�Fl�Y���"��1۴+��2y%�*��s�u�v7���e��n�wi�R@�mfu��_j�#)�cHB2vYx�r��#D�����Hƺ�����Z�8��jXZ��L���u���YT9M���pfMȄ���6:·lK�[�c.�,�,�R�:+@]V!d�:	I�v+�R�8�)�hj��3C�]��Ձ������d����23.��٫��U���� �u GĒ��S�r�F�9%��ɨ�-&�\�t�4QRU��yk�%(����c-͋.T^/Kx�E`�".���u�|����h2o[��c-wq��5����+���6�mn���<^,R5�Q�9r�
4X��I���[��k��[�u�\�\���k�y�0bўu� �� ��>��8�v�{#���8�|����׹žν���,�΃�@��h?��q��:�������\���G�(�@Ϟs��.k��ب`\����p]�vl_T�']����*s�A��q�:5��@����f���\�:�)N�s�z�b���\��T�
}e.͛�þ�ʍ���"P}�s�e�S��9�hsC��_g���3�~�E6(,��/�u���;C�O�Qs�9�ES)i�^�k�[���U���2��s�����|��ڤ�.��k�ᵞ�,'��·s�i�]=��z��D�W;������O8��ؾ�,c��r0�4{���f�6��"Fo���DROy��#�1j���V�}�.��vr�n~��'{{�_xQs�Ŕom���QP8��Qf��!����5�/,�lel��ȇ�[n[nr9��c1�H7n��1���GS4�g5��Dg�Z�{W���h��>��q��%2V�Qn͍����I�<�5����p�nm�g0���8;\V����MȪ.�ok��[R*w���k7�mW^���4fNO{p�q{B�o^��f��_����y{��L ЂY�I""k�K�%:��q��*�ǖ��U8�e�O@�y���C���un�q*�:�y*s�A�@[7�VB�N=@4��{��ڵI=�?Oۑ��T�O�|1�!G�*�?x��=޳���uo�)�Ӂ�����dI��@�<=3�AX�Dflyt��}	�����1���U�/M��/!VZ��a����oz>{7'��>�g�5z{;K�N9D?Q��fS3�B����Ւm�m��={�>\r��V�q�Af��cļ�b��t�(c<}�ֹ�nܳR#��o����L�̀:��P�o�&�ʼ��L1t���ם`G�S���@œ��{���-@^��2�7L�=��W��{�c��#��Q�N�ec�x�t�V���^F�L�q~�y9=GUŏ�ǹs ���r"sz,h�n1�_J\�,�z�h���3H��ےݙ`h���]�W�yR��W��;/���&�n��S�Q=ث���j��cz���_�F4`ڿo�f�Ԟ2��<�Q�(�O�ߩ�jƭM{=+=�UM�~zǽ�:W�>�Z[]~�<x��L�|�Z��{c���>�	ۢ��j����എ#�-���6{��p�z�c�^��������z%�J��Sy���o$T�ї/����"Β^8��w��V[�A�JW����{^>ɕn^�P��htS
�Tո���6��C��;կq��fR��.���v�O��M��.Q��W/ܭ�ϳ�G; ����4�{3'�W� �=�*�/mZ�p��'��b�P{Ӹ�n�K�JE�l�aV��7=W�{�O.5��mH��rҲ�1�S����ˁ�9?��m��vE���m�g4ϱ�Q�4��{�1�b�v)=1��}�<�;8�A�\w�iۇi��w4��}<u��h^R���C�Q�r�b+����,.����Ʊv���0�����[~ju=��
�SՔ�E�{�+%T5�Ά[��7��Rv�i;�L9��o�����\k�r�w.�_�1C�px��|fꦝ]�e��]��a�,Yh=�:�v����?�Ո�:�v)QKj�̭M\շ�񲧺�?t��W,�2��_��uT�=��w�
OP��6��� �pW�Ԗ�3�HQe���Z�Ϗ��k�}Gҵ3�>�y��w����X���/|�>���V{n�Sԇƥ�BF����UM�M�A%]oO�=���Қurc�M�o���}�Ԓ�c�;cs��7;o����Vw��R8�#�c5f�6��9�18�Y�1��T<rۧ��h�P빮Ȣ�V��*�*U�,d����X�*�P�A���8�gkr���l����S��&�O��w.��r�Z!��z�D���~�.j��O��k�ف:*�dM��yxb�^$��]_�R[I�n��4��u��{��W"�ҋ3|`�wzFY�w��y¹�sJ?e@��}}�v�0;i����Ōx��M��gfb}+:��Ck�V{�V�"�����'^��ό~0��c����
�|�#3gwv{��%{�'�0{�bj�>z�B��7� �s��VW��NQ�Q�Gێ��s"�!y��W�py͗�	��lE�%O*�� ����|Ӻ�wV���a�C`2�V�*�Fʛ����*z��t�(�.�q@�;�B`h��Z��Ե�x��J�CJ��{z�.�/��v!�U�
�������n(�"���㼋���%���_�_���^�N�(c9���s�<HIn��A�/��r�{P�O5W�7���,����6�ro�u�P�U�v�͙�ϫ:���݃o�]�s��nb�Zj����Ȫ|�}ѣ�w��1�F�<sb ��Ͻ�䵛���s|_wiz]��=�{�ĳ�ʉU��Z�C���J�ʬ��s����,�׷��?j��=y��ⸯgn�c<�U�����B��Җ�4|�=��t��B��Rdf�to�j��Ҹ����KhJv����Y\yeH�'�E�p6���.��k��U��ϸn/�պ�YS���	�73���t������{������-;�=��x���$����S� Q�Ϲ<qn9��ؐ��˚w�%�}�o$�v��d8[n��W�����n��*�9��;ط��&1�~�ne���<yAM��.�>��kK^}9�V9�:;LON���G{���ѥ����.�y;�7�	*)U]xR�s�֓�YQ�Yf����ʽ�����ӏ���k�G|a`�Z��)�z���ŲI
�)ZY<|���w�V����\�zZ�)����V9��:>-��r�6�Q4s.Z9ழ�ͻ�����{@�К3�`�qO_�N����o3I��{^���g}:s]ú��z�w��8�BZ�G�d�h^R�:�|���������
�z���5]�r�����
�{v���wmS�T_t��Q�O[����ݺ�U�A�>}n;C+vcIѥ��[M����~ƣ�Ζ�(.����&�.6}�oϵ�5��g�[@��Q�Y3w�އ���x��{f���א=(D�uj.O����]�{q�t1{>����t���XV{!�q��W����un�`���B����Q+5ч���f���W�-��f�`�˒cv�v����z�1�C��h�7��ܛW�RP�!�mX�ҷ����"�����^��ѷ29tA&s
���Y����v�� �v�ծ������W����΂b؈�8�\b��r[�r�p�Vf�[��ʉ�"���|�7XC#Y��N�'�w�ổ"Ͷ˽ؙI�γ�ZB�Zc67���u�&�".#��y�c�q/%��F���
���m^�v8�iW+���,=�xC��y|2�bf7ݺ�$�&�����1CO)i�Ý��%F�@�ԻeCu(m�k�bY��a�\���^��ٟ8_D٪�����;Պ�xu��P1˽μ����W�nu���V����ަ[�؝����Q,qO����Y��k�)�Tb;J����8]���3��X��Z_��Z��F#�'��Q՗aJw��C���E��mF��<�`��,�V�	��5�U��xZ��\c�Px��\�0��x�G���3Uu[���zxz���\z�s�3Q���J���6f΀�lmj�F�u=����$�̾��Ȝ���1@'wŮ��E�Y
�w.�f+�t�rŲ�p�d�t�&lٳ�`��l�k��Q��w��(@���0�k[�@5���j�'�T:�lr�*��f��"�\7yb�[�ê`������kWf���H�SU��p�3��#<�6����{Kwt����z�4����&=2�rS���ڱ������;k�s/��`�z�I�M�G���3I����@79Ӯ�)��ȑb<�_-(=)ἢݬ!ش�'1E_+��d�$����k�9d�u&��6p��ua��ɛ�c�����I��ւŹi�g騈໮Es�y݋I��%���TF���o^y�w^y�noyڹ]5��M�uʼr#b�ʮQ��Œ1�;��WB<V�T�.coZ�Uzޢ�����y�6�t�{Rx�[Ւ�T����"���u�K�d�-�oZ�;�Ir��[�]"��ߏ<ת筦�B���Z�<�n�癷jr���sF8�v��Ƿq���Ɂ�k{ ��y��u|g���%{���
�yT=��r(��0]B�rs�]d
q�C�t�gԕ���I�������G|������7�z�\�IYIo��:v|d�s��[�ߺq��Ҙb>��YCg'j2'��[=��g��t1o����\\N�aev)��X�y/w[����K��3;����q�_^���acC�{�lu�s��Ȍ��ׄ��2��z��Y�V_�m�0p����p㇧o'M�C~���h�]�(i\b�#٢hɉ+vmA9՜�u�bHxf�xs���}sF��N�:k�u8��E]� �������Zвy�S�U������I��,x��^�I��c[}vAcu�;�N9[o.
��b���d�#Խ���/�5}��f�9륔O�S����t��>�B��v�[1�S��n���G��k�b9�.:�n
�!`\��9*n����t��^q�l��1�J�jY/<��v��o���UC-��d��ٴ����}#{ O0�:@��n�V�Q�Lf��ף-�v���z8��X��7]��y�Zx9�����+�.̞��{����������MTEoN���O���v���+=v�&bfcX)O��j�k"�{�h�=9�e1�ڹ��'g)���٫��QfG���e��aa��}�𙓼'm���'=}"U^�����|�T5����ݵ59s��Y���)��i�X�|�1?{����_+�9p
s���9�B�(<s]}����<���$��~
yL]7�s�?{�eR���z��N,��L��bt���pή�f�^6}y<p|�s���Z�x?}'e���<��+S�v�ȘU*˽����=;z�
��^SW/ro��;"^���<�����}e��{�5�JN�^o�n��e��)y��7�W�3A)V�!�Jz�����0{k=����T0�u����̜���ۻ��z�����K"��-�l�п}�)ǹ�W�=�_E�hk��Y{�A�0&���'�d>	���ք7c���bI&���^w�9g�!S�|uӎQ{���	řӝ
��VI͖��O��
�`�}<;H�rN:���#�q֊e��	�b�#���:��߯�c�OCٹ��b��݇�������{{z�QJz�N�e�{��q���Q�R"Z��o)����a�ԡ�s�n�s{;���6.�𕞚JW�F?My��h-�sx�K�-;��[1n��	�.}3R۳��d��u��1C��Qc����V�Fw������Ɣڝ�94OmvؗM5�&g/�}����}U���Z���'�⚳g������w_OT�_�E�/辉�5��]9���.���'�^�����<t�1�^�b抝C���SΌ�u��/��S\h���xё����ֻ9<~����8�x`��.Ȼ�k�Q�Sxb��kO��<2��6��+�K�?M�C�t���^y�4Vi���x��ٮ�o�1=����*F]��#�P��eiO\7�s6�Kɫ�LX8��gbh�qr+$l�BO%���Z���0�f�Z��6ZY��3�-�N�.F�N�Sɨ�כr]wH{[-#X��s�:p�g��-8{dk9����S���7w����j�H����
beȡ&�9��G����l�����q�l^���N��Yٯ�<��f+j:a���obbF=��k[�{;����="Ӝ��D����Ӡ��P��������)c��t��S��ݨ&��zW�>�����؛7ؽx���z׺��/���ۉ��p�)w)z
��݅�]O³�h��e�	��Vw�.�ġ�T^��+݈��>LE���k�^�]�R�j/ B����~(c<z�qUܡ!��f;��Xb��{��t�4C���S�{��>��5sz똋n�W0W,��j���s8Vf ��ee*�)k�v��}_$��|8G<ݻ#}Whˡ9�I�N�벓wγ�=i�=�ouv��έk���=���.�j�:��rs-F�M�f6��6�R�|6�7*��n-\�V^	�LC+$�����p;�57�WY��K�VWW��vM��*�g����3B�$�r��r��E���C1t�I{���V?S}Kt��{e�ˠ���j�Hn���Һ��T=Cˏt�-�����I�7��sޑ^i��tǯٮq�W���҉%�R��LY���\����%f�);U�\#���랎�
��Y�#]5z�C{C!���4��%�5ǜM���}_}�w�����?Q��=�8S׫�Ɍsos����p������u�7��h8��j��}:�j�uB�}M�8��τ.�{�wV{k��j�hV�;���cl�vϨ�}S�x���N�f��1���§}qj�6 �������m���S/�r}Y�E�®�ND|s��S�lf��s�˝8������)V��U��駻:�U�$��.{�7^��������֡��+���7���?�
��������+����n+pyǳPܾ��2Iq2�ӴН��@�?p$�/����\k�Gٽv�	�"{-[v'���Nю��Nq��9+2�4�UVI՟��%�?~���E	�QQU��e�����f֓��Y'IkH,c�d�^��Q�C����U�\�G���\c\�9
����>�hS¦<�Fl��6}Aő}����ԝ��K����{x{68��*ӥ��gj"�����DU���Cb*2/�]G�4}�,�XY�& ��	����~Y~2��Q���gcG������㇍����B~���'`w�r�Y]Zߗ�_����-�MQ�X`^�2t���t�r������x�C�F���|��^ޯ���@}�^��,���ƹ����z'��V[�Qۈ�<i�:Z�]�
��,]ֿ�\��ж�W�r:'�[�5���S^Zǡ3��ش��Yަs�,WL�:R���gnhUΣ<c�$iu���}�x�����~�l���d��\�A,2t�*#��%�y��w���l�NJ���@��T$<t?F\��֨:�/��5�~ls>��I���N��<Y4� V7�&�j���ج��G���t��׍�������$a����6����^����zC"��^>�@q��.�>\u �B��f���;��^�ҳ�I�&M��Dw��8�n�*y@�w��z�o�GiHwڵ�HE\3�O���aǈ�\LǪc���?μ#�m�����JC%~�!�h����e!��'��6��25�4%i�Bu#���C����y\eO�sG��HF87���g��F�#NC�>�ZW��_�O�i�zmˠ���v�[�lfb�Zy�������.����²ۑ��qH@oO�w�m�uǩ� b����͉��y�qN��v��/vT�qɉ2�R��'�e�ݒՋW��_H���*^����,������G�U�(��Eb�o��V�W��
r�
3*�,�e��|j��`�PӠ�%�ׯ��km��w��Z�ZT�m4XHBT��A�v���g�{��W=׻Y�k4�e�!��O@O�o�v��`R/-h�1�W�� ����c0݆�*��TVŻ|�Т�Xt���X���v>�G�����s���׊�iO�U�U�t�$M��eq��fd���Orǆ���Eų�zed=7�1\N*J녭-��2����:�6J�+�r�[a;:c��O�
|e]Ӥ�+Oi���U�e�8��c(b�5,�[�O
�%���4�l�p�V��gpzU��8rp�sx�����QHx[x�'F `�Y�j�k#\�q��o*�8���,�,���cMe;�ge<����0������Kb��u��D���v�gu�!`���n�����T��/u��յ��h��j�8PC�%�a�ͺv�*E ��ĭF�E9qhͬ��/��!�=� ۦY)c��n⢦�����[�$ߝ�;uq�+�͗egd� 6�6�m�/dF��%;	�۬�X1�#V�ܭ�Ջ8	��)٣͏i2�Z#�tL�d���j��.���[�kyI���/8<&����B軶* ��n�����̡�g�S�)֓�9�����ʄd����r�b��kv^7d}�ď�� (�F�5��®U�W+��ەwvۚ�s[�;�5�׬\��x�淌kE�W����zض����TF�EE�6��Uwv��y�͹^#W6����h������x�^�����+��s_W��>:�lo׋^/Ƚo}�oRQox=V�cA�^wU�|�b׍m�7���BO�M�|���հfcqc����j2���)�&����a�IrQ�ٚQ��5�9�"R�VD���W�N�jF��6�@Xt�n���ۜy��}3�ba�8t�Dr�q�SPt�^#z��>�Wd<z️5��&� #ډ����s������lq�=���;/awzF�@�+uHHl}�@[������M�
,w���ߴC�E�z������x���~R�Q�fR�J��_=9[�r����9=��6a=`�
W�w���a��%��=r���2�	�z��F�y����V�����*}��	����dw#��r'wa0�o��h���\Q᪊��/����=��>���z�'���������Fڠ��z$��*����3�O���}$��̘9;b�ڝ��k��1�X���R�����w��m�ܛ�>W;s@xP���uՌ<�[�K/��%��^dҤ�+9���T̍}%�_�؂=ˍ��Y�1��2&���3�f�'{VOF^������$�v���G�2�7k�ӄ���F�dZ�xG{cgϨ��f����)�8�5#�hT-2f�A���*uU~��k�F� ^.>�����,ѝ^#5��ϟ��ʾd�kN$.U��Iq���l�fǲ4��˦��b3��S��O�Ta�T\�i2��I�R���b���wu9���b����=���|E�ȳ�&�D��g<���7>�|U`��~�
�<�`��1}�hu���L�(/��t��}.Y}��w�}�z���^�D�f3�"~��HH�%�Ỽ�Ws�=�^g�/>:lR�1��E�,ܸe�8W�G��h������A�����u� b��.��
:r[�#�u���h��8iMѕ����{�L'X�T�WJ�3�	�Zr�n���T73Z�����A�5i�N�:�AnE�Y����/2e���>�I>��"F��$!=����>CM[�*�ۇ/;Ƿv<!i�_6��m����8G�:xʠ�x�{Һ�~��[g�d�RR�$Y�f�d9��[#�g|���*����@����؅��qi���+䰶�]��xn�U�{7�Ã�I���A�s�Y&ε CL��j��u���d��ҙ�]^�,�z����y������{5.���*1�^;?8�'���8'�p*.4���VO�t�"'��v�큍Q�Q��4�ɛ���6� ���o���|+S/�����I����B֜�S��GI��HAG��]�
��^|r�/���J�ᯅY� M�*�1�/�ؼ�{
</v�U�4LjN�Er�W�:�r��h�kD�17(���P>�|t����I���胆s���[��kqM!�=�6Fl�,���ya��fN�<���.��fx�Hz:0����6ж��ޑF{�_�Jq���$�W�C�b%� vǋ�;&��<e��|��$\\�;��M��f9��g���yi��Ĭ;=D{�{7ϸs�3:�d��8��=h�㠅����$c��xL� �ձ��Kǥ�}�8�p(f��wC멁����E�U�Y�^W&{�;���H�0����P��2�]�gc<�\La�*(���B����Ć�C3��٭��#	xߔ�2E<�h�~�P�Y����>��PI�~�lMFZ�>��d]Xo(+"7f�
�ÞjZ���+�4w�\/�H :K��RDi8��T�u��%���+��k�5���뷬�ۉ d{���V���0ᠦ�\2Ԛ��n0�|C�ށ���ev�&ry+�-A�Yh���#W��&�E�������c��D���y��#�m	Ԏ~�sHy�M���ٽA���2+�S^,�;��4�dA�k�Tu_��tng��»��m�FR�,"����^�#S1�5�����`���O4ϒd��bU�4�v= W�He5|��yP�2�j6����8�#�¨&�@�XI�&d��&F�@�v��>�5g�	��#��@;����Bޑ����Ua���~�c��	����æ����!ҲH|��j�����=\��0è�����Ėh�d�=��1�����r=�j�ӯ�m�(ef���N��^�n7�:����]�b��1V{�u9Kh�v3�v�+��Wg�T�W>5:�sfR�ʬ�{��=�25a�K�|���2�,���'y,��k{ޙSy��a�\}�MB�3S7JN�6�=���ڝ^�K��i�>7�GƉ�*F@��ʌR����|zG�<�{��|�c��t����L���J���X�˛����a���N�"=�j� �J ^����*Զ�ȟn�Gq��$�t>'Pe�J��8Ii�̸��y��S�F�ǭ�Nj�{�z�B�'s,��l�z9�%G�� ��k���0�f�U�|��{���P��]���C=z����2���;�\A�ȯ\a����=��A��T{��Ό?�#�o��TүH�.0:��QY�@�D���te��N��[h��`�\Von��?�MBT�B�ō ;��:��ڪ�i���r����@�od���Gr+����}ˎ;��@�eU�>��&�*�2���ъ�t�e��g�^��/�$�9̂h��!{���j�{+���W�M@x��V�"�!���I���*^q]����ĉ4}��<o�ϧ�$�gK0֝�,���f˫C�d�7X�t��3��!fu[�z؆�Bo{<���I(�"G�**��@��R4ǁ�.:��:�dQ��/���N�u������<��#�ܫ���:�����f��'�'�8p�����>s&�>�����M�i��
>�ǌ�cʾ#�؁-,�a�����9��\����B�����i�`�L�������,�R�"�8T|�aW���� ��j�ҍ�H3\��Zye��*�Jn�IAd��8��6�V�����P#�N���byZ[��"�?���"9uz,����!r8��K%�=�������F�%g�Y'��4O��U�$��hx�g�٫�Ƀ8�{���B��K�̥^TF��DFL���6Ѝ���o��g�ɪ:o_9�H�>����ɾ�1�}��U��dr�Vg���,0EW�2�^�^����������#���"�0wˎ�7����N���GO-�|�V�7�8��w�
�Q��)	}�c�}^����8��&�Hd\A��#ظ��L�*r����y���!Y㟇�~���D�7����妒���4}:�����[7���ϻ�q��z�#�t �.E�Ȏ���푲�n��"y��#l�{3�1>��]*Ĕ�;�)���ޏ�}��̥��s�o��&���l�̓�ܓ���UM����B�5�-�2����cށɓR5��+���_yp|���jjL0�rg�����	TW��	v^:��J-T��d�:D��y8��l^l�S�]z��a��Q����I�*��&n�q��43�7|<4Nm������玫#���C�
`9�e�5���pɈw���WU�#��\�Y��qU� �l�A}�S��;�oyvU;��գ�M߾? �	���1Is��5�B���G�>Ӄinu[圴�<. L�H�����Ru�6h�:�u]潅�G���v�o�ȯz�z�L�!���v����a�ӥ3c��#_��f��~5�
_�1e�C<���c�eٌܒ^֒�ޟS��E�5��θ�;דu���ʞ��}�a.Ŵ=oS�:Y4��v���#XmU�\1w�2���f������®�X��D߬L�	1��������	rq��fz|<.�x��gZ^�HHl}��9x����ET�^�b;`3�g��:w�o\�l���:����TA�5y��KqOԆ����q�ˌ|��'^Ѝ}�^�#�����Lw�yue&Y�pN{�]���<�wm{|�I�PI��M^!�f�	��#g�Ⱦ]1Z���o�i�n�?F���~bUyV3����?k������F8^�>����#m(#'�^&a=>'��ϯ3�f��?L�z�̐�Ӈ�^��
��~P�gv���asq�����06,�#3'�8W�|9*!��&G	��S*T������K�L��kJ.��	�^�V�h!y�+$���L�oj��b�ģr1úo2muJe�Cz���D�%�e�Q�
Œ��}F*[ݢ)�(��Js�mw���P\�ls�_	W���Ư�m��+��Y/����[G^5��°��qYu9A�s��lw)����xL.�5���B�S�q���uJ(��[�`�mɉ�;l#�Ȼ��D5�:�5A,�2Tʘ�.�
�G\��[��+z<M˛���.��(�wj�Z�#�o"�5Ұ���)ձ^n��P�,�5l�TeC�Pj�b�k�(΋�ջ��c����k����m�0�a��X$F����*_u���XQ�6���ϲ)��g5�9����5�Kl�w�F� �&Z�(������������6�j�x}[W���1�[�R����I91`�5ȸU��v�R�u�q_�JS)1�Ue�|<�;^RYn�w��^�]&.�`[������:�4��q���js���	i%����մw�����}}BN���E�5=/.+/IF�f�V�����4���n��'�o�H^��~�M�2<��v�;��VM�L`���Cn,A$��m�bfȈ�H��/M��x)��2C�#��WRF�*������z�W�n���,h�i����h I���0>�aV�sb��b�8�8a\U lm��s�:}w��㝰�P�Q�:����p�h$�7��թ#h�U�-�d�r嬐4���f�ڈU�ʚ���q����]#]�ћ"����Ww:�Um���<�υl[�+ƍ�Thōz�+x��޶��k���b���]x�6����[�[����޵�Z幎c�U�s\�'9mxת���j��o�:��x���W�[�j+�<��\�9͊2nQxۚ�\��^���;���m��z�������p���Q{ݷ�\��W67��Ty;��B׍p�7�Q��
vU��۽���\�T��-�r)9x��p���h���{(ĺ��u�7O��nC�Q�ř�v��Nj��8� ����\Q�Rj=T����ڢN�.��+�q�8�@����!�ԢF��y�f�m�t��!������f~��6v�9i�4��I�S�Nf�k��Vc}r/��tٳ䰝�$R�)G�������4p��̴ώr���"��B~��s��S��t�u�.^�4�B� @����G���fA4|V^��dK�sy���wzD�֗Hn)�4g�����"v8�}��ݲ��yz��=&K	I�c��ӆK>�1t<��?jg1�#/��_�v! �H!���##�M|�0%is�,֠|*>���<�{����B�/��I��BC�dR��Z$�i��`jt��֥��/y�+����;Z8M
��ht-�����V0�]iۏ3��[�^�lbk��6�*��0'�323�aGfT�>݁�x߽@���u��4��9Pb3}y�>�ָ��E���'|P�y��R
����o�v��oj��������3�.Z<���ж����o������jL�gN��ў��\IA�ˈJ����훚�͓�xx�kM�P&��h��z,���#T��|���y�o��sP\3��(��D��"%ǌ�pM��E総��+f]��y{�� �z֬�hf):�֯��Q�r��lz�����gh�H��t����΁<���Ma�xW��t�9�l�ܻ�����T@�U�*~�4oV���Z�+��r:�^�,7�Ҽd� �(��/dGԙ�����|xq�~�H��\����
\��\wbx�LcN�wN���r�=�z�:H���n9�kq3�y���9�ɿH��Fm�޾wx3��Lt��;��W���:�ɬ;frn���<a\{-':����6E�ޡ��=��|OK�D$�+Hf�e,��=W#遫
��R�m߽��l��yH���Q��r�� �󏗓9�[���8(���<9�Մxz.F������j���M�DN�*�e�i���̔��Υǚ�N{��Eiyॸ69�f��<$�z2�/4&ԝm�������@��T����ي�{=◾4p�Y��6Ǌ�)*���<���⟝��3�fܱ|@�p��BX}>�1*��L���P�Hu}���Nk��8R4�g�L��#��p�1�8&���>����j��ә�ڭ��&�R�L�h����LZ�Rc����嗳آ�,bٟ���Fms`�Y�J��
K���]��Q�����i�����w����Å�8�Nn�M�_�~"쵟~}�p�,2_.!� ��2.j;���s����5�xB�جZ|q!7�3�N�9�,����p���4[^<v�Ec��� Rư�|��C�����V�u�p�w�"�Q�U1LLg��K�Hu�Ræ���[�^�[�y�,��y���RbA@_��p �������{��{��sz��	����Q�t8г��M�Ik}#͋��r�''0׻�����8՟0l��C�>��I#��1W��v��|��'�E!��f="=�g�pOGq������]�w�� �{�(��V�$�W���KZFu�9��2���׷����	Hm(	qm���L�(L6.����џW�/��O�+���A�V�"� pGygθ�F��D���w3C�v5wՁ�2�h�o3�����*��9���+w��oT3�ݧCj������w]��ˡ��ƍ}KOy��C���=�����(b�C��x�GmBA��F�t��R��[��h]�
8�>���= �hSXY�J`cY��_u�u53^n8s�I��^%i�m�z�Jݐ�f�i}x}�B�{��G���N˹I��E\u�kT�C��	�%���/��^كfO�v\Y���k�Ȟ���,���z�u�^ڀ��y	;��G�4��Q��2 ߫7uEk�9Z�z��!>������Ii0��I��}�O����^F����e³ܬ�Ɔ(��o�#L6�����:�_���|��Ha��.�������f��֝�yEZ��K��H�hW��a	��F��ab7T���F�qIa���C�;/�Ht�1;닢67UpřJ.o3O���������qQԜѼ�j�%${�}�W��>Ӟ	�,��A'�|����	����jy��}�亶�L+�ϲ!����l
�������QQ�󪶟�uRWϜo�vđ�JCѰH���hwr7蔏O���s/�`Y�q�!/oB<l{��y�&��2���9	8]���[GL��Xhς
�gނw��P8��$ad_�G�ɿo��Π\�H�**&�H�u%������H�6}y��7�^�,�<��NE5)�,�����$�G�A�*��aT���$f!�g�L��6�\�4g˯х�~�F��3��K�0��J�>���?@�-�)a��"\x�8&��E�uz�^�M���x^Q����TyRYɜ����P��K�������r�y�G]�\8�2\��Bۗ�����t}��6����د:�P+u��)Ǎ�(c�������6|k�Nyq�qdH����5��g3�{жb����Vy��|�A��5�-�x����a�Y��9S8�}\r����wu��f* g�>L��ZY���D;�Q��ヺ�ێ��}=Nj�Px�{�n��:q����5�w��L�di��PM��B64��2p����"=]�o�z=W�"�,��B�{�N�wV$66 �Y�H�=W1�����?xxW�'O���V�"��������=�m�m�o�����-;!Ői	n<y�۵�8�/�ԤO���>�}^�Q�������Hӆ,��u�9i�#�R�N{�(r�P�m�]M�{�<)�8�}��#hY�Z�q��	�Uj�n ����1S�c�u��t�K.�)�9���DV;t���yK��Ot��g"5�<��$���ے_��Zc/���)V��\V�)X���j����1��m�>���R:>�m�p��(ɢ/1��5��k��<�O4��G�yA��D��l�1���j(����ɹ~�;�}�d���.�����s�0h�HA�d퇈�;=�[�^�}2g�o#��6	��Z�%��5�L���JP�&H���[����$&�VGA	��ӊ��__g&�(j��Ј��/�����3~Y�WY�V������O::v���d����b4�Y�'������_�U�=;}�A����5��Q)�����	��2 �%���'�}]�y��׃��"v<j����H֫P@��JPkI
�T�{���?xW�И,fŘS��op+�4w��"��y�n=�,�eim��V�Իn�1�NoT샏Iٮg<��U���ؠODV�&���F<?|9Y�HveHӍY�G%ag=�3�H�X|ˢ/g��{���Pc�q�!&bP�p6Dt��E���q�\\�^BR�u)�!�ςt@B6,��I:�R��֑H�秢��q�e�}������v	_B�=�����Czf��7�z�I�O��cނ`4 (,���6(�����y�y�!c=#�^8�Lbdi�A��7�z�Wk�y;�;Y��Ƙ���<��v!yq'�DkA��*ʜ7���i����>>i`��L�H�L���h��߂�y�(��'m	0���C�%��M�i�A��s틩��y����B:`�*0��O�,����<g�p�(�F��������Q�};@p0Vz�[[���'��u.��8j
�V�]&[��y�9�?
a�C�f�|�����w<":;X1��q�L���R	t{�1J);��Gf�/ʭa�0���}SW[�;���"�>͆c��X���X��eg�x$���_p����|/c��L�X{�cmȽB��b���ӛ��^_"}+�M!��#u��h�/��WC3�y�lmK���r\|f��N<]!�������!��(�ִ^-]S��ov�N+9���S�L�H������q�5g���^
��'7��aG���H�7�#|�|YH!����lx�_%�N��W�WW��ϸz�9�y8���3�G$��a!��$F\�f��m����^���ˁ��i�K��8�>�2il�*:w*�ߓ��z�^�6�h��8�ȝ����L��G�o��ȟIF.�M����+����N��Ze��ꃨk�� ���AC0o7
w����S�8us���eh���9t�8�r�Ѫm�g�u:�������ȷ���lcG)�FҜh}&��Զ�H�\{K��y~O�7�+&��x8%�%l�_o��"��s�Y��c�w��;I��^���ѻ��Z�Y����\���Ԏ�����o��l� άEQ�%:�#*(tn�������u�n���M�h�7Ϯ�
�(�xxn�Ak:�;�5���.x2�_q���E��wDSߥ-g5���&�n�o)��G��vi���1�L6���8C��"	3Y2�O�Q�CJ�>�O�E3���&��Zk��Bv��yr���I(̣]���
��Jm��5�QңR�"����͖y�����������u�����3F	�p����P6դU8M����J����Ĕ7�u(uܱb���\w�s�0���o){��V>\н��K�"��%Pgz��@��$����Ƅ�J���e|���ӳ�y�BTe۸,G�^H���5w�ma%f ���t/%�j�<��C򱼪r�G�aB�)�+�4gU�A��`����1ܭ��w�O���������;iR�i%��7����K4J{!xi��A��1��l���B�,�"���[�Z�&v�Yݏi�H�$�e���%�&�sAT��+IB�՝����.ԗ+�"�*p����F-h# 㗕K6��CHh޾/z��*eX�}}@���wŘ�va�3t��M�ڗ� r�orF��P��8�Tzk&q�<�QF�b�{���>{�w6L�D����R�uC�V;���|��cz�<ڜ��+9��C�Ì��.)C��9b�5��o��� (�[�ܭ�t���o�j5gu=���^�[}=b�=W��r�\�k�s�*�r��|/^wG;�󻚍⫇�r񫜬h��m�r��6��z�=�U�9�N���x�b�j�m;�r-���W��[�4�Z�^1�h�m�U��\�G3��������[�y�[�ش���抹b��ns%r� �I�@ "�XΣ���;��V�z�e�N�
����
mh�7p�f�8��
��������5���3��f<���!K��-�%�.'��G�2g�$�f�
qH��̋A�=#ظ���{�߫��W��4��2i��Z���V&�A�z~V8\��o��_���<����e�0�~�Ph�K�.\x�򸵫v����&���L����I�\u�#g`a��5���U�uN�y�߸�M�}hl\A^�ָ��8r(�+"Z��e��//���������]t3�z��g)���'"2�Wo-��L�)��sVR��܆��8!����m����ZPс|m}BdF�'���Xoɓ�j}�|��4y�"�����:�N�	n�	��$�!�x��Fkv��ī��^C�>y�	Ozv?�Сxp �iu'G%�@��e�.�/3�)����t��|л�͊�Ս�M��)n�b��fv�CqfvU39Ẇ{a�3�|��yP��GC��h�~z��'%joy_�,�;#�dB�9�hv���8���G��j���e�d�#�ޑ>ZfJ�ǎRgR���9 {�=;�lz_C��y�5�D�z�ZБjLhCb�ɞ�'yw1�J�������R�kś0�����II���U� ��^�=j`^�8����k㶡,.~�&���f}~>䗎����e�Y'��92���Q�Ýa�0g�.�y��ܰ��i1�C%2o`8p	[��4-n/)g����b7f�d��k�'��L�Ȧ�~�!��Ɏ	��SF�	�д�@���a�ͤ%�H�����Z�Z;����G��#�@>̴7ءs� �tܮ�����X��OQ���r�E@��=�gJ�L��u�Ne����2��98l��5e;���{����_ύ��8]DVzC��6�5#�O��n�XE{3ޞ��=C��a�&��hhBbZk<`���_�j_��8{��_���Y���g-"�2&�8�	�D
���<Z�����c��Ó;�Fj
�g��!(G��C;kRӲ/���D����g���!�/>��R4�΋<lؕ��r��� OD�����$�˾j	k�/����j��q�̡��;�[��9z���Bcb��)�$�V9uMn����:���'����F�Ж�MB�;\	������Aѽ~߸:L�{�c�<oނG��I�2��l�QމOٸn�w��q�.9=�|}#��p4:@'#iz����bZ�#f��Y-9���\�2pվ~���p<[e�+ż8��gY�ٯ J��R�|Wo�NVr<�6�L�ƛ\�6a�owW����{bj��lB��O=�#Z�{kR�ܽ����p+�"�bL�m)��Lz}"F&N�Z��9��b}��v}~v��r���\p�B)܌��1�:�-q��	�Sˠ��H˷�Aa�QU��#�� X���1��Vo/�=�z=��=�ˑ^S:xj��F�'�T�TMu��Q+�w��?u�1�E�#�q�հ�Z�d�p�J�F�Z7�Fn��vn�|zl�B��,��ϓ0��dX�r.��U�W\���v���>�A2sU�Cǹ��[�8c�	��$��ά��q�;�p��^�G���@�S� ��[�G�]��}*��.��c��?@��qt��D��G�L�r�x'o>�s���/���<�?m��%KO���_3�ߠ��\���AssMկ4��eҏx�d̤���ZZӊ,����Ck��c!P����K����R*a�#Z�	g��㥥�z�|���n�h���+�R���wH��(��G�=Q)�w�U�pwj�(Lz��2OoF}����@�9�Y,ɪ��Ws5�sc��6��+��a~����'}*��r�N���S��"M��6dz�mz�*ֺ�؅�|�9�����{i��r5��(%������;���UzǢf~x����������<d�!�L��3p2�4g˯�0����^v����;�}���>��M��鼘���ߏR&��d���I�\D���-YNb�����n�	TUN�k�R�Ve*�Du$DxWH�����A��e�^��1��[L�͹�Q�u�2��eC,�z�*����nĨ:�i��eJi�^�F]-��yA�y"ݷ�N�����X��gkV�RV��W%}}��BS���^<��=��Hg�>�q���K+��t�ϩ����<r�qN���T�Px�������~��g��a��]ɝ9I�NW�TȍZM��'�t DZ{ݽ��=�lx�
�Р`�o�cH�N�$^��0�y��3:�ӫ���=���0=�<m�:\���t�)�z�d����^���̄���yQP��/���]#�A��[��^g9��"x�"Du�gL5��㖙���\I�Ǭ�=�'��N���ZI ��aR�B���4챴+e_6���xzg�Y9kЂ��Gj�tـ������%8[۝uo�F6'<O��NZgވ9
��dm�p������-D>0jA��b�v��\-|3��{r�a-õ��#3���A��5SN�����OeaB3��=�v�z���wΓ�jV*�1;��<:�ˡ�C�����v��ڈǷ����m9�xa�)>�V��ɷ�$eC&~�	��!��'��D������^HA���V̙�ނoՓ��Nj�*.~�q<^�sꛜ���a1hM$x烁��\YĄ�@�\X�na�t���k|��J��Q�qf���L����Pg��ȣ��{���ֻ�O�q�Bhk�r��V|��<��ң��=�˗;��	؁|1�Eo)�&�"k"	�M� V�ѫ)ӷ~��y��?Rӳ��#6��7�*�F��@;�s:={~���i���������Hn`�s�pك���@l��yO��cɕ�A�-A��fR�TC7ꁳ"=�g��!�x�ꞹ��u�alP�'*,�17��vn������q�z��f���n�߷ճ{ �IT�qm>�v�S�S&grjw�^�8K<��#쬫K2�7O���Tq��!�����lY�Y�N�Ԅ;H��1���<F4�r' {� �RH�>��	�d=L͈�::A�Wy�vW�G���.0=�&�������6'2]GG��z}�k9~�B�����	���T�����v��"��X�P<{ˍ��^\I�qkC/T����t�-&P�,"�bK:ҥ���רQd��	��=j;������⌃�^8eT	�r2��:�k��L�<��`�;/7��m�"���^�!a�"�	Y�V`��k����#n&߷C�.A�l��:�P���hU�Qԃ���Ϳ��'�7��糗��zr ���:�����>�����%���L")w��j���Y����n�P��7�u�YW	D�ñq;������x5U�_'�)��{�;pv�y��`n�gV�e�O����I���#�3~Lè��Ƚ�#<=W�����Y�Az��D�2�4%g)�8Ǻ�l���j�
8���Wk��kuќV{��bR��a{ ף���>��H�:�]��n(��yqd��i3��	>>,�t���=�Q��!d2p�ykSSˈ־�A��
6<Y�r���>S]�t�׶,�U�$-��Py#��$��a!�ɚ�;=Q���*=�>(L8�&I��p���}����w��C[s���v��, ���>�'|P�o֩����"���Cث\��o_���#�?1�}������� `�+�,;(YIa�RT)��
!���'	-�:�W�y��V.y\9����n7% 7 [Y{��Ӻ�H���{����_���qѡy�yVm�"
��L�w)�Rr+	S�c'�}p8�h�!����C�j�M�����,l�k��c�fδ=�|�z���G�}���l�p;˘q���?~<���i�8&�@���L}���''��qdL�6v�{om�s-!^]L�Z����2+�Bqqmz�^��ܞ���{#��ť��_8���h_��<���z��}��lv�>���&���L�E	Zc���Vj����@ˑ�t���íq�&�G��p̖p¸&� -ZO!�N�!ی^E�w�G�׶<a�,���0}�[�2t��n�F�D���|ɧ���Z��>���Ck�x�mJZY�7�h1��P����}�s���EGw�Hl�lR��Kk�z���]�|^��|�T�e�� ��kT�����mZ���%�d��6�Y�R�3o�^����[�Vv�p���f[*!�I"��iW�^x������_���z���kmm��+mm��m��|����_ۨܩ|7�Ct�,�l��\jKԉ��IU��T��
�Xߗ���M���y���Z���t�K�"��cL���9�ѫ5�ݡY��UmI��Yu�nɉ���M���?��~�6��v�+�H�5tH$<�BO�5B" ���Iw���u��vX�?���>}�,�����/�W�sy�%Y��I�G�O�߭�εJq%���LwP�x%��������>��z"��,���r(�o*O_)�F������f��*�����rHD���-w�����jd-D�Q�mm��k[W󕭭��O��}�.�6�j�Z��ؚ�6$ߴ����$�A�̙ҩ-�f�uϣ�����-�JW��֘8��cl���le�O7�,����ʴ�j���ԩh�<K-*��}��Y?�u��ٲY���ϕ�lE�cRN�y��3��N�V�0O�u8i����������N/�TQZt��B�}_&�&�4]T�R����T�ޑ" �W<	!}�
h�_J�­*�#��ZO�fܤ���1I70>c7�" ���yJ�������S�4�"H�,T�Xbj(�n�q�����6IL�j�K%jl��3�g�QzKY5��-�W?{$"r�G��a��D�AY>n�>�AN3Ä��'���'�ml��?)����9It�ǽ�7eb�'��]\���mu�;j��=D��E�.m�Te���HD�)�\��B��%�������H�9��`ϼ�%�����krm}���؜$�9I.�==�$̈́�(�"��,z�X���wY㾆>#���0�Ě�{�ߝW���4��װ˒����H��3��:fc�_�D��ۻ&q����)���Ȝ6��,�u��s�=DX�&��'IP" �IH{.�9I�$�+�z=�f���Ap��b�3&�q��hfc�-j������1��)��X�����j��.�p�!���