BZh91AY&SYV6,T��_�`pg���gߠ����    bD^�           ���"�Wئm����d 6iJ��i��!�ZM�$�ѭ�ƴҬ�d�I�*���U��+X٣��e�m�����ʉ���ƉlĀ��e��֤h+�5M��H&�l4���fUUTVٙ��4b�V���[j��`�
{</5e�w����5�V�����u�\WNZ�.��"�4�ox���j�4������#ce�c�gR	KԦ�x��%*�m��u�j�JՔ���ŉj���Km�R�i   ����2s�M��q�>�P���v���vًm4���s�C�׵ uK��]	��ڽMh�{�tM��cIS�lݚ�1�u��6�f�Vئ����mw� ,��2���h��z���9������þ�)D�����}�[jzҬ��O_cc5!�_=��T�ٗ۾�>P�	U��k��Ҿ���_>[��UvϬ�}�>}zeUR�{���Ki��c2(�+"�kl�|  3��R��!}���>�����-�e|�}g�m��K��w�N��4�%_z��Ͼ���l��oOJ�)*�ު���}���f�ޛ��m'�u������jW��U�����QK�ｆ�޼�[e&�,�mQVe��  r�ԩIw۵9󾾯���T�Ѿf��>��T�{�ܤ{z�-U�+�ҥ�kJoos���Wv��)�y���z��헧=w��	Kct���:�(+�z��[X�2����ʵ�Z͛U�٠kC� �ϯ�;���x�R$(�/z�Se]��mל�����{�M��_{5���ל��{�˕�m�g}}���KjZM�v���L����Vf�ն]������ho��j��kE*��6j|  6�u�6ʯ�w|y�v֚���5�iYKf֝��T��O[{�Ǟ�kZ[)oS��k�wN�Gw�����s�������s�z��{Ւ��ݞ�*N�M{��ש��M�Z6�6����&�|  v�}%^��{�� u��ywA�[9Ӝ��������B��k�|�(#���Z�ע��;�{��p��F�;��z�@z�BL�F�T)Ce�� >����p�^��9�n�@(�v���mU�Sl޽����^����x;��7S���+F��]h޼����teTQA��� ���|޷�� �u{ ����-jwI����ۀ+�7�{���뻓��@����M�â��mǔD�f�6����I�|  8��Sճ:����^ԝ� ����� �{�ƀ�w�����=�(�y���{t�N׭����  @     j`�R���&  CF�"��F)J���`�M���a2���d%*��    4�j��@��*20 �@�  i�	�JJzmH  �� 
P�ҔH)�i��Lђ=&C@2dѣ#�?w�B��V �Կ�_��2�t�Q���sun�*�߄|7��3�~���]{��
������_����W����������o��O��������?�h��h@U���UW��TP���^��?��?��?�"�[(�S
��?��O�`]`]e``a`]d]eMae5�5�u�5�u�a�U����A��5�Me��YYGXY@� u�YYYGGYXWXXX ��Q�WX	�u�u�`XP��E�A�]`	�u�u�`CYGYGYGXWYCXf 5�e@�T5�ad`]edCX�Me]`daea_YWYYSYGYGYGXC����+�"� �"�*k"� � ����,�k*�(���
k �:�:���l�� k��/�#�����+�#������*k"��"�"��k(����/�)�#��"k"��
� � �(��:�:�2.���������Q�����XX �Q�d@� 5�u�u�5�u����1�u�u�u�5�u�u�u�aXYXX�YYYWY�u�u�u�u�u�e>2��#��� � �(�
k
�(�+�5�5�z`aa]a]dY�E�YGXSXGXYY�E�_������*k�����+���:º�=�.����������������0.�)��#����)� k"�"L��.��&�������.�	�����0������������E��T�U�Q�WYD�a���A��E��Q5�d`_XGYSXS5�u�MdCY �A�D��u�u��GY@�Au�u�u�u�}`]d�@� d �aXS�Q�Pu�aN� �D�P���D��T�D� &u�5�u�5�u�u�u�u�CY�Q�Q�Q� 5�u�aZ`]dead]e]dCYA�Q�A�A�A��@�� 5�u�{deaMe]`]aSY>0.����L����#�	����k
�
k!���:�:Ț��º�:�:�:�º��	��k �&���\A�T�u�dSYT�A�D5�oY�� 5�M`GXY�@�a@�u��5���u�`�5�q�c�5�`�5�`�c�\q�gX�u�X�u�cY�u�d�gY�5��cY�u�gY�5�gZcX5�X�u�cX�u�c�5�cY�5��u�Y�u�c[�k:�Lk:Ƴ�kƱ��Ʊ�k:Ƴ�hƳ�kưk��k��NƳ�k:��5�cX5�o5�cY�d�5�{p�u��g�u�cY�o�5�c�5�`�5�cX��α�:����t�ì�Ʊ�gX�{q�]e�d�_��2k:��Ƴ���k>��k:�N���k��u�cX鵝`�5�g�:α��ݰk:��k3��:Ʊ�k:ζ��:ìɬ����k3�k&��kγ���i��x��<c�<a�&�k&�k.�k��z���������͌Y�b�?��M���R����yΧ�;���-�3x�nJS5<;4d{�C/vZ���	�t�h; ��m����?10�噻��nRˡw�rH�R�o#�D��s,�f�+EP���H�h����$�[0f�4`Q��n ]=uc��tZ�f	/\���b�/$��0�+l���6`'[+l��n�-�.�J�O6��h�nYx(���RE�pܓaӚX����R�RW�KzHܙ�ս�(<�ӆ���[?+�1���VYT'Fc�ISw%��l��"�q�Ն��(ٙ�,E�@`goj-Y{Cm�὇i8�_d��eۀbv�`#j�Ѳ�!�XwkB�r��n������p�U��Ga�rl��4$�"�+%�� �z�m��N���ݛ9����oH�f9��{*5j��I1jd*Kh�3��1@�B��Q�*�8*�N]�,�ʁjf�do6��v�Z�Y�4[�m���^2\�����m��
��m
Q�4�G�GZW(�~bh���nI1��� ���b�J��v��w���ČF�2�#l�f�f�sk/@q���`H������O$�ya_�Mw1�v�4lC��X��]c�Km�Ҙ�w,:�&��m���+w���S�%�tJd�� �z�$d0�'RW�*W��K1�u�T�� �Zěh�w%�Y-\�sq�{�\[Z-��;Q,T�vM�nM-k3dm��$�V�Y�t�M	']V�--T�b���3G�cw{�+�T�6>�60~tk[��Z��xhc��b/E�y�y�wV����.�����y�JA+5�8-uv���ϐ ��KJ��Mm����ul�N�7˕�VSj� ���<%u:��z���ۻЮEK{`����%��b����;�I�V`A�d�"�EŰ-��щD�fH�a�Y���+F��䳵�OQ[��&K�E�Z̘�-��&�UD4.L�,,t/m�7!z�(�9P�fA�j���`���đ�+ep����G#	�`�5dB��+	a�d���h��Yqb�k%d��h;�e ���UEc����Be�v�4�d�j�n���n�h��V�؆��'qϓx����r���b4��fĶ}���k�vтn͸��u�ˤ��#,j�#��ʙ��X���i��a�xoAhض�`)Zf�ķP�Zs��E�<�>'y�l��*�I�#��Z^3�b���w���$�'4A��ʼ�A^�F�d� @m�/0�U@˄��cRn�EД�8X���d�Qj������=���;"�$M�@��g�
�v)�\��Z����d@�DI��U�����V�M�˧.l.�
T�Gf-(��jt�ytѹX��-c�(M�tӫ�j,Y.~*S�;���"�1V�e����X�D��]��fA�*�At�7SD��l��ifp�j�S�V��ݭ�,��]��̮6N��2-���B�m������GvN���uX�؄�T!����eX�:��,�T�Γ*ٚ�݅/)���j�nZ�(�t��n�֌stݔ4����Bh� ȉ�R{Z;�wi@����\��wq�{)��:r�k�JYwD ��{6��u�~�I����6�ֱ9F�mS.������eFɬ�ce
F�s\#Q"��vX���Ŋ+�U�
,�zkY��:�r����C'����Z�i�u8A�1/��W4(7Dbw�`xAa���zkZMḰ%���65�)Y����u���64,���R���3i۩o5fPĬ2��4�ݻ�P��M�ǖ���ߴ�p� �ա�I�m�Ya��r��@<�v7nTY*+�!��,(��ڹ7%��t�YA9Z��E0�E���-���r]YKDj�hݽ�l�[R��vy�VI�P���3D����K��Ҥ�h�6�T�ɓl�*�)���ڶ���U�d����e�ף*J�`��ȕT	��'u�d�ꤒՑ�1�I,����'�� ��ӵ�����\.�5U�K"SX�n\�QJ'*~n�JgJ�H�(��I��j�(�b]�&��%ʺ�ݘջkS��R	,G��Ajk�[�p������(��4DҢ�Y�Ԋ��[���,L�I���42Pm���f���k���X	hSnkOM;Û�������{�BB��=��KF;W��`�1+�ClI<j�5�9R=��b��r�{)YR�injy"�sS95���o+�5��d�Z&}i��q��+t���"
�zs2��Y���9�l+*^�xjՆ�4s^������Ֆ^�6�Z)R���7�S�Q,*nm�C&ӛWK l{�+i'r0��"ۥ��[�de���9�ICL�Z�d�,\�@-Q��̿�E�kF�)�/a��*����A\ӡû�M�ƃo�bK�u��g5ٹ��l��g4<D=���Y�%g2����j�l!�Vj�`˫��ص3K̪-#�.U�l�ȵ��v�-U�5�ii��1gZ�E�6�Q�x�p޷m���u�*ݖ�R����/�����u��nM�e�:S�l츶nɏE�^&8q�v�heT�(�T���1,��u��ǁ�-u0"�-���6������6�S��g5���|q�u�Ҳ�U-��b�a�%F/�U&c�����y9��t�˥KAl��s�CH�|G(�{\��]�����y�����qe5���uy��U̔VCf�su:��H5	}�^c"��v-��]��ʔ�j�o�2F�R!�)Ƕ#4�|w2����ChɌRw�Xں6��2鋅�v����]�͏f]�4�`v�h�10��^�ة�Wx���#��ɻ ��q7�<5 �͗���C�P���N�B�V���7X�)�FJ�����Ջ_Xnd�y;���w�������QZ'wV�5z
�Co-CJ2�i�ߢ�L��v���R�sb��w��I(&�BDfd�p=`��Lsa�$,�%�\k-q�x�ڻR�n�͛�㫹�6����mJ�v��(����J����c���K׎����e~w�J5�|mS���W-����͙��k,mnjx�ID-N��i��)�:]歩l���@;eʺ�,�����R�ok��Vo::X�ɤniǻ�	Oni���'�&�m�*A�[�-�-�B�hϯJ�eI73�j��V媩b# �a�#���J?���E��=UƳ;���t^����؛N��@�r$襸P��Ɗƍ�d?n�C7]� ���~���j�v"vq��qY���A���4]��^��eh��821�pM��ӄ�)f�̧"�a�y�v�sb-Hh��:��Yh�Ȱ��N��$d��(b����Tn�۩YT�YŇ�;[��/�wlR1�v�T�+wC��n�;���1��^���Pᡂ�ͭ�^[I�m��p<��ǯ����U�I�Y������[��]�Ypn�b�f���v!@ʒ�˲�l����D����_f��[�j�e�b̗*n;�jH)�����X�[s2�M^���N��l<��	j#g�l�wj���⁮�|�7i�����9���W5���aj���3��`۷mJ7��`:J�����[�V�`9YE#ص�Ǚ��ΠwI����*�Ê��-�0S)MT�/vUY1��d=3R�Ʋ��)�cu���X���4�ݳbY��7���:l�U&]Y�$��h�!<���m���[N�ܖhK/o0�X6��E����d��T�4K�Gb����-E{vpe��ݽ�D�J��t���"��Q|�f���h*Ǭ�/U�g�e��*��*�թ<�wi⹊b V��7!L�N�U]gQ�_4��l];���ָm�.e�@H0C���2�Ȝ!�Fc�6	���m[r�	W�e���mS����D�H�TV��ɘ��"e�U�M؞�4���65��2��$�+�V(�l��Q}�E Yv5f斴�̖�s`�q�ĥ���ŵ�q�e�[�&^\P�&�� 	�r^�)�]��r�b��h3=H�l}o�����)���j��z1�J��[}�;N>/2�se>�Q�C�Z5 ]5H�wx�@�B��/^f�n�^�r�em�6�c͉�B��Ry
���Z��љxFX4I���K{3$9�[��ɻ��^�[��*v����J��oz��c���'���z�{:��v[��	40��s���}���^�0r���4�5�H���&���W�ն����d=�!��$�r����IbN�N��;o�7��2�Sj�0f�A����J��{X泛P0�z���-2�U�Ƚ�?nL�xq�{j��N&� v�.�@D���4bt�_����V;�Я+X��,ȁ�e�X6ADйo&mqlcJ��7y+q�2(��/)����f��	p13sAY�.���	^��l��o�%K��C/��6��{�H^��n�l��Ԣ��n��H����Z���$Q&UQ�� �*A8�A�C,�ԫ�V�4�oe!Ֆn1�a�hm6�J�#onApܗNQ<\qSR���I��)2�����3�0*�8��I̔�DN"���݆%�%Y{Xn�[�aT�щ�Y��P�^�,m�&�G��*�E�y�d'0Źr�v53��D�{���Ѧ2��r�J�G�Iʽ̂�7�*�"�E��f����sr�Jx0����0�����ڊ�1z����g+�%���qu��c�Jg8��Wg��ܤn) �awA�(��a��lÛV�{�8�3)�fJ@�4�k5TqiD�2�WIm	��U1�5aXByn�0��GtL�T��hk�Ic���)e8���]���P�A�5�ѻ���!�OD���mS�[�.�c��Mna�����7[��)Q�Syq���6�16Awmj):˰e�&���L �7.ee�V�԰��-���}y�dX��^�em�Y��-�,'+��^6��o� eZye��(�yz�SVE�)�ŷI�Y�v�G���R������/i�X�yz&�-I0�ȶ�8/C��,u7M�ݩ�j�j&�9�FԯŦ���1���X��YX~�I��o:�<���8.X�]�VF���n�ͲZ�t
�ۖ��x%��h8�^�q*�m�Y�s[Ė����ֻ�gL�3,e�pf@HZ#Jɦ��� �VY�r[�pP�t��V��hR���q���|,T�.V8-	%�J6�iD6�
�?`wG[��xxվ�ȭT��Ỏ��l�w��g�ZSk]���7gt�@6`�B�Ӵ	��R�*�F	x&��v�zc���X�!�:�ɡ]�ǣH����!���]���5E�$��!��H76C�vVڔ+5������FfH�+W��zʙ19�1��K,PN��j�t�_�t�0�u���.���D���U�*�Fc5Y�����V��PRb�иs2��m���f\ɪa�fdB�zT�i�V�c�Lz�b��c7nڄmd�lj��)�8麽Ndxle4Fxf(�GQ�&�;Am�u�f������ q ���Z�4��8�i�8���a<�@�͏47�3Q��Իj�f�����]2�(�����v�a�Y�l��DGCEfc�� 5t�v��e;�SNL����T�,h��̴R��#X��ݎ�����j��Xr��h<w��V��F".L�NZ�̢u7jj�d*��F�eK�a"rdKD�&��Υ˘)�e��V\(��F��܄�*Z6���ڂ�@Cn��ݭE�������t��݇�Yq�����4!�>O��p�J�kB��vצ�0�m����u�{����Xy}�QT����q!�X�c��8O3{�N�ud�cH�4��8�Ӕ��i�E=���e��7�%�b�2�.�f�a�S`��gۨ�*��1�ڱ�b��k4�fV�K��eM�Ao���N�iO�)�^�X�!)D���n��%��>N��¾u�z�<S>5,���CL���]�@^Z�A"���Y�w#��%�e�3uh���I�:2�t�Z1 �vwQz��ȋ��fSQ|�^�
�{�x؇:���eT��"&�klYD�����c��L�����نL��L@�N��ݠ��XP%��H�X�s(�
��?fA躕z���U�8$<����9�8���jƊ]�p�gP�oG��|�p��T `W�m���S�\:-E��LA�������||�vS��$��I
�fCp*�dW�+�6h
�)�8S�Qa�'�� �Lo2a��bo3���8��mΊ��VQ4ðL2лr��T�7G�Vqnf,-��fS.���	�����@; fnRzqU]��(�k��*[�^a�	���%�����-��u�@�NZt��H�'wnbT/�ˊ3�[��ڵ��)XB}"�b'X,�DO+X�ќ6�޳g��6-�� �k�̧srLۊ�b�<�+J��61���R�l6�ՖY� �`��;�X�w�6;d�d�7#�9�*ц�v���VXͬ	���/���t\ yh�:;~O�^���k��i��[�ygF�����D�g3ײ���!.y��r�N����R\�	c5`rR�hn"�ø)�N�@m;n $c�]։WWf�[�e��q��8�eX�؆x�/j�����q�S������-��/^S�B��`��Yz��V)oq�mH5�[7�ْ���M	����ΦQ�3��B�iH�VN�8,�R�ޕ�c����1G:H��Q�`�4�A}�z�83�����`��B���1�g5�j����,�y��e�;X3z������L�z��,����9��M��+�r�;�f�}W�z��ie�Z�,�@ީd�TX��d�?O���}�?@?�F�[�a,g���O�%:�����2������m��s�"Uy@e9����E�J�x�5�*�����x��i��m2��L�eP�x�@G9���Gֲ��.ƌҝEK���P�O �s�>�9�l����t���N��HV��v�Eɧ9WS���YY�P���5�+f�p|������L���B��)����n��$n־�}&�������]58���S��)Z=ɠ��*��l�XB̥\{�1r�=�Ȕ��;ugCW���J��qڧ�T����E��=Jh�t�\���k�X)>y���!��>�0V���dK5i��ܳ�Fژ�6K5u�'[�o���z�s秂��D�l�9�bl���V�b$n����Q�Q!�w��ZRm�赠�ݺ4!�^p֠���� ^M\flRҦ��N;�i�TN��*�V� V?�m|5ĥ�6��oX�tvC�%���	�14"���ؒR]����Y��c��u�הn�k���5����W�-�<������]����RBa���PT�n�>K-3i��6�^�h�����^aUց��:�ɍfJ�P���˽`N�iyҭ�m�7�}�KZ�����v����Mb+u<ҍ�ãl�"�S�ɥ���n%�Y�X��ٺM\��s���ס
��)Jٰή��nN�7����� y�be�䆾L�zJ��wj֧3���K����*l淗�����ѕ׏��na}`�kocv����:����;��u�r�n�28�ά#C3G�"M;�sY����%s5 ��ڳ�WE;C7�l�k�AM��	�d@^�Z����y����cnL�	V��ݧMp��G	���C��$�s�����op3��\f�|��M�J�.�����K�m����6ef��zڎ�>8ګ�9S�ۇ^f��ʫJuvs7D��\��o鯆��a��]�܏�]٫qK#�l��\�s�|�>J��L��g:�%82:�,��p�X��o3֒\��
�t�{��8�)��6�e�F���m��L�]_q�R�X��k�|6�#���
�:_r:cGKlkS�B���U�{]�����Cr��?NԹ�{��jA��4]	Cr�բ\o���*NS&��׎,r��;�=�}����*�F�o%�7��
m��ʼ��j<CS:c���azE��\��5��3_:x2�]zbx���G�+#5�!5��i]_��.^)��{jv�fs��fZ%����Y���������0���p�$裆�$U����M�×7y+ݽ c$��^B~�T:5��4�*P�t����M@<�7wO.��ӡ��E����|9Y~j�*cq��	�O�l�H�o��3A/7ao*��9���j�aM�k����xD�f��V���Z\mb�X��Sp����*��m*��11%U�r�����롵�ȏ�� j�m�of�0u퍔e��>�Ǖ�`h���&���{��t5�nU�.d��>.�g46�N�9�SJ��Z ���7�0Rj�4g׳z'�*i
/n��5��J�vbb̽��2�l�r��]7K��e�0ow)��MK5���u_i��l����;�\E���tmLw�+���	���]+7�9�'Ir����a]����51����C|oa�NT��gQ���|���-��ks*������%��jv!�s�:k���w�f��N�U9Ӎ��K�'�3i�ZZ�:�����8�"q�(��J�kK:�M��0X�]
+��gs�Ц]՘.M�}h��{J��1u�7���:�}ʁ���$��ղK��9\olV�
�"���w�G���i)y�����؋`�6�R�����Z���:��칧meE����ш�2�������M���o1�Ə��VI|[?����.LF��z�&�����b��[�6�PP�L2��2�!���5�룙-t7ԍ�%�K�'}���������Y��%Ê�����9�CŃ��Vs3|�N�7wYHc �y��+	�����I���ݣ���D�[1l]0�T{�Z��j;і:�+��P���u�C	.X�H���2���W�9�
@�!�[����\�Ț@]K�L��R����z��i�Z�b���9�J�3M�s��^���)�[��pu���v��I��I>'�`X�F]�)eS�����:�u��d�bW����C(� I��ㄻn<賅I�����G*�k��]r86Aխ��H��1�Ԝqi�+�ܩ�h���3�:M���=�WX�r�f�tb=3tq��R��u63��m[�S�f�Τ�MY]r���q����l��b�O(�R+��1ٟL�`��>{/��o��]��;JK�s����	i�;7]F3�c�6-B, ;��;}}ɷ�Xn+�B�q��s���^��DY�R=�SٛNl��i�a3�7Do�'�+n�議�/��N]��H�+��J'wX�dd�k7G�A�#�A���Θ�gXG�2�@��۽�"�i�D�S�q�s7o�()\��,��9�jS$Z]�I4����[m�W���ּ�m.5&Y�(�ɷuͲ]���*�O��2��U�S��a���"������"�������:�aX��er� �$�oT7���|ٚ��qŕ�ij�y�	ن�.��۾d���ɪ�X��QK��+���TGR�*����Vi��w�� �uji�r\Zp�[4�b�d5�����ӻ�C�����V�"��,�:��<���5�}N�9�}O�A��7	P���Ζ�:��H+L�k��	���S�yl>�4=�U�����F���5�5Έ�c�L��lX�N�|��H��S�֥��^�ޢ(��r�+sF% ����hH���usV�����FT�����c�(� 9k�\����N�s����}6u�
�3��wf���J���gU9|Vy:�;2�1-[���:���:j�b߅-o��1E�5�rm]�N}X�s�̓fTh�^�����
J��Hu,�^<�O5�>]�+�0�L��M��:Jk����j��_t�b��l��**�N�AU�u�ѝ�9n��2fIa��2�&�U�Ay3�&�S�[a1�`��ru.5����ۂ��E×�����k�*p�7\��3R����h��NEj��*���yDb���hcПfG��������Ⳣ�l�ڼ�H�eugwLP�BXA]'Ü.�֯��Uգ��>��q���q^7��-�]�w�Լ�@B�;c�M��LP��Qp=��ቫ�z�}q�.KOI�6�p[s,�����)[�-���܉���:�]�4�Uxv^��R���(j�h�G��2���ν˰�]X\�qѨ�����*#e�X˺t�&����J�X�Q���t����0��ΪQ�����`uX�\Q>�-鸳�vԮ1.�����u���K%�
YK6f%������6�7����VX���ͣ�k7$Ư2����e���lZ\�b����,�Ǟтԉ��Vʗ�(=�ή0'ó�r)�r�ːQ�ѷ�ٕ����>�®�^�U��ƣ�w�I.�vfA��Ge��r�p���VW"%��i����.�=wQ'00H���t��Zz�^� wR�];�A���.��Ք�fGj��D�t�|�� ���-��/��cy��������q�I��Ҫ�`g�`�*ފ�V�历<A�r�f�H*� �t̩Z����^��z?h�+׸�请D���7�!F��s�O1�.g�@5�iDq/3��U}�uk%�쇔�U��]�dwָ����4>5ӌK�bMYmL�%��*�T[�B��}�h�S���9�棙G3V6�r�%ɫ8��h����1��D��Ѩq�mk̳+d�R��W���6j4���n�n�fW1��ӗC�h�2;w���4o��*��+����ǖ��U���ѫ�]��Ǵ�h������8�ث^�������<��]���2қ�bQW� �ި�r��׵N��~=�z�]6��_�c�u�`wÈU�4U��)�X/�S�Jn<�]5+�����v)a���X*��ہ��(s�NJ,vy60�廠*V3P���f�<�L�ܛvw��8�QB��e�_9����E���6$
-�ǲn����n��*4wL��k3r􃴙^:����ֶD��B#��I�F�̫׫���oEy�a<s�n�k���#@,ݤ饀+�x{g��u) ��dX�n��c�S�eb�̾��e��u��5Mfփ�v��gU�mBv�\�g3ub�d�p�~�7h$��:��V�mW)��l^km��sZ�ox)f���=�ۡ��U�< �kF�DLc|��{DbwJ�l�{s3v��nl7J)�u�0�
�	.�:���n�{�^+���j���7ϐǥ
��.Fj7����Zq�h�����>&k���gnHӚ���w��v��3�mZ*�鈙��6�'`Ty���=��G
�-m�-��o��͂¾PK�s-d"9@�iỢ*�[SD�.�5��ks8a��6�pH����i\B��5c[�kWj͆g��q�];���o+�CrS ��˩X]j��ۂb}��|�]�Wj��'S;�]��s�\�Cq`sPE:�	���7&E�T]h��$V;����W��h��U��	ˠ\��4��qt��Lf,ݺ3��bq&��NM|:c{���&@��i�X<�_gon�twr:�� ���ż���j	[`��Rɜ��q �Q�Ƶ�î�@�k;�7���U�b�s��u5+B�aʺ
Lj]w�#Xb+Q��X�}|*2�4g�=o+��Cn���HRQE)mށ�FsL�C�U��Ffє%��׳HN�`��x���Y���;���yu�<�T͚Y�5ΞX�#)�����F�i�Ncs�z�Z�˕�7�~Q�]�clh�[ ��ǐ1l�\���Xj�(̷�ڊ�ha�l0�u0-:3U��(�	Q�"k4�'�n�,���ob��M�6m��"����dԵ|{y 8�p��K"�(�r�DU���dR�ܣTrg&,����uہ���0y��b��SSx%�c6�j�~��%Z�����'O*i�0;t]�O�!�����{���>�R�g��bx����z��<�]o�D�]�o2Ξi�8��:����l�����pTw�]��p�4�����Ч�1[��pZh9˵��f-V�MNfW����%ix�sfrΡ@b-��rN#wo%*g@��i���6&ƭN�!���)j�4��pq]� ��@T���ҩgf�a�C1�q�[د,!�23�a��c52�0V#k��Wa��-�Z�쭵`5*V�g��� .���.[-�tT]��h��DŲv��z��w����\�I~qx�Su]к9�����^�&��}�n'3�:�iT�<s��@-��ˣ
ܝ�3��mn6~\ZV \#
��e�nIp]r�w��q+r�w)�����ά��qKR�V�l�U��R���H`�Y��Ƕ��g�XmU��y�%���q�a`V��b�[i�4N�|��č�xݕ���i�+[<��[��kk�nE�)\/{k�^>T�*t3i�9a�W<�Bs㎈��N+�X��ҙ��;�ݷP��o�S�RG	���m��Vr��5:�ڹ��4��f�*䁽U{ܗVոfAXj�V� �FǨ`Ð�pؔ�����+Ƴ��j��Ո���i
+�����:7>��֎�q���8f��5N���:�H��NWl�6䕱M��J�AHvd�nI[�8�]��cۗ��{f�;C8Q��� 0[ܷ C��-ʰks#B'!U��y�ܚ��΀Eؒ+r�\ja�Ob�z��x�8�ý��q�w&}xu�6�ސ���m�#�ȇL�Z\�$�IRI�K���`���Y��ۛ���P�Dnkp�4��V��	�'oPjb��w��V7`Ō+$�\��I�blY�AM$�_�2LF�&��$��$Fa�E�M(M��4���"�	Eʁp�ܪ�ʺb�&�P�(2�b ���t
sR�')��+0��IP��q	UH�n�R� �Ir-��)�0�i$$p'$�����?j�(�JBb �	�I�Cd&#k�c���T$���l���w �NMTW␦@�΁@���b �H&�L!A.��1F��D��7?/�/ܟ�Z?��6�Q��ҒG�fP��*7�J��-|�PFhK�wa�H�,�ӎ�-�6�`��#	 ��d�c�D�1���*PT_��PpK��pSnR	�UZFʺ�h� H�FDU�FX1�L�{bC gP�D-�l�ʐ�_����BO��	��j7�~8Yf(A	��H$b*J"% �ΆԨ��0�HH�06N�'�e�*��&���'�H���� t��[5u}���F��:f��ɓ
VJH6��q�����fC	SM~Q�[1�d��D �@�La�h��J- E"�H�b\FR/*D�5AT)���`u�}�W}���xvx"���ۈ ��~?����?��D�\�f��go�y�⦒��Ï�p�м����G�|6���;J��#2>�*��D,�������J�
�o�	˼�FK��H��o���7�+9wAU��bŲ��n�p��)���C�vJ�����An�]�hћ�yXsP�̭��8=r������t�S��H,�n)sި�;1=X �WdmN�f��[6�u�˳p�ص���{��B(ø��T�w���Ϗ���-��m�ǙY$���u��fW=���K�.��+5v�4Q�(���r�Q��>�I��:WL���v��JA���\�-��.��P۱Bs�*�~E�9I�8�BLvo;+w���� hǩǔ:'���k�Ōɻ��j�i�\�����Ff�+6ܨulu�e..��dq�Zr��H�[F �	�.�}��������2�Tw`-L! �*���賨����ݻS�YJ_�w��:��֡���uTa�bttr�\��˥n�����9r	�wة�W=ޙ3�VUq����[�J]�!�L�L���m�L�4�S�9�,ѭ�����|�T#"oq_g�+e�3"E�|�]�q���n��R�`�>�ʧC��؛S��S���|�j7�$�Ӭ�o���];�F0��3���[S�����׏�Ǐ<x�׃Ǐ<x��Ǐ�<x��ǎ�g�<x���Ǐ�<x��ǏǏ=<x���Ǎ����M����5i��y�2$�D����#�h9]Ӄ�DK��9h�]a�Xs,0�i<|��*��%eu@�ܮ5_7ic͙Ze�yR�����RN���0t�;�*�V���m>:*m���M&������*��۳mh�w|�47�qq���_d���u��)�ͦS��-IɧS�Om��X�PR���d��nD&,��bT�h��~$1{бR��p�'J�f5e�ζ^��P:0\���F��4�7�axC�.Ftm*����5;.X��
Q�81�>�a�꽻11��,�K�{\�Ӌ�[ð�̹��Th���;:����ɐ���w6�8��a<r.��t�������[��z4wwdQ�S�U��$�d5*�]e7e�Si�X���).O��tԬYx�щ�9[�6m��zg)Y�r��ǌ*Yyyc6�3�ze�i`|��Y�[9A���yœ��8N���]k�Ϊ��}�b�r���h2%��n�V�d�{����z�7W�n� �r�څ�<��P���;]���Z&'��:(�F3A,���.�1D��?�	����Y�q��G��
�Gx�k0��!�h1m)*GNP�ϵ`R�d#�.m��!�Κ[���k�|�xAT%��Q��=&��s2*:)����i�����@p�Xq)"�y���9�dQ,㮶�U��^���~^<x���ǎ<x��Ǐ^<g�<x���^<x��Ǐ<<x��ǏǏ=<x��Ǐ>�x�Ǐ<{mmmmmimmmd���%��]�h2@���E��U'�m_bOr���G����C����+��s����6��A�.���`n��(���c+�-.���mM�^q�?��E�q��ﻴ�}Lυb��8t^��������]	�7L�_}֭�dd��]_uV�r������Agd�rY����P�Ȁ�

�(:m�,��Ke�,���TD�N��KA�E��J��7�>p�[��
�>�k����W���z�r��{J<;����H�H�?G���U&Z@���]$��d�%ىj�ȓr��Y$n=@`�j�m@X^"Xͽ����$ɷx�^�SY .�pN�,2������N

��-:@�N*��W[ �j��V�98��˭��A좣y�7Q����G��쪋�d��]@�i�vҲ  A�J�PU\O5I������Yl�������1�!�a'^���Fw*�勍�[``nQ*�N�g
�����т��:\��Ł:�NP�6꾦��޴y��5[ۖ:<M�WWS[�wEʞpd���y�cW5�V�JI�]��A����
tk
ar���ۼ�3������\rjɛ���Z���9�pQ���v|�&��f�b2IS6�7}�A��:=������Rs�U�֕'�/S�ie���>�O��W��D�Ƿ72�\�f8O17~�����B��t�8',wR����u�I���Bs( �W�;#��z��į�кc`��-tnð��>���-�Q�U�%��w���q r���yV*[U;n�s��������]���S0��c[K[k;SckckkSkǏ�<x����Ǐx��Ǐ>�x�<x��ǎ�<x��Ǐ^<q�Ǐ<x���Ǐ<|x��Ƿ����ɥ�
���[�K>���:��S"(PE)HG�-*�X5�q���Y�@�2��͸"�2<-u򾫾#L)���	64��Ts/�ض�g>a�C���+賺Sv)��]���:���7>+8���h�VuV�,(�p�H������ ��)���-Ahe��rk�t�N^ϥ��p[c���+unmliEG��$c���U�J=l��4��"��UK�w�g�+��Q=0N
�]}W��<\�O��f&�k�t��֕v�.��c�e���̖�Υ�����A���=×Mv-���r�(`
|�f47�X&�Y����0�+9� Եd�M�Ƶ�����BWmt�X��I@�i��ʖ3"a�\3/)
B��:.����]�H%L�[}�&�}K���s m7�l��Hλ���Ldgh��-5�E�gL4rSu)[.�ǽ��tU.�C7L[Usk<fr�dZxR!y�.�B�h���%Rp���y^��b�{H����ϳt���z>i�Ω��		�c�\!^Z�{��Z��4�f�r�gF,�I����qz	ޕ�b��G%�Nj�_*�wHBb���>M���I�ʐ֊.P���<:�:WRU�xgfxUhu�fg*r8�X���(m�f��
�=�����<C��1���-���g/��.�P�k,M�+i�;cS[cCkkkkkKkkkǏo<x���Ǐ�<x����Ǐx��Ǐ>�x�<x��ǎ�<x��Ǐ<x<x��Ǐ�<zx��y�o�+���t��
�V=�*���9T��C�+��i�W�ajl��m�D����b�8��sQ|h>�Yj�\�
HA��Z ll�0�QD�vj�zU�gW
[
����|�ჅsL�s�U�h ޔ:�Л�C�P朙(=4���:���m��Հ���cz�<d��v��t�L0��e���k�E����]��1H��Ä�<ݍB�,�/wue����;-����-�N�aVh������D�@�D�ؔ�w%͌��N��a�-���[�S6�` ��^�-��+�Xmh��M�$�����,�S�v
�-�Q	�MF
��55:�X��ݶlr!`���z�uD��6����R5oq�� ����H�E�ʻ��_R�gC�(^ih�\.��t��V(k�z���&�f�/�G�m�b[W��ǇO�����#���h(�P:�t���l0p�;5�ޔJB��|�:������ B�m��X�t�,{��wGKG�'��]���0�]r����v�J��H\#�TC�r&�̇�΢��^љ�9��)��l��w{�î����@^�٧��'���+��)\S
��zjܓOM����+�I��-�w�
F�ҏ+[p�-
�2I��^���M0�C;Kkkcx�Ǐ�<x���Ǐ<{x��Ǐo<x���Ǐ�<x����Ǐx��Ǐ>�<x��Ǐ<x<x��Ǐ+���}>�O�ײ�&Rz�K����O��Aq9[@�"�ݝƱVR�[�W��}ΐ�1�2�8�Jֺ�,��.yƋ�>��dք(۝u�a��؎#�����m*ovs\N!h�T��e�����弐����yк]	�dEiQunt_t�j�bݺ��2���E��&GF�Z�r���%�rd�iV,�;a����bώn��zR��oK	���\��@om�`O�R�tL��"�v\ٕ6�[<�=e�YJW�Zn�� �N7:�3c�;���/2m�'%�"�i��Z���׉�{jD*�\4�(�Nv��ң���l����[F� *X��Ö��)�e�+Ga��o��F�M��tѥJ�b�+&��
�u#_&��p�OHs�T��i����(rvR��nQ�4��*P�:�osr�qOJ�����q�:��yd3��H��fc��gh+�a�����m����H�q��8u%s.���ئ��P�Ub�a�W-T�{�;7`�F_X��6z�^H҆�'e�+#cv���z֭�v�R&�hz�#�N+�> [|��=��.��^��������n㼜��]M�\K��~��g̪U���Z�mX����\G�PmЅ=?�?__��x���Ǐ<~<x���Ǐ<|x��Ƿ�<x���Ǐ<x���Ǐ<~<<x��Ǐ<x�mmmmmmmmmb���ɓ��.�Y�R�@H��+�!t��Y&�}(
q	1�T-�.K��j\�R��#o
<��v)�%k6�4�
[�m���ҚJ9f���l��̱�FՉ>�� �6��a���[�;{��^����o�]A�F	mm<���2`Q���Ќ���o�
�ɀL�2��yIg=p��L�\vʺ}b�%g���h�p�y��e<�]Z��M�[>��Zh�N�#�2=�y�٩f��@�� �H�g7��q�Ehd��
�l'�ٮ�V�����`�o�e*+���5+f)|��T{�_�21�o2e��H#NX����L{s&8]O��;�9\ew"4���d<;ǂ�>��rMd�e�Ggz��,���on� �y�͚R���>о��L�x�ε����P�ݣ2����Q�*�i�29c9���5}4�0��qݠ햴�}(Xt,�j�.u�u�9h��z
aZ���vo�G�������'3��M&蘖��r�OP���W��p�O,H������/��n&wkL2A0���b��(���j���=���;!;�(R/zDNֆi2����p^c�z�.v�O�_K]�ô��qun򸄗�S���t�����']�Ī�fkn���[CSC[S[ckc�x��Ǐ<}x�Ǐ<x����ǏO<x���Ǐ><x��Ƿ�<x����<x��Ǐ�<q�Ǐ<x�������n,,;1nB(H&u����W+���Udŕ�q\�S>�;]�c`h(+�oo[&�Vvd�43�aj�$�������t�y�X�{P�[�)�p��Y����okD�q��� �7��Cz�&�;G*71sȭ�iS��p��;Z�a�b����2���$�m4֮�w8���cf�������NRa�F�De���9^�nn�@a�ͦ+�RGx`�*�`nK���@e���:�bG��Ae�I��
� ���8+������v��j@*�l�h�C�v�1�K�¹�N�;;D޽t��],61ջw�pF�6�5����a�"�u ��$�t���+�Џ�i+�/�M C�Rj�]k&庆��7e]&��V-w6�����ljp�ƪ�N>��O,�z9�3��t���:e�uVp�ݑl�c/X�r;�/�dԻ��=���V"�EL}-޺e�u��%sqnZ��)V�L�v���}V�A�w�5��y����$���L�&����:^�j�=me'.�s%�VP�A䏊v={o�o���ٝ�Ԉ��(.��n��4�VH�V��33��҅g�U`�보I&}Wi�K*/(�j1��Flv�s��-vVpt����1r���U��h�hYM--�-��m������Ǐ<x�׌��Ǐ<x�׌��Ǐ<~<x���Ǐ<|x��Ƿ�<zx��Ǐ�<x���Ǐ?<g����\�J5�r���m��9g���vX:.��̗,��K�=�d��e�@(��y�g��%V򃮏���h��0��Z��d��k�E�ʥ��8��#��Ksl��h�)����
b�R��h������a���oU7Jνn��`����7W�÷��Ɲfeʳ��8��{5�/�uL��óeJ��[僫-2�u��˳ZɭjEʭ���\�=��μ3����>:n�d�ټ��\�A��V\�
��yz".��$��[�ڱ���"�a.��oV6M��N�p:�_C����l�5��U����/�;���rܚC��,���P�;�΋kT�ZƳ�x��.Mz3�ӑ��wP3��<�SE��-�5���2�1Iõ�t�J�g�v��� Ot�RY(Q���h�#�7O��oQ�`ܓ��i���ee�:,�c-X.����D��U�J�u-cv�U�N��3Bn�"����%�v��ڙ�w�����w�*��ј�l*���vZ�#4�Nb���YwY��kW-��wsB�<��U�Æ�;�fL���y�h��h��{�[՗yR<v]کL+M�Wp{Ї���ѻ�F!jIu��+3�=�YLs�����t�}�.
#��3[]M��H���|�4��ͼ6l�v�Z�ٚ�o	�դ=+u�S(�Ѻ]���qo1�=�^+2�&�z�ئ^�
��l��|*�X��/CҞ��!Z���˝	�N\���f�1K�,�5�]k�frO��b��:���k����f���=��,M���c�|6d�D�]cJ�L�ۤr�y�	;U��2Һ��/U%��\[,�b�#���fh�x�������QM)ӵb�dK��7)!��4clX�[sfEU�Z&!֣m��'Li���ף':��}�β�d�ot1kyⴱd���yX-����#�'u� CngTkk�o3�c�3G9g'2�-h��^�j9��b ��:�ټxqb�אr�I^�9�Sj'Op�����G�Z��j��GL�u��`���;�&սwp:��fj	^"�o�Q��l]F�l8�η��Ar��{���1��V����<�+���mK��ǳF���KxH�\qI�;�£�e["�Gۨ79T�7YzG��!W�]��n[귢ӛ�SO�>$�W��s�!d:g-`K��+
\��68�Yh徑�*\b�#;/���F��rC�SN��7�fD��	Pn��/��D��URx�un��wiN�r���w��D_�����o�����x������5�߳;�e#T$Q�[��H�2�H�RQn�I7L0RF��I��&��PU`�$)ӕd^���Y7���r2"�+z����z�;�Om�ȹBZ�P$��W���$�f�@��RI�|��Lޣ#`,W�\Xaǹ.c�Mk.�;+wжʧ��n�N'{p}������{����ѕ��`kE�g-(�*��TN��2�-j�o�t<3m�Aq�/VoN"v�U�b��ɷ$̩x"@�Y�|�U��v=	�>�0ЬM��Y?TB����!j2�+��@�p�h������3����"�P�[λ��E�W5�L�r��Ku�,�R��hV�sq�k��-d��w������:���}Pky��.T~����H��q��]ړ�L�2�6Ό��O���].�Q��U��/33��iU�'[��JķxX��:�,�)Jq��f/���^(�9��!k!�m�6�˭�ep�tm�[�)���9t{�w���]�<��a�����������aլ&�T:� t��~��h#����=b���j���Ư�������]���,E]b��B�9z�4j�A����ҷ��\M3p_Jr�ø8ʽ�`�a�e�
m�q��%�]��ǎrz���Ҙ�Ɓ/1��Iɓ:N��+�+��P�[���f�B�1�dH_&�2b*�f���_�M����Dƙ�[�M�.��M8[0��!�a���a�B	
e�"����b0��h���D1(fu�du�ٝ��	�1�=T���ԧ$����B��w:����]u�C�'Rw#�'P���:�b���X0ް�0���"�"�&k�L��]MU_���]u��u�(��
b�(��`ɤ�I�J�@�����0��*�
iX���*JE�p�%4�9� �>���4��Ef`0��QO�TTM%G�ȥJ����(*�����dUS�d?;�:��+�p��8���}u׎�<²C�:̬������32貨�yaq�U=��S�U�`�rr�2�H�2��&��ɢ�"jR��{||x����8p�2�f�5ԙ4'}cK�g:ȃ�0�����)�.� ��+�;���&Hu�)����ߏ�Ǐ>�G�ʐ��'�y�����A�w��D�n�
|�è�(���C�^������Ǐ�9��:������w�u)A�/����:��I�9L��{x�~�_C�O`��)_�IAO\�<��9�#J|�힟�Ǐ;�"|��f❓A��
o1{����� �;��)��D�GϘ!�ܾ�����N4�H_����c���%�P���\Ho'�10�{��Jy�7lj�7w�ͮ뷇׃W]s��{ � ��G$3�_�QW���f��G�T}a;	��t7�>�l�����gT�z� N�zo����N٢fcL���\��<T&y�'�*�ĥ�δ#�O4F��$Tij���@����1�����G�}~�����
�+�0��,Nzk����} �@T�n���+�}��uYQ��','x�>�Cf����c�f���������bG�C�ۜ@��W�]m�ߺ���ܭ���*���d�s���G��������Ƹ�ӎU_�F��3�y����i���[�r�ڮ}���c�[���*=�s�>��}������lIQ{�[�O`�V�;U�g5��ch�������@�q�kr�oc����azDGm���X��� X��!}w`��z��NT<����ޢ�=[~g,�',zm�����`u���Ͻ�����DY,�{+�P?u�W.f��mf�$;�f�z\j��<���Z�a���~�lH�Ϧ�e:��>0-'*���J�-�28�h4�DTJ�r�k���V7�ީu�oqeb�̓��p���fbX.[|�r���H�v�b��(ԝy:͊=4�d���ǂ����I6vt3�D��ۈ᡼+=�Z��w�$��[�#���ږt6#}���v�;�r91���|���������~�{������نK����urU#�zGԾʊ��']��6�9G/Ը����>��Ww���Vt��u�N�����P��C��B��]�ɯ�:?aK���渟��������{����#���*S��=�e���l��eTtOJ���#��Om�b`�l�nӷW?e���+�	�B�NW�m��ˈw1����G�^��z�(7=�;v��j��ޗ��3��Nc_/�ZEN�8���ytz��<qo�t����N�g���(�wo}��a;�V���A"r%�fM�K��A����X���{^����G�����[уi;��xa�����Pku��U{l-���b�RY`]:�ɴv�'Ji����S���s2�4�U�8�Nh�u�k0%�"�t��(^�$3I0Ҋ�d��:j��=��zNvLV��#�-Mٳ��)a��B���ṩ� �t����
��a�������]~�����ێl��|�+��Ϊ@M/B7���j���H
����X�t�X=�Qn��'������Ax�>�Lz�$��`r���SWo�'{�|Oո��}���Ӭد���g�簄�<*�����U���?>���P�XY�GK���۵���������ƾ��rnC�>���x�n8�_�вp�h�����ÍfghE�O��|���#ݍ,�'_�Y�|�]!V����
/{�,���(��ys^���]���j���r�,����a����12OWL[ʠ�����X��dع���E�l������{�T��/$�+��c���L�Y}�}���r���^ޯT���v��&�!����r^�ܦ�۶�xa����;֮7U{)����#"���{�G'm�:V��k�o�lY�EP��,Y�h���׹:zt���JW��I� �G����������7�R�#8Ƽ�ܱ�B���{�8}5_�o��;5-]C�t�Q�*��'wC|�J���c�*�?�*���.��i�q>bKݰygï�y�f�s= _{�*���뼰�������Y�k��"84�j��{�;ވ���*�g��.��[��Q�y�3��5R(�V緢�����罳��9����w[E[i��K��v�#k�����=�I��cnK96G�G*ϹuҾ��co�>�դ�s��"�s'��{\�j�J�?t���mw��;��p����̞����y����Z��-�Ϛ���`�;�����wĎ�:X�m1؞	�����y�e��V�j��������҇G���9���X���3ޚ1~}����4"��q�&��@`�>�)��P��k~��,ˏ^Ĺ�Y�晓վdҎS��}F1S=���mOL��W�]�j9P;$g;�Z����o⧩)�O�)�Ot��]Tvfv����~v��d�z��7v��5��K�d+�S����κ)�Y�Vt�j`zMnX�K�
�SWQ%�����.�F	��e�(!�ۣC���m�g$l:U�����������x�k�����{JS0hg��A�W�#2 �6���ϝ_��j��,��T�)�J��q���C]��AD����Q�|k������Z�!2y�޻�ރVOP{&�(�֐(�g%����=خ!�V񺥓��=������i�<Y�E5��̓+��	>�^�&�P�� xһ��v�T����4�zo�RR�,����bf	=���	�L�ol-���z�ur7�1G���\�g�;��V���i ��gi���i��#z�:{k؁4*�:ߚ��&���5��)9�\���������W5��{��{�@�5�*y�=����}R:��&����K܃�<Z�~���M�ߗ�8}�p�������Ms���	�u?���M��O��O��3`�;9�s0�}����L��$���- 4d��=�I=�k�Ɂ��8w��/��΢��F�������:}�/���[}Sڍo�17V�
�t��g�p!w�����
e��I1TB�����U�˰�*{���36�[�o�8k�WaE]�Z�qe `�̵���;����q�������!�v֤�t��w7���d_V���A�a'P$u݊���&�����s]�E�ۘ	Z[ɻm�7���.M����EC		K��f��9���6����=s>�]E����w�J�c�5���X�#�
���gA$��ׄ��T<�^�Tc�����s�﹵�<�u�{�3~ZE{*��'l��3��O
��J�����r��䜬�Ydh���`x�@f#!�[�"�ߢc����vޘ�)R�����Q��4Y���FO�b��8h��i$�x��ۭ��}�3̼QM�\��Y�?_Ӷ;�Y�A���U�`�A^�-����$����� ��:2��O�ݽ��kX�T􃢜�x��?I���]�i�-8�Z2,Y��}W!���AX���y����Z&�D߹G�=���t�z��Jr)�8�S�V����S{��{ԏz��<��=7�,����3�==#�S�˪���*��%�\��c���BkNw�B�^i�c7�aӔ�y+��zn�Ϻ�\�!NbݭcXkFcd}ǩufo�Y֫e�V�Ī=la��k��E!U`�6
�+���e�9��^s�]�1I�6�< eyx��4��o@na�ޗ{�y�d܀D/���K"wٺ�9J�l��
��87k��:~���C2�v߽�~�qvt�M�����=.&�������P>�S���i?�=��5L��-rx��I�u��^�itLLt�/S����g���)�7uD�w��|穘i��u��M6���O_�2��ۯTt(�����2yw��|�y���{�b0�sy����KN3�k���bE�l����=2��+����/=��t�l�W��ud��D;��kС10�ճB��!{ >����f��C���~����:���9SB�>�=FT��n$g�`�3�q�l��޺~����=Zk�RF�HǱY��E�����U��^��J��.��9�.��~vq��j�6�ަ�-%�^ss���g-q��G>_r���zu+˅�p�'�����{�q�j{rE�zZx����t��q�˃n̋ޙebx���f!vē���rx��W�t���F�a
��6&g��0o�S�.�U�4��M��C؄&�|�����u{�B�QGP��!�!�u�зܕ�\�/D�A:"�k����\	�V�{j}��3C��Wf�\�sr�chU��v�b�﬜��yC��5j#_s�\{��;A�!KQK��XS��lt��z垮�7΅k�s�ޝ�
d5jf)nٲfVz�Q��	{��~�l�$�B��^���U�6T��i椵�M=�Z�N������f���ڞ�+�3dϢjdUv��#2�3�l�2;8�?�Kp^�d�w��c�E��o�����_ϡ�6t��y�ŷ��6�uu�,WUilN�ޙ^������_��Df���4a���&��&X�F�x���b�!���G�=�r¶�W�����L�v���7��I�i��/�mzwǃ�=�i�}#zf����ʿE��v�'\ȳ��쁴|/j�j�EO��lN��q\w�5k�:�t>q��C�ZO�	P�����v=�m^nU��?c�3� L�0}�׬��ff�Wҩ�^���>��ˬ��}X&�Ɩ�X7��r��f!ZNͼc��E��z=�����]�=�uaDu�X`u�����dD�-�!�@��{��
�ї���s;_d[M(�=6�_ݴ�m�Z�Eo7���f|4�v��۴�%�a�H�	�d Q ��`���(�JgIR��s�a]��c>s�����g��"x`E����<�
&�^}{p��'���geV���OI=����w]X~���l�\�aVa��y�!*{�� ��d%y�9o�����L��E���=��&����q�D�z?v�^��A�I픗��>T�ӷ���Ȩ1jS��s�Ԏ~��Nc��#X���v_?'
x�$�S�w''�:]�g�f*=�;a�98פt�S��F^�>q������c���a�pVP_uX������a9�t�4 4��է������������7~l��W���&�0�t��_���-�J���
0�t�h @�G��+�&�bW�w�ӕ�U�\���{�X��Dk]���J��;�K��\�L���_������o,�0rM����I}�5���/C���i�=�Q�a]�޳��寳�2��a���zu�Yu��?V��~��3�,�l���W6NB%���س��e�	��{a���]B]v*Κí�rgy����R� p�Yj�r�u�'gL�}�1�:�W�Ҟʩ��>�Vϟ/x�5�;T�g �������5�j��sҽ�*��:�z�x#|&�ܮ�Շݵ�Ou-�g��q�����4��ך�'/C <T��a����TW�z_�o����ջ��[Fs7q#�EO��m�\5�Q/~�����N�8&8�U��|t��yx3 ����Q����ϯ�퉾%�����V�� T,w�+�[��c�g��jr��Ok̿Ph$�zm�����],��I 
��?#�֏���s������<�z?
�)qӷ\����=:����;n�{>���|��Փޚmz�������c�Î���eE�᧿�V4�ǽ���s��a��_�o� k�(��+KW��(/?�}¬y����50��T�������K�u���w��բy]�=��S�� �v���%A�o�oOK�^Au�4�F�=��>pEӗD�ec]-��TW�v�i��ep������a�t�*ά��o�ڊc���]/9�pqd�(�|3op�V�M����$�k�ˤl�\���v�`���$J���6}��u~��9�U$	o�w;�[6F5H8��Nf�raNK�wׯee��^�wAM0c�A@�ƙ��,�So;��Z��;s�m����e�jj˵uQ���|���͙��#�B����k2�LHpֈhȀy�"�
�v�v33Vv��6�)1��L�2�a��[G�4VB��T��&��3\	^��`��:�΍���鰽��I{��'Zg� ޔɉr���.C�k&a��d�8����$
����)o2�Y=S��ƞN���D�+:f]Nݬy����d���L�wY�U��E7�o�CɚD�vC�d�\��]ǔXu����M��a�O �NN\�����,ٴ�$yk��_vn�F��Dͺr�8/K���O�tE�X3m����]3iI��ɲ����˖z��-	�:J����kdy����$�hf:Uz����Pv���oÉ�x �|��xG>��~8���Wch�.�\��4c�R9��;�A�3mr�y�&Pp<�5epg�(!�Ր��!������|�� �\�OaN�9������W����oHEu��Â�[e6�W��mI�o���b��3��f��D��9�𲲮g$oY��U^�U��7�XCo[$h�杵��5h�jڝ�l�(����Ų�=�<#�����C�E*ZlL�kv���̗r����	:ؚ"1v���^0�J�0N��U�5ur��2I�w�Ԍ.VC=m�|�nDo���;�����?�P���Ô�z���5��v���МR /^��Qި�J�e�=�ݧ�9��i�Yw&Z��܏�_f�FۈF����gs�Js�:j������⚓�������9W�geg>3�C��-�Z�R����˕�e��I@z�՛X+��������Z��V���� \�<RɆ�*��b��BN;;�^��[`��$��BW+<�d�߰輓�P�(G�r5��������9��FZ��gۻ�74�ˢ�T" ��xj3��f\�F)h�糧�U�Va<�Q��#�v�=�Um�v��dWig-D�?A˷�J��x ��u���m�6�0�<�>���Cս�+{.����	9��}E��\�^H��K�6O�EW���SM�,�����f�}2�
��E�e�X�T��:�qIL��8dx���s�lp�H�D	]��Xu�m) �����J'M�`�����c�o����_@��B�s��)�=����=�.�Z�\z{~>�x����R�#A]�b�A���ܔS��f4�A�IS��<u��P��\��/{��$h*���+$�L����O�x�{���>GO�b�`�ɕt@�Q�,�ǧ��^<}��J)�����@��H��:�(g�o��_����O���)�C!n���D�1㏏�<y��p��;�22\�JF������B�I���Ƿ����~��R�r ��2�����7���O''�<�$�2(G*O.�:��""�߯5ޯz2Bx�hk��0=�2�S�%o!��Cf^��8���c�.�ck�A,p�y3�:���YB�.s�����q�a�3�0맾��d��잉j`�ϣc�_�����8��{�{��~����i� "%i3�(�g��z����7�5�G�׿o�e�j�/��>��h�r2�`5�-"�{��\`sR��1�Ì{˙��;#sn;�a#�.�Δ�&u\�\<��k���N��M�B(!�q�a����K������t��u���Uzl�LZ���c��i��y��9�&�a^�	����(]�����	^�$\�(�\ܞ�5z��E�}jzK%HuE�gE��j7�����N8 ���^śD�,��W_�i�φ��.�0�sU��d���2e��YB��<3W�ßtД7�[��l��J%m��J��^΀@�x6���L��<�;�'v�<�1^s�Bi#���!t�ř�@�\4�h��eM,�d��9�D5�*5��o8�+J��qO�z����{��K��������,ńկbg�ga��9��ZL�b����<ߚ
,b��h	P-x�N��� {��tN�'.f*UІ�����%�&�-8��Ӳg!����_�N9�	�4�?Hܭ}�7"겵�e�HGF��3�:�b\�+�>��|\e��c��8c.?x�2�ZwFb� �����+�o�s�<�ʆ�_*Ǆ�B9M��u(��ή�2�����݇6ۮ&�S�	�"g$�Kⅉm���1`X�Q�L�&�L�2d�����%B�@��**���-���Sz5���t��xE���r6�Kz�`:�vwIwVo>#�{�8�َ~w����&~"�>L��52�x���?9�uJ�&kj�f�O�3��xWT	�\q�8�c6h�R�y[��
�M��쑯L�BXm
���i�[:ʶx|e.4�PǤ�#L���%8�=>�2��C��Zx�Ö,�����eJ�W3������ׂ���*q"o� {���o끐0���,X�
�'-�3�R����;*����p�ˑ��|�����'d�[L��\"�Ҝ��H U1�:��k�g�z�WG|��jz�	2)�u�j��X�{/Z��>�+K����
��$	���:�|��픤�s��Ω�k��6g���8�>8^�Y��5�)]���ͪ$Cμ�� �/B�[a�����Sw��xx@��y��e� ׼dK�!��q}�1͈q�T���:N'E�9q˳w���$8�T��D�z��/'�W�b��
Ƞ;k[V��wb��装I��1Ǭ�>�g����G��ۺ���Ou7�݋�T(�cU֡(�lv��I�o8��7����&Pp����*ei`����B&��.�����}�Z���������"
�l���Cvɸ-L{K�Z��^U��-�6�9�Gf������m�&�*	"B,"P���	
��yuW��俖D��f����Y�O�%�_/�;��}�{���8X�
A�Y�}h9��M��7@ډ-l�tCp(Y�O�nFhJs[�ޙ��j���U{�Fe�`�͇n�h�����r\&,�[
�-Y�hQ�M�lJ<�P��JbKƘ��
�0Ɋ��/V�����ⴳfx�v=��i����k���tʹ�/�8�m�,�nq�p�!k�Տ�|�r�e�ع(�b��_T�~y�{�5JR���b�A�R1�Q��ZpC�hn�����h�H޹-���Jn��y��R��zsCNΦ�u!��B㏾>`NW,W�| �X9�Ea20�N4�U��`d�9��y��mj9��y�8�j���JLe[j#�3�i�R����+�~�AC��`���"�Osf���,��b��jV^)iD`��ӵ!wh�B���DxP�w`͞!�>zSȗ�Oq��IH��g����+�ٯu{�3�yλ.�q�Q.mD�'� a����~"��[-Q'�i�˽b������:w���A>�ϥZ��p�.r��	�(tq;tB@�P���'�S�AM�����w.& Ӣ	7h�b��9wX\'���uV�N~e2�7�L�_h��U~���{~����Ti�[���4E���(�;��R}w+dyݱ��>�0�z��͟�2�C&Vu;}nJ����Lw.�U��z�7޺�����W�o=����d	�W �dŌ�0/rɐ�"�RnX�HKk|�9�1�j~aL܍W� WT)x��{�����C>��G���GPʻ9�νe���9�h�D9�wO��� LkƁqB<$%6����t�:b�I������E\�~sW��^U��ZGu=�lji��!�Uz^>u��U�H�����8yF��>����a\�����d�oy<�\���4�LSt�T=�:h�!7Q9B��i>g�Gq������P}�u���A+0%f�F ��
!�_8�Pi0�.?D��s�9��U/�V��M�s�:�s��9y��ےu�7��0��р�W!�V@3V��2j�h����0U�l��hgg^k�,˺%7v��Z��Z�YX����Y1�?���U"_W��Ns�Y��hr�	�(sPd0�`�A�%:aeP�;��9#��Q�y���4d5e��ng��=��3����<��"�(�Z,��J\P�^��'�I��������U�l�>�T����xK��i��"e:kT7<��e(��_#B(�\���9�i��e���<*�Ân��\WX������x��v��֍~ӥ']�l��v���1l�+���D���f���*F������|�+sT������G��ׯ�u�6� ruq�v:���J���ڌN��DEl;��>b� ,@i,1�I��eBeBab���]{�����)��P����[B}8�b�Ԋk�|هlT��{�ӇwT���
��F����Tb�C�:�s��[,�9h��xW��:� C����/�E���+0h㷗3�13u4Q�Υ4������Lk`�34e�.���@��� ?O�	�z����ef��v�ky���U-i�B.3Z�v3SA�p1�̆v͘.�YM�	n�������+���ϻsf�XIo����t}߲�P΁jl���ʻ��<K����{�2�����G{/7rt¥LPi��])�	p���f(�W�����ZE��-����͚v(������Ov]:��T%� J��*�9u���&�7��c��z��m �5A���i�s[�YHNEOm���R$i��PE�i\�+�[dRQj�و��R�.�b�C4���P�� gva9���g _���%)�^�)�,vM��b�"y����8��H��%��04���;��AR�u8��N�6x2kʉd�i`�)���Y�ƙ��/����^0O�z�6�d��?��0�:�ң?�h�׾M����kB��b�m��t�%#�f>s{TF��\��f�=�,T���
jr���T"�˻@�שs޵ӬRa��w
*�˘�s)X�]�nk�@WqL�,���0�%Fd�����d2�y��� �i�	���ಁ��̊̈(�ȁ�����~�5��|`|�Y�;�;oG̹�b�O�m�R$�s�)�z(�%k�s9-�'�	����^��Q�n�y8e��E-�*yY�q�O�]�M��P���5�t�x��PByՐbo;��֒�-DOC���֞��2���W�K�:�-@%ﭺSA�����Fy8牎=%���'��*F��9ۮ+e��#�ڧ��A�V<55wd�8�S���[�LЧ�]H�� ��ߟ^����"-$h�8\�Z= ɀ�܉�+]\�M�Λ/�;ȹ|{t%���^�;"�
,�Fu�8,q��ɹ״��V�{, ?>j��gqy�<)��e ���yb+]"g:4��[P�;�g�Z��k��m�ݥ^����?�%נ�Ӷpq��p���ީ��\b��<��"F��,�8�̓[6�w�jKn���y����g�lw�I �'�&��2�@��%:�������}#1kʴ���<ʆ��Ia�M.s(��B�S9(��s��Jo:�(W܉ߠLMy�[�|�����@��]��xٖx�;�#�Y�&Kw
�:��EN���q� ��&��b��E��a�
n3,h�v�=�4�re�I�@�I�m",T����`�#{ok���k:>Pi���0�S:eڭR�I_r�`��r�HD3�SA�|F�F�B�U�Y�ftffu�~TS��0�̈39(8£2"̠*{������{�㞞��k���&O�RX[L�98�`{j<d/KAn$'JuBY���W�B����0=��e��.EHi��ӕWY��Krvf^��N(k�Y��Y�+��ba�n���]F�ewܯr�X�ß%o�Hξ�j�K��.5�ˁ���p[�+�8�,6�غ.��ͻ���5�fq�uÙ��j�FY��s1zbU���{��)V�1�`<��&4�����k��օ�"3s�=zw��l$k�W̮@+u40^x3#��@�5�?3X�}���4�^���b�5��dm�Mۻ,�׫B�ْ��t}�Qjl�h�м�[r����M1nsLM�Ȯ�lS]\�q��8x�(��]�����e�5/���L�G��@ST:e�2Ae�6��Ď�Ž\��C�<#��y׉�e��T��+�P���CޡR� (�-n]����\������)���s�cN ]��oxR�7ʓ
�L&���)=�oG6�?%��뻁8�$X��+O��]<|��1^�9�>z-_���6�XXβ���p{����o��gzsD��V��E�3v�����t6�� QJU�����%٦9 ���ȸ�F��LX��{������H!��%�Y��ϸ��X~����@��S&�냠���&���3凌�-��� #�\P����H�dܜ��lxkN9�V,�|��u�]��f��s���)��UI�aQ�UfQY�@�	�Q�<����y����ߟ���xg}�l�LBq>��Υ��V���\H7�r�b��YRY5�/Q̹�ֶ�y�Նy�ü�mDߍ�E����*%ןm�S�C)��or��;gv��z	�^ƌC��"�6$�sw=4'� �
���(��8Cʈ�
�l��<`?=�.�<0��Mۭ<�c޸:�<�zqZ�O0�o���SLs����iP����%�>0�C��n33w5<ZG��s�$AxZq��f����\ِ�P�c���_��=�\|g���lwS�a�C�/���Be.eG]Q�X�>� Sy�)�$����L>��ś�F]�7�����n�����I�	��
�x�q8�z�3U�c:��W!!� ���p�\�5t,��\���f'L�m�G:B����4}�Mi�Pw��g	LQ2mS���;�dEh?���"����g�^�LB�)Y�J�jr/�>��qM��;j����)�t��ځ�x�T�71�b�B3L�*���+2�ߖ�Pԥ��)�aK���� � �O�
�9���A��2WM�y܁,S��#�Du9u�ރO���>lM�1�>��bN�i� oE�>nS���m+�.&u�5�!���k]4�C�i��B�9�V�.���T��vdo���Ŋ|�����%):��sn,~30bQ,�dV�L`&AeT&e&TL�������~�Os��+Yo�߈�ݙ,�UL��TSosl'�_��c<ב����;ϽR-�GEf�ۓ�:#׫Ʌ�ˁ�a���D��A� I��p����l�R�l�k���m�6�boK���'����[��`W�����5��e�\���=6��~�?:R�����p�.�>{����x.D^���e�,4����o�R�>p�gK&<���/�~����?�$�R]�w�B���GS�zc�
��.V�ĥ�!o�*e�Fdϙ���G���~�
3�d�;�lrP��AdGc �-
���.we
�_l?���N_�:8�����D��D\/	��e}�Z������W��7�c|jj ��wae�k��@+�,%���z���>�Gй�N��H��\�Q�s�v��mp��e�f�ZdhFӤ��ݓwF�F��'��|�b�MyČ��+6}�}!�8�fXc���zF��.��3���}n�z�R�]	߀L�gXE��ƄC��� 	�A�^�1�mֈ�{�H�H��S��U�S�Î���:��9�/Q�w!���.��sGrs0n�ݷ&wk>���K�=��ў���yV>iB1�Է*wʬ��Φ�W�!�S�5`.�ح.tKǫti��ٽ���N�u�;��W+?*�~XQI��E�D~�+� ��(L( ��30�f�l�^@�tWO5R�@�:���	a�I��沜��?!���\��.�گ���B��j�Z�x���6�]$�03i@P=��E��(<2l)S�&���wM1]�x{����O~G�����}��}�PĻ�D1%y������c{�Nu�";�I�P��~Hٰ��UEȦZ�*�	�N��7�s�7%K �.�G���|t��t�R�v���bq���D(/�ׄ���_�B�VGu�JΞ�8�!i��D���/���Z���x9 ���Er��A�:+ȵ��۵���ݑƒ��5wZŮ���Dz�!�������]�uЬ؞���
��o@k|y�ח&*�|�5�m�Dx�u<\��� �{�1��<��]���f��'���ȕ�,�N�qT�:� �b]�ڌ�m6n�����s-��T���)��jNx��⵹+Ai��I�Ʊ��n��xO�������ǳs���Y!�#lE�u��q��n/��ۼ<�Sn7f��2�M��UZ^��{P�5����0oZ&�ܤ.�����C  �ܩY��y�i6��v������Ǜ���b�e���$H�����t����w��7��5͊�5`o��w�ˤ`���{>�
Pwn�YָVi;��UJ��4;Or�<����zv�F��^�w7M���UH%���7�튤�1��3Q\#1j��:L��8�Q��s�,ۥ�]lOhu�PX�6w
�`��3�{7�NtJ]��hec�H�(s�uU��RVY�1�1��R���j�к���%�y"����ͤ��+�^�%G���r>��=T�D��=��m:�O ����[�j��O]�v��zX�.�mi~�r��&{�e6ٻ�D��C�h�7tfu��!��>QM��x����U+�Y��[K@؝m��iu��%��
�]�.S�Ym_BM��"9:�?]�P�㥥[:��d%])�����nR)�6�L�9�ڛ�������F��0�,����`'���%K�V�1���.�ݣe���!oD�=@�D=���ʓ36L�o�5rT$��O*�d�[f���m�;wf��Ӻ�}�fK /�S��d,x��;;!�¹.S��-�֌6sflAnv�@��|t�h�&�*ڧ���wL�0�,�7(�>m�3=MC�.�E�� �~��w�mt�C�)e�\�x�' ͹M����D�+M��][���XA��z�ݜ�"����n���熭�"Nh�BI�-5�D�B�	�*�
ة�U���KK���6� �)}��]��
�*)�P�Q�yʲ��,�@��BH��G�Kt���
Yp���Z�mkH��ؐ�t,"a�v�Z%ec��Z�9�R1��A>�}��78_�U�T����ot�ZDk[�:��V<���rWGo�1<i��4����N�_D�*�dS���)��/���HE?�K�sM�b��4�p}�bB3&�}X�ƅ�<�i5fD�8���[�E+��\9��A]y|q�1т�w�u�Ԃ:�JlGU=���:y�<������C�
L[���c'U��[��
�i�w:;�Q�l��.3���f֥C.��._oi	�#�¢�%�"P�j�!�p�,Y2�a����n���]ࢦ���X&#$��������n�;�;{9���|�4�V�ԯF$�
��M�G/�f��y$̬�.�X���:�/+�>�Źr�V�jt�-����w���7��}�VJ?a^R�����CG�k���/�r���vx�����r�(28���ڄJ����ٗ��j>�݅�ǐ�w�U_�69���X]�Xj�ɂ;�Z�P��]�.�آ���˳��m�=C��ow��z�o�49	�fQV\�`�lG��M�Gl6���ں�%/���R4�9A����l���Dˮ�=ȑ���fk����#��o؝Ǝm�nжl����q���V:wm��=�a�tr�5���;��|�q��8�>�/���s�P�"ѷ�Xl wj;O�T�e�1A���d���%��FB p���%
�LI�vS�I2��1$�c��I�,�4�� ��0�JH�@�D��R� 2�I��F�j@�gTq�M�\0B�1"�YLq(B~��؁~
#%>����z�:����~T��#�;#&�J�%��w��>����} iZ{̥��!�O`�iJ+�s����=1��3ǧ���T>c���Hđ�Mх�$��L������ǎ�}��&#��c�2
����"�2ih>H��P�E53�N�u��eh&
H��,������ʩw�J�#�2����$�������ވ_�!w�]`�SM$ICA�2S�1�zu���]ҏ���쇽eQ���eT%	����ACM/y�3������~���/�O�f�u۩J�L����*\�I�=<}~<x��4$IET|���!M�PSE$�ĔxfRW��@$KI5!@Y��U4���3��I"�!YD{f-���{�6��������4�
ǵ.S1�12�)����[5��j�V'Ɋosm���4AT�)0��8�q��/�A�����˺��䨿�UBeD&a@:��DLd@&EeN�g�s��ί�g�VYO�ʓ��\�W;3/�_���M���.[�0��]��;��^FV�m �����]F��ڻ�U=<�H�7�MB}�=�9�φD�����p��4E�P}3+��]yg�Nq��n�?�1Ar�{ˋw%r>N��!�[�q�db���NP�7������w*��O���l��a�B���8��x΢s����8E��=j֐��K-|0g����K�~��H6�O����j�S�����$�2��%rLZ[S��,�qZ>w&=��Q�[U~�Q}Y��WG�,�HO�;G���Fc�/'��L�cz$����c��Σ|�b�b�pD� ��zS��9�+av1iz�,Ȱ)���#b���B�v�o3u�غ6�LF�ka�nz�5��Y]a2����T�@�"��)�ȧ|��lh)67TM�!ڼ���*�KΥ��w���lQda��¢�b�o%�� �L�>�S���9˺\��f�'fesz]�
�eH�SNby��2�lN3{	�=��O@{i���l[��v����UƩ�μ�Rn�"�=�-jG��(�:,����uVr޹��Vj�أ�z���H+�����nt���Ry��w:��Y9wz������9¹Z�ǭ��Y��M�����i>0��kj
K�v��Ob��-���H9&^��7|���}����Gy�[�z��f�R�A��V;�PFa�f4��LM��gw���W���+��� p��(3
�ʉ�!�"�xx{�Vn�S�{�La{���q��/W\�z��"��lh�B�oE�%�r��<���-�Ď�Nmy�پ�_߱8fB�$�zs
����Sg?g��t�f��;��B�jXX|�UX�v�kM��7"�X����]'ցd�y��Mi�-���&�ԣ�[���[���Ϗ<����8���Qo��:O6�B�B�/��hC�=�Xa`��ڻ�02�O�${�ӤbE�a j�ni�v�Y韮���z]sQ���:K����w�rޔ�uشhV����l�z*;�״5�35m��1��[�e� U�0���t��4P+�%�~{���{�ȡ���Ǘ����z��a����}0[����XE~�"_U����Pg��t����<�� �������P���Zo���(�/��ytb�ۅ۵��he�-��>BN;]5i3��DzL�"a��6G��#�WtSJ���ǎ��p���o{}��I)Q���!&Z��8�q����dǍ邀Q�ʵ��j��S�(N�(-�i�@>}�O N3�KT@v���������T ��d@/�;c�|$��V�c�����;1�}��9Q���Ѽ�Z�=���q��4e S���n�^t:^�PF���woP��Ū��v���F���G�y�CnC�kR����b���U�Z���-Bؓ��2P̽t�33�w>|����Fa@�WT$�Q�e�@fTX�f�3�������ބ�|s#���|�	V!�\#)�8��	hհ<zq3�^��P����wp��r*p���o��Q����D9��2�d�z}�0�����%���CG�� 
�7W�7r�G�,s���N��r�Ij'(�`���7P�B0���uHկ��C����Ms[���6F�Coi]6f�1ۭ�K�T�x���R'�vd�TI�D̫II�R;�/xl������U}N����5�����N����,'� ���UM^[)�R��,(/tSۃj������Z���1�)x���wz՝�r ��k��I�L��D3e�IU���m�L�t�ڛzYO2|b)����I�e�
�ga��V;0kq�[�s�!�|�x�7/�iG7_0��{Wp�j��{6�<6�R�!ΓVb�pPn�ӾGb)�}��bL�z���\�\���\� P��=8pw@!ˤ���R:/m�[]h�6]��!���6�I�Kl��-U7���4�3�Jsq�����G2�A�	G7-�0�G�
���ٚ��h.�dn|����T�ޒ���UꌳǏmk�4��5��GhMޝk�sY�R\M��!�Fs�έNx{0e�����r�1�uuX�av2���E�{�˟ h�;�f��V*�ﲎ!ܚ��3T�4�w6�Lޖ-�R��"��D�`P�9�o�@|3��`X� �@�e�A��ŀ`��P̮��>~�k?��u8hg����Z_��@2*'����� �Sga�Y9�g��z��j�_��g��Qk�,>�-jyKll8�딵׆�"<��R3w�^`T�h`���6�S����y>���� HL��a#,#�=9�q0a�/�ZU����I�"sj���vO��\��it�5�A������{��"��-$s~L�`���s��\"�\��c���4!�����#���U�]�&�,nV�8�����òɅ�F�I�Ēsp
�XУ�XNZ1W���w�v��|���A�Emfν��n@D����3��vԖ<�C�t��9k%�� ���ڄv�;��i}]�3�B��r��yc����m��cK�ʠ��]��2�����|��C��XE��F�,�yvA@��L�`W8�Wڔ�v��P �A��=1�fO7P#J�k�Z�Z��t�!�mض|&�T<5�pܡ��N��t	�#���en�̤��!2<�K�]�7J�Y��b�� y�1H�Ԣ��1ƺ�\�d�f��I�b��V6@L�l�-���QˡE���g?s��K_Q>O�qI~�:��=�e�X��0�wS�c���<�>6t��_9i��;.mB�KnؚșGVL�/�[L��Q�HQ�&�.$A$�a�!D:���j˸�7����>�Ɯ�;�	;o,7]B�}�p��$����1(m^dS�D���p^�%īce7��X���{u�]��vde�g�D��00 L�̊L�e� ̳0=�>�tӶ�	��V�L��V0��	��z;����q%@�9��(�}&u�8�|�t�2/��R	E���1���� j�]�We{�Hí֦�dG�C��_V"!"|��/�Zg�����Y�9�[�E���/^)��*�9�^=.���@�w�B#�V��0��cU)�Um��/Y+�G���7R���%�m��Me���n8�,����"�ϣքSes�`���{�eg�'�"��s(�_��i:wʢ�_yC� ��oӠ_�.�|Q�+�!��|Z4��gI��G�j�U{���p1_��,��P���Q#���'ڗ2/vv�g="������Fu?c�U�٫_�3M�)�^���E+$�na�5#![��!��W4]���j�4�9"�M����L2T�g�޴�axW���-"���VР=A�]��4�?0�A���8<{E95�ϛ����C,���5��u��M�x*@��,��Tx�^y+�5k�3��'a��\���f
ާ71Bg#��������͡2i��0}���Q��(grt
�%�3��K�)J��x.y츬J�x~P�e#Y����N�[�y 9U�Oxy���㞼q������t�T{����mؙ�7Z\+��dxA	$�/�^(�N:t��;֖R^��/i���i;\Ŏo$of��uZ��q�7Bn����㏘ �[�,���+����2�³*̣1`̋3Um^�)Z���xZs���@�^tb���-�g �o�D.�[�w�RB�����k�]�8cr6�N�� ;�;�3$<�z��BJ�O*H~��R35\[hOŕyq�m�6/}��{��@�����Ҽ/^w�-������`TQO��3� �`s�s�E����dޮ=��Gs�<��|������>/r�^&s(;
��DH�ts��VAi�ïZ�G/3@�8�{Zu�"6d~w������h�[�9F �gˍ��/^����Qp����ۖ����� ��q�z��2��}��̝� EY�?:�6�:1���\��O�|�ݍ�&m��uA*9N��
�:Q1�hW[��`R�
\ NAee���.׏ָ���oJ`%���%��)���y�(V��
9��A���vwU��2Iva��Л�<sU�t�ކ�"�bvW�����b��%��8�?O[�B�K;��O���r�U��ֱ�`���û�����Q��e�9�y89�2�l+�	��I���*�7�����n"�{��&�����NV�����)s��>r������"j�^���E��)����&
�����M${xӊ�l�\C9��J������G����U�d�,��>IoJn�ʮ�V�u6�����r��3d��M�����U��6�{����ks���<������:�a�E�s%��?}�����	�	�&�Be<���� %���q��Se�	����&3�7�T%���l��y�U��47�L�Lq����*
���|Yb��o66T�Ը.��<B��KO��̲r��hx�f�j��nxt�V���7�R��nz9��j�GW��h����r���+���0����@��7�ߚz�	��v[�|y��K_�xSx�4�aBkՒy	hǀ�סh�R�R&)o�Ho�4n� )_�E�]c�����[��ʥ�\1ՕK8C��	9����]���~�dv�����x�����!��\U�<6�����y�g��强��J"�to�9�b�Ɂ�D3��TL4�hi�n��P�5?-d_��gw6b^l��4���Dڦ�X��e:u�;�&�z,�_��S�;�W�S�4ע23�yy�p�8�V�f�b	���U~xK���-�=�Ъ��N�R ��ݭ�*6v�0��7�k�����^��^w *�HޙL��e�x��h��aEE�ǅ�<���i��j��qH��\�@#�����ş�AXC�f}PA�?r��y&Lr`���x�B����8���\FYdJ���ݧg��%=#Q��^��\E�CWz�xn��	&��%��6f�c�j�	�-�����Gv�d�.�����;b�ѵF���n��Wk�I�������������7�x5�a}9�v�`,���0���P��Rd��P��q�0g�����u����*"L|U�;:"Dq�ltx��Ȇ.�:z����#���Qf�r�e��xL�{cr�>�^��N�Ų=?6�ZhNgW� �I3Qӥ�ozϱe��	a����7ꊾ7껷TX�~c�Bf�L�@3�&6���B&�y���5���=@D����}��%��{^��e�&O9�g��wݵX�
]�� ����R�t�7�D��8�,y��!��B;�~/~P�H9�oMb{t����9�T[_����ƭ��a5���s>7^v�ѭ���
�AG-��7�Tv6s�H��<�0ۮ��J^qK4.7��O'�,�V��RV���>� G�����xx��&��ۚF皁2� ����!������0��yg�{��Stc������7���"&��I���U���]��3�'rF_��V80���2!��`P�NzfW��îFD�c�����F!/�ͽ�`P�y��)�Q0\��)A�kh3<@���w�F���\=��ԑ~t�k�|J���<=}+��A4����<�"�-$�Xׇ3	�!&����X�L��dUZ|(�qjT������C�����*"��q^�x�}*`2c�ݢ
��bT�^��Ǧ���i�Ke�!eTR���&�]���Y�f���ip{�sw�REwʴKDЩ��\�7U�^tYnW�6����/wk]X6��w��D'.G��1C�rq�&Bd}���CI!�T՛t�ΟU����S�L:��:E8���E�2vD��Ζ/�ͯID�����C�+M�ʒ�*jϜ]��][��s摻}y+e�T`b�)��04��*��Ż�bY6�K*�m-��~�9ׄ��b͇W�WO��2�X4�'|k�3�-�vP�q���S����|�8aT-��n�\o��2���@SM=m��a�V�90w���D['�M4�R�\�h��&�:��x��^^�B��5HI�0f]zI�l�:E\�հƠ8�q.}�h�E R�2y�W����"]�NX���)�Ф�~|R���'�����q���ܠk)�dO]i=���<9�P�����>g<Ĺ�ʢ�=��Z���p��Hݘ\瀎�0�R����Z���D;+|	Y`�#���LQ����/����T���a��%<ځ y�,�Ѽ��˔Ɋ0Y���ֽю�oygR|Z��f�D��5��UP����!)o$C>�r�Q���� X��	���,m+7��W��}��,V�qY�y�����	Cm�&m����b����Cw����L�ۥ����,��g���U��'��_��_��ѣz���v]ӂ �C&���<�-X�9a��C.�] To�*u���y	����_�BK�>� 7WyfD��Nb�K�J�>��w:�ܬ��T��X2o �K�"ެ����I�7y��J�V�W����a0������0Ͳ�]�K�t.��@z3:�wE��Q �֏����$iW@��l�N���j}�x&n!e�,��/Ur0��%b^��n?E��.`��9����U��ߤ:e:�&�BC���9l��G 1���
S��<`Xi�U)��S:p+�]�WC�j}3�[[����qC�����n�$��x{j��XDˢ�%��K',�爂�!+���jWG�QZԷ��K�S]9����A�^ȑ
<4Rkl��c�X�')Y�-�g�s���`c�t��|NN�؟OU4��MGKt��>G�t�S�S�̱b�~_��2��e Q�L����V�v�������k�|�B��D�?b����is��W���F����;K���.ōV�A��-"��}T(�w6U�hz�1�|5�/LiІ�=v��d��r�.-��;�˩��7���}��b�"�e�M~$�}��h��vL|�k|�=�-�(8��i��/]e\�\Ȫ�$(�B���|ϴX�)�Y#�[���fk2b=��i�A�DPD�����z=�\��
����5�/A�2��zX �{���@�ī~WP��@�&᷃&�]P�8�&�ŃugZh�qfq�5`��l��ګi�"nGȡT�e
y1B�h�W�I�F��`Cp�������H�>�
y�d�u�v�nJ)u����tr�J�1�q��"/x�z��c���4V�h�t�)a���D:$.��u���YI��Im`p
9o�4�f]6U�Yh"1��O�l��n;Z)�:�ꎇ^�J��c/:���k�b\�.l}��K6t���wXq>�<p�N�j�� *-c�����ƞ4>��*�ׇ���X�M50`%�Z�I�����H�Nmn>޽����lc++̭��s��w(b�+��� �M���̞���ϰ9.��^=Rv
6�R�;2�}��pl�9��ɑ��[V{��h�e���[ �����z3�
n��D�b��u�V9l��we�0�)����3[w���u��`z�"�������#��TGP��T�1��mSi�=]8�n�D��XT��RT\�>Wޛ��G������9Y�@b�QT��e���5��'U�DqL�d�j������82�u�;��&8��J%:|ș��C�3M�պj7;ٳ2
G�����Ks$����\���C�vS$�MW��i��}t;$��]ͬ�o�X���嚹��조�oQ}�5f��(�4�6f����̒�0�o�邘��Kvmv=�B�Q���3;1	��ӧ�wkd��80$��
�aV��Q��F`�̅@O\}�`ӛ��\/$ "�^�K�ط�0l�C)�ze�ه��@ĕ�؋���p��7��ֹ�?r��_t���Ybj��xض�M�;/!��}{�Ms�QCm��ב��cI�v3i��]NۓB[�XQ��������X�em�tX�en�I��7Yo��.��L�3gmk�o4����z�S�ˏf1o�j֝yռ��LQ�0�Y+ܘ�jw&�F���@��Рa�([}#� �%��Лol�"�9�(�f�1+r��E�3[6>�ƹl:+,�P� R9���޺"Σ;i�8�f�f
Vb���cYy���Є��M,���[��p��u�X&�̤8"�᪰��zr�M��;S���R�[�ͫ��8�Xˏr�m��$�]�U�u�����=v㥐��sl��0��(�E	���N�����&d0�ǋԱ�ݮҲ.6.��O��uS�n;��s�dͼq���ۄ�#D	��ˉ6r��[4n����oaH,�\��X�}n���y��Y�PU�Q-��l���fN|8V�w��F�r7|������Gx�k��JǏ�w�Ϟ~:���b� L�h�r<Ϊ)�ʓ30�q���}u��M)L_�g�r: �^YJ_2'	>A�e�?=�x���jH���z��!���4�%EWs�D�{�A��<x��}u�ݨ�J�������o�9%=]��5T�DH�8믏�]}v,�**Z��6�h~�PU�=<x�x��߻��
�+�cT�QG��E,Tݖ%%WRe3�ǷǏ>��D�О����d�PaU=��5ADD��>?u��c�;�(�j*(���CQUQ@PV�Du��8�����Xݢ�����b
>a�UTU|�"�bZ����2z�
��*"Z�b�j#��i
"h���72�*�
!�:b�HԂj�B�e�Feɳ����M]m����cg0�wO�vBe�O.Mv��W����fˮ:I��-7"�*6���|�?�b�� ,�1�]A��F3�}�ߛ��﮴W�~����a}a��Tր��~��+��P��^�b�6ޮ�3mx�X㜑��{�޾|��q��|.��<ϩ�Ӏ��.�lL�o={K��D���iO0+��Uμ=��D��2̜�K�ʶ�,[��Rqi�%0� ŝ���ܽ�]�T*���⮛�mE���+H^�ȍ^��B�Ϥs_
�23�:�
�	<�����Y
6�\=Dr>��Y�)�e3��������
�z�BI��-�z/m��,ŧ�֏ ��O���t.�lO�/�l���Z�\�uD���8��
�U��g���I�0"����6��.x���62�ѕ���j3r��F��(j��fB�@��x���`_�߃���'܃��|�n9��o�߼_|8��g���1���B	o�l�����S����̲�h���,Y���]���㗛f�U0e�4ϏG�_��O�X8�F���0�[�ؿwsg������\$��ݲ��=\ڀʑ�7��޺DA�ւ{�	�p��U��8C�R��W�&y�I�lS+2��Z)L>��fhc;������������o��h�&�C�s��ԖI��(Nɀ���g�甧%�Ҥ�{t���^�u+u|���;W��vҿ�m�swfCUv�����c�'G�ǘ��a�a����鞱�Ͼ���u�V ���HN4Pw�&�9"q�܏��LeBxr��	J�2E�Q��Qc�&x�t(ԟ��t��1̏K-��j�X�z��z�7
��aTݙ)�{Q3JoKV^�S��(�l;�>���H��<�B�TPuخF8��w v���sa�����ι�j�)��,�aAtճ1�l��!uMX�OS�1#Ҽy�2���R-�q�Yk\1HW��P��Z��9Y��=�
�m���3�`��U\v�o��j�1���� і��c�q�㋵nűyΎ���1Q|11���+����Lu�^�q���&�Zh��P�*�\��H�%��vu�h��ϯ[�ڨ]O]�y�,�oH��d�(�e��F��Q��^Z��#\h=�Xr�Kw~9�=wQ�����/�4�W�Wԥ�Js�禡}Ҙ�>�s�e��b�����&FU�&�:8
e�b��{3 ��y���!���)�,�l<�F���o��d���zi3�ƥ�Z���P/�:�w�������������N|o�-O 2D8�mo�C�Y���[Sw����f�7��F�YE�ɪ�hĵ�],m%�[،�"�=}c\pg	��Z��8<.��ˬ����q�;�e{[�=�t�7�$��r�`�F�
�>�y�������2��)����	�V���N0*vW>�;[;�,��Mw[N�q^F��#��=�ڹ���ݩf �ɬ8Ok�m�&č�d��ї��b`����3:�C�l�f`�g�gWL�X��W��t׏Bٲ���_��
k�+N����	�u�e����r�,���P������]����ɵF3�Mzs;�����p~��8�XP�toJ&�8E�j��*ۍ��!ُ-r��[�����q$7���	���(6�A�d���X��!+� .R5BXIF劭N`��"&-�l���\�T��ٍ]x�ܝ�^�<���=d��ŷ��=�H��J��:~`�o���{�Lw;���I�'����n��g¯�Iݡ�uTQ�;�5ChʆOh�f�E��UeC
���ؘ�oV��ʑ��P�<7���m,2�∸pu�\a�+-�bY6_�ʦ�m
�E79������9�P����!{5 ���<�G���n7@�x�Zx�-�I�8�/K�te8�����{C��*+}ff=��&���T�0����7Ϻ��5ܵ4k
��fUu8e��1�h�0���V3o&��Zy\�y�kCT�z�@�.�L��,�O��f�Nz'��OFF�l'y�.�^�mq��{�����*�zb�q)�ؖ>��c�M�U��>�F8k���P�TŪ�<�y���Ur�A�@�Tif�A�Պ�ц�^5�t����=�Ϥ�g,QJ�x��9�W�5h6�Rƽ�w�*�y랖8ҝ��ܡ2�]�ST%Z�ݩ����\)of�==FR̵
LM^������e3�tg��@�R-���/pko�xni���E�#�`�Rw�=
:5��GlP��ȳ}5{�Ds��~~��sy|��:֩�9�F�Țy�KWO�y�ݹ2�0#%��3�"�\r9\3@f� ���y���g� �	���nڠ�G���V��qϤV�F��a����Ǉ>���b߯;6M'>ne6mK"
D��W���Cܥ�3�'1���߆Κٽ��ƕ������Z��׺�F���k�h�	��,�{�Ν���,V��:ޅOs��� �md��
���+��� �+�Pt#�^D�`�a|ß�bc�Q�t���{Ш�g�x/ӹ�ܜ
N�=Gxc���[x�{9�|�|���3�y<��W)�	gJq�/���K�J���Sy��X@xz;ʅ��R%E����/ȵ}�🾩F߾���S(�ͼ�sQ6��|[ͽC�4���M�hMyTU�Y�v��s�fb���� ǌk��qZ�w;!E)��������#������|�J�O $E޲�`��:�f��|\)mb/��/7-T��y���-+37LQM�^}�X'��Ո�Rȿ��JD�(i����^�旇���|��$:�����qW/}��K��{�<stὬI�[s�m���p�ً�DF�-Ś3��Y��Ө����ic���烗\�����C��7��Ƿ�7�ؚ�d�{w�6�!�EyTD(.�&J�Q[ɡ>���ޢ��*l��0%�cR��Î�Gs:2����|�ؤ�޼[#h��qv�i�M[��%賶Kцu�A#����toT����v�C7/l���#z!7�f��R1�ݣ}B�H˫���zV)ZB0I���W8`�w�^���ǥ�sB�� \�h�b�Q�����1L���T@7���co𞗑�9�)�s�(c��fJ��\�H^�C����LO��'O4)=�aspO�X�ɐ�`�3�豷�b�7j�l#	��lح�iծ�i�e��N�yj:�I�~;Q����kl�@dW�y�+K&��\q�k�V���=�~���<q���$�:J<�t�B|B}2S��{k�0{��+s"�r����;���j�r��[�UE=iݙ����tqע���ql3�c��<�D>��jj܉;J�~F���Sm��	���c�������1m�`�Y�5�˽��k�7����YޢO�J�\%�>9e��S�תx�i�V}="a������T1V�QE�������N*8��=�^l��gz�[I]u�C�r��:�GkE�X��p3����:���m۔X�O��^m��,�}}��1�)c��s��魫�ڵ֠wۭ�{ô�(�w��ˎ%��̮u��������dC���Y0�˝�9����q-"v^�P�O�o
��ql˪y�����ı2=�#nڎ����� �NV��v��9��GE�	�r�Gb��0�������=�_|�^�D'���T���N�J$�;�A�x+����1C��8��?E����{�C�K�>?�ne�w�ߘ�{'gC;�j=���2�>2@]7Q�vs�y�D��+�ѡ#�7����3>2���ջ�L�/sK4ϠV��Ed&�n|&�7�2��r&�4�4[!_�.�u>��������!�.�&~�����2����1�S��*�g��8��ڑD���o�>B��P���E.	I��ڭ?�l�i���a5�)��2�\�QM�VV0�U���R�m�[E�E��Wu5/K�;�h��@q�QkBe]�3��j׏.#��2mkڎҲ��Uvl$��<7�����-� d�d��e�i~�o}6�􇑪W8����y�1Ǌ�}ˊ�S�(�V{|�vGtv-4��&�'d�stJ����N|'׽��d9t��oA0�p��EX,;b�捨�tj�B�V�������V�G� �ltwU���¢��%^0�;�<}{V�,E�nT��dF�*��X��HݼI�6z��>Q��Ե�n�/0K�[?e�e�twY�V����R��۹K�wB1�è+>�5�'���?RP��12D*1QP�BC$�9���~E��A�g��g,���zrh�|y!2~�7��*�EW'!D=n�׿'��-H1Я�TO�~?v�����;���a����j��R-H��;<ݎ'�s��Ǳ$ `@��\y>1 ��s.6z�m��յ����/%�CCk\gM5P�(vN���yډ�lZ���n�^���6�ulj�!2%0jlwM�����SM��"���`+~��ܾb���b��v�W���5\�n�׌��mM���X�u}���1a���,�+�t�k0MȘ�%���a����ш���F�9����W �@] \Yv�{�XZ&��Y�Vn���n��&%�P�2잡������W����Cj���@e�c��'�~��k^���1�K�Z}�cV�����hp�w�0/Tʸ�0�J��U�T�S���N#K�\Gy��1��m���>�� �V�v�S�j�i�y#��*�Tt�x���v.��]��v�YJ����ƞ���u�"f����M�"�= jy��[м��Y�dڕ̶O1F�fw��sջ�D��9�K�\밸�g|z8� eķ�}��2�\�Ǜ��b�m��
���eԽ�[�!�f���U��d�S�Un��a���|0)�P=�n��v���p��/��.����cPIٻ��bC�,�&fbh0��o�}�T�>�����s�7fO���!U�������xZ�Ι^�)��e�(7"j0[b�0ﴻ�)�ZK���}mY��7���cCCS?����%�Kr�/�3�;1�'�%��Z;�b�n��tNQ��a7j�ʶ�����_Ӟg�`��G��2~)�v�w�z��37�������-{dԵ�S����H��+7C(G�\�HN�{!P�w�37�l�{�iW>���1�"�s�7�F}��D;9�W��U�w��|Q��>��H�]1)ߴ��9�ȩFr;���8uL�B��Z���0�P*:5*՚����r��E9�6�4#9����UD9��N+�S�>�~�ԙ!�����A���9~]�J��Y�G�H�ײ�'Λ�s�K����=ᒽ���65�u�� X�z��'}�p	+�C���4 ���O#ѦEr�.2���e�Y�W:k�dc_��s�Uz8/���^.�E�1}�W����K��TP�Zh�&�\\�#{���fP���"}�
����8�0�B>TkEz�$��y��j����-�L�1-L�ɐҢ�����ɺT3]8��ޗ�����{Tو����^Dg�j��)X�=gF������^�|������^Jq=�:1��jv����5���l���itr2�\=e�N3�5��X>�1,Hb[Ag������ub������%f�
�k�Dl�嚄���1�+�%r����x+�?������n(%���GG�������ɢQ6,�õx�<�o��=�R���C�8�.�#w8k��O��8GMId����l�ɝ�$�&�2+�k���R7��,x[����u����~���W��2�̮sP����=!ݭ��@�������Ġ@�~�V{GW�u<������3vi�D�J�h*7iިV3��"���Fˣ����	����邂��5d��B����jl奐��˞��'�Kho�w!v/.QaV�����8������2bKm���z@�Q.>�OF1l�R$oI�ہ#CȬB��+����\�>�߶"�Z�e��J*��°�ڍe��#~�4P�6�ٞO~�f�7�Q�]v0.��:ؙ�3��U�-��-�T�Y�T`��':b�eqU�@P3��G�O��p�^��&�ҨYY.����=�>|� uMV�h|w��R^E�"��p���&�"3MVd���Ȱn��zڷ�g)�^Y�����44 K��H��+t��ݘ{x�f��F�+T8�0��"��uy����G�Й|rT������;�r���T�<w^.�g�Ől3ai��2��oq]��p8�o Ƒ��gX���o?7Xnl&͢�ΰ��)��by��tt��ߟ5CIf�:�oPI{����0�ҷ3�W^%�o�D��a5�����-ʛ����x#Z�Ta��Ma�8?�.,���|�=CÒo%�j�Y�2�w�%��OL��p��4�ϊb!��iGE��f�&����0x�ސ�9����{�o����$Vr%��r׫�4ɦcK��yĖ~03��q�����R��{o���v�۾�$L.]�G�s�D~XD]�=:��zWἰn��j%�;% ?��r���e�I�r�n��_Pwls�c'c<������m�tf�����\]+�11�Ӊ���o��͊#O�4W)�:�	'V�	��S�4��1��=,��e96�3�����Ϊ�fI�o���$_kˠ������)��<`�[����7�}}vC�,A5��l��zF	��q!7�'�֐�m�ľ{wƐR�Mts?x����aRwaay߾�r��E�݁Y-.<�v�7�ʭ׃׭Ӎ풬طŕ�� x ��a<e'D{�����Vuc1��P=vZ�.���0G�U��	�*�e�ams��L��=�������mC�xԃ������\�w+_�޼2�k:ja��p�e��6U]f�SE.D�ņ�Ngp�+�t�$��&29���/���>E�,^�f�v�1�xA6!���[���@�:�=��0�]/�,��yݷN���)�'2q�cb�֣�=w�i��+�vcg��6�;�k���֕����(Zy\��AvKۉ+Y09J�L�ͅ���V�Ⱥ-,T�B�kK��btK���S�%u,������Y�L���L|�y2����vt��j�-m���3Z2���@�5�,I!<�Qb����m^̅�l�iTq����b�@���c*��z��Mf�@;9ٴ��.:H�s���v���{�l���}d܅�:ZP�4�B]R	��P�C���.f�ae�5�I��|�O���r�;�ސ�k�}��z�2�pެ!	��r:j����V�q
�sw%�oBȝ!��#%��C�T�8���+o��8,�NNq�\�.xf�F�\p����I�Uq�T�9�܃k�+�VH�g�6Ru{uʅ�^듖��9��7��(f�ަ��l�0��Pg'��q��8�6��R���x�L���5i�`PZk�N-�|*�j�,r&)+t�'X�D(�W: m�=`Hb���I�����Հ�t�dK�z���n���TU�C�yEE�a�nK܈ފ�'��&���)/����xOw��y��bm��X�m��V��c����8-}�:��f���v��DV�_�EF����aZ���G��r����bDz-8�sm���m8���N��3�=֯����Hha袝a^@�5�`7��h����O�;�&�f4/UW�[�o��J�7gX�Ƽ��M��\�-j�ō��u�T% ���la��ܜ��Ƭ��oA����h`*Ip`��^#9�:���B"򢳼�dfϮ��<��5b��5L�L��e�ك;"�裖�]���.��YV�uB�N��^H��5"#hk�R��N��/�۽r����n}C��������ۦ�R������e]KN�UʐnO�P"�Mq��N�we����mV��#�nj<Ǔ�	 ����B��e)I���9����g@rgi��y�ugQVֹ�PX��A�ɜ��U�&~}�M1�G�Ѫ�'q1F��F4�p�)�1��>s�Gn����E%����]��n��,,��-f7�ͨ��v���u���]�B�\@�u^��fɪq����Hq�kw��-f^���b��݉�ˮ{�m3�\m�_4�N�9{�e�i�M1�G�*4Y��@ӊ0�J$� ��2�6ɓ"�B]?�@�$��iDBseԐ\�`��j�
7m���F2(�	`��2F�I�ф(�%1;03.���Ƚ�������J�ƚ��Q�fa�ՙ�L��_�����u��2����2���r�"��(*���dUue�'�>>�x��E��Vf4^�3]fQL�MYd�MY8�ۯ����A54T�¨�&�**�((��&��"<޻��g�O>�x���2�Ea9Dc�U!U�QnaSs���0�
g�>�^>�a��A3
f<���2�7��
/��M$�<|x�x�^�Ĕ��Su��QTU�Eng0��(�h'�Ǐ��>ﱅ�a��Uu��n&QA�T�Fa��AD3�ۯ����Q��q�z0������j(�+�:n��
�)��l���rji���d��u�]Yo~u�E�P5uNߔx|P�V4[u����^M�m����n庲��5��:���`n�K��5z8̪����E:���e�Xɀ�����#���Rw	9oд�ntАdX��p�f���x���-�t�_�%x�Tw��lmPb���d�*�\��)��5»������T7�1�S�W$]�C�yHg��Pwx�d-�$Mw��y,!0���M���h��$Ӿ�ּ=4؁ɶ�&m�\�O�|�%O�"u\h��,�M�775d�5�2��A�1�"��}m*8�J��zE��x���~h.��bzV������]�$��oh�Mk�s�����b,���ϔF�!��R�)>Գ�hN�n�`?#�s�.�T����׌
X�T�DF�t�1�2'|�k��
�aE/�b}
�q���j��/k��B-F�^�{��w�׻�`��?�بE>^41�@�I2�����=	����f|�8L�F��ҭ������r%�5�5��!�0�I��(jS��-�,}�T=�j+8�[p���ʗ}��6��hw���*C:ݙ.�քm:D۞���8�^Tm��o�0V;&��ʛXzXĽ��1��:���Fe���t�z1N�;a�r-�ʁȸG�Yr;���f�kĒ�~ݭ��47O{N2&싴�׎��V�=�bg�"9�e��UlDl�*��"p�]��G�"ܥ���K��ҕnܼMl}V�ӫ�^\���P�+�-6ܡ��
N�N �ŗ[�u¹����ߨ��E�$1A2Vި3�'ቚ7�j�[>5�cZ�[��ʘ���r��	a%�Hx�P�ډ6�Bٌ�6�s�9Ͳ�xyn+�x��C�e���z�k���|����n�-$���BQ[;�6��D	�^\���v�.%�%A��eu�|�y���uW����ΩE��y颮������N�؀-6�Z�uD�8�N ˡ�S`�~��y1j�ɵ�j-֘EvV��Ȋ��]� ^�r�5��D+�^\��t(o2j[��[ȱNnoTu��]L_��T�\@�����*s�۽yJH��d|�h�s����]��u��D�o^hQ:�HV�>�9�j:�G�k�*amoe,�a�C��K�;���
��uř� �x�ܬ�^�K�Q��jC6q�l�9�I����X�07Mȶ�q}��+yS
L��ȃ��k맭N|(��N�"V�a�1ڽ~N܌_LkbF�n$mlY��꡺�����)܈|aM>�`�O�_����Y"K�quѼ��˔ɬ�$���=�+س�Yޫg�HrL<x�~rV]���u�2+��x����W>Zk/��B�Q�G;twL��<���©D�=vy��H����;�S�;yk/J�@C��pAB���rs�s"��C����gFe��T���z+��q�$
d�;`$��Ć8�2!�^u�w���?O��hy?O3�4���?����/���׾��Vt��M�X|*.���t(���{v�{Ѧ+�e46�3�[.�K�u�_/ag/�vy��d��5I5j�W�Pve�6��D�N2��k=�MV���W�A��6�Vy#��G�/��L��7�
��	�����23�kH}9S�oAǮ0Y�ez:h�/"#�=�ͦ|�]_{�|�X�	|���]�YgK�E@���u���ED/2���e��KP��r� ��+�J�S���Jk��;F��������lOL" ��T.K��Ig&%n��I���kG�W9!	q#��o�>�4��?_�5�����*����/~=�ja��맔P����<��(H����8s\5l�)\�����+�q���6�}����6��)#�R]�}Þ&������W0�v�0�h%t+,j�a��#.���d�����~?2Շ� �o��7�X^��cߘ�lO65��s����dg��v�S��Df*=�i��1�4�V�>��4B�)��`m��έ�3wO,�,T�B0���.MjG�f�K
<y/ς;�.�WHƔ�1�=Zo��g!����JwV<'��r!6Y�'-��ǼEϱ�39��ކ�<���>��}�ۭ�������,S:LAb�]�[݇�9�:�B-%�b�qA��Sb�̫~���e�B]�9���E\�}�<��$�l�U�׽�f��&��|���~�60�z�<�Ɋe��
�ui�
��l�Y��6�Y��|	�N�c�۫���<��F5#~�`"}*�ڨ��@Y��^�ǎ�r��ҥ�"��N���Z֑��@�X�(憘��}��V�%ۡ�n/��с��w�]����p����,��/6�0���'t\�@,�������q��C�pf�]6��)MQ�i�0�q׫�0�^��WB�N����qgzaP���*�ޏ�x�k�Q�|�2͠�C ��ݱ«2����.��jz4��4�eԼ�|�o_��C,���� ��=H5CF�vg>�k��v�N4��7".�r��F�p��.�h��kdTI�@KB��e������-����#����e��4�Z�]�~Y>V��1f�	�)gG�8��##<��G�����d�&���K�a�,���[����A���3 
��m�*��NU����;��壢�����)�0ԅ������{�V��a�F۳w?m�8����$���*q�]I<�[����@�r��Y���0w�3?����ol]�n��7,��OޱUWwb��8'��\ې�x#��h�2��r5�A&滆C�q��gqU�4�8�n[�U�y�����o>$�$�	�`�?F��D::�����:/�妘�񏳄�L�v�Y�^�������N�7��TP�b陋��>htkTHr|Dk�*D��x�6��9a�V)�őŻW�U��Z��������ފt�@��Db$zj���?����,).�9~Y0^k{F�K��!z��P*}�<�sEx�kĭ�z��Vܼ<�ӽ�n�C�qƯ���>��2�0����g�D	z�R��Y�d��Qm�*�p4�<>q��Ş�v5���G�@�ٺ&�L?5u��p`k�`��&K�5M�%>^wt�xnG��:"U�+�\�9����&��t��1=/&��g���c��/O.u�1�ygrvkPE�q�ʒ�~�G�eE���y95�iA`7��Bㅤ�9]~.kt�Rz}���;eF��b����pnO��)>�OͩA��^��+�+e��~�f<�G�Y�_�&z��eo"F��5�:�%�z�@���dA*t�~�scq֨ƾ{/��#�v�y[��s�R��m�!=	.=��T�>̛jj���X�:��[NGA��*F,�Og�������Tܵ��6v�%��/�X�P�VP��z/��;|/c�CE.6%
f��ĝ�1�j�D�y����4��֛F�=�X�YcpMQ��9�ݝ������HƷ�����.�d����Z)X����]f9��4�3ws�����ޥ}���G�ag�G�?yTS�ƄP��J5y��ߏk�j��K�N3V�����r����](ezjD�A���0��r�Vдߕ������exp����Fy��Z�r�~��l6A�z2���	�DDo��^�[�l4�x��d�h�p]M�ù����[Z|��z����K�_��s�'��X\�f���v��f-�&/�~�Oq��k�qp,,@@���0(cH�B�Q�H�yt�˕m��*|�����'����1��Gx���>*�ѽ��,����H��VE��R���~7/����wh0ff0��g|��b�v�y��J�?�v�e�0��-O5�S6�`	��;�?������ڮߍE�#�qɶ����(7�����4TUR@��*l���FZ��d���X�i{x�˯��#�ksZ	eGo��*��m39�8�p��%r�}4Z�X�^�����.��'Yї�rw�x�&)-��̛qT;�
7��=���}袠�u0F�D�3���g󅞘����SʞPf�;�y6;l�k��(�@d˗��އg��bߵ���]�޺�Y7+ y�ê>g�=#]�T�x=���L����f*���_F3���K*Jڎ�\ڼ.o���W��ͽ�s��2��ɡ�I�0h���:����0FלO<�.%P_P���m�*�kr��| �}��|aQ���Q���8�y֥�b�O����(�mf��p1�wU������� 0�S	���&���7��M����'>K��c�j�����]"G�N7�v�$bѩ�ڳ�Hk5$лD��י�;V��$ڲ<O����*��޷�y9:��Z��q�6+p�C�T'�����\���,3s����>O�_�.o�<�A����xD���x�}2�R�U+����M�)Fk�/[���Z^%��-��Ϸ�ok�-ِ��<`��-a�ߝGX,?��#���R��
z��eܽ��qN:��0�.2�=B�_�t=U����"�Lyt��[�D�$U����y���ȿ�hm8�	dO��J��!��
ރoC�r�SièBh��6<��3$�u=o��:�!t�� <�v�PSפ:c \3YsC#�/�m��y\Z!ý�Y)�ӒL䶬�C�gh]���GAP�b��e8����Kt�ϭU�ɦ]Vj�I�^��&��������C}c
�˖��Yx�V+���H:�N�v��)r�j�:L3�<`��sSgR
GOV�6��WBX���n%�}��p�3�<k5G!8�g&�S�x�=������Xg6��."�=�v���C���}�#v-�F��5x�)Rb�c.&A�����Jd;H�%�r�z����*�Bd�Ω	�f!3�]�s��D����E].Y��p��E[u/���d|�8S�Z��kV��LʸȖ��p�~��o�|Ħ���R�7���@��v�r�|�S�"w�#��z�����&ԪD�U�)�bɈye��*�A[ɶ�Z~�w�����Q[�Kje�\�]p`k�j`(^�c�gb����ENc�[��4�˷%������U�5�%K{e�:��i�J��[�脟	O�[b��e���חM=c�}>�tq��yy!F<��P�=��~�G�B����`���rz$�\�+�#4s4t,S8�0�f��,�W��f`�0��o�Sd94v-�Zڦ�5�2<a0W�)Q���N����K��l�)����	N�R� hi׭P� zJst!��6�ʆ���e[9�-vWws[�F��:N$q�ZÉ���Ƒ�_D�4�X��:�8HJ��;����5��oӖVk�;���Ty@k�Ż��r?�qh�����:��� �~�`�}I[9��׬��T�P_KJH��̺�㣼:�P|1v��V�b�W9b}r�gj]\t, ���3(�A2p��U$۶J*5���^T�uv�K�6u�RC��?�n��,kM9�s)�V�Ɩ�7����h�w��Tj5���Xj�Ƈ�2�0�%)q��1n(2I�jA1,@�+���\2`[���� ��F��Lŧ�/����-�8�Y�FE�����-��9�6���/[{�tW0k������8^���G��4�K~��y�N�l��<�$��� ���ݗӛ�D���*��������a�@}��D@���WE�iwm5X�����Z���c�LFji��AuAJ59X�^=�L��*p��n�r���^�J���&�t�U�A��L���_Z� ��"E�\�5�
�Aр�jL�a����c8���e�o4�k)����.�f!�ْ��~N�� �$d���>F���+i����;ׄkc�\_vX��vy�S}��pˀ�~� Bf%�p"당K��(�M�sf����V=�֑>[r�����YGEߒ�]:R�̕� C[�2D5@09M=׫���
m�8����қ`�}W��x�5uc����3$��~͹��U3��R�P�F��\��A�r���ުL�y�m�x��s�]��Y����t\	m�7\����x�IK:����2��b���v@x�}63=I�U�K�ɝ>3�u��.�� ��nW�op5�sV>w,J��v���TWE�� =�%Q��3-�I��{��m9���zZ��gt���Ãɴ0�Φ��4�w
[ӸN�����tY�������~wa�?䙘a�Ƙ�G���9�e[2���tR{a~:n�9�
i�|�m��S\�aM:�m%G��g��M�ިj݅
$\M��1W�P�^��>�4�������yO��*9��R���)@GԄmoP�)��ϟ�|!bg�k��T��;6=��)O7�e�B(�\�;�-c-�$�Y���;����q�ջ�9u�q�&-r�G3������d���`c��
~nY�S�����~7�D����3YOC@�޵0p���e��|tR��:Q��?�P��]?���j3���\�$:xLR�5%�ͼ%�ޢ�qe�l9w+����Y�V�X������?Q�;/�s&��A��g����R�\��l�r�MhFӀ�Ǉ0X;b00H&��5�b�8�5v�F�!�v��>���^�['�I�H�_�H4��W�m5�a2t|��Y*�����m��߉F6�~�S�|%���ٳ�����а���-#��6\1�t���i����r"�]v5*�Zм�X��8�LL[����^���g�0��R�-�V�f� 0��༪�Et����s��3��B�`�(鵝5j�wA���/��΀����z��O�3v��Q�5���8���&�2�{Q�v;b{�J�.�sK=LK����.�OeiX�ͺ�0���);] ��=�@chq�$ןq��oW[<�뼾j�*���rW�<�Ŕ�p��4!�+4��m�e��z�SJO�n�`ʈ�T�:y�K��̜�R�'+VI�+)m�MKJ-��w,Qu���iـ\����=X�y�z�j���4�/3���X���Wb�A,R}��6Z��E�y�硴����}[�E��S��0�|�����tyҤ�o�8c�Ҋ�}iI�:�b���Z����C�0#������5J[�J�M�N_;��xf�2�wN��;�N���ӉVN;��:��\��ΰ0��<��M쫣�LK5 ������iu���NyGt�!Ɉ�ɕ��:��A�����.���`ILS�j�=���m��zvؓn����4	�k�SȔ�n� ���7lзA���yb[�\�&t<���K������4.������h����vw�m#�;���F-y:���{y=SML[�`��b��O*��x��������t�A֣|�y��o0��-��X`���&�:�U�w�����p9����w��z�5�B��2sώ��/E�ELn`�ٷ0c�/�SB��[Qi)5���K���f�C�T>`���C؄=N��E�����U<��H=�%�����!w(L�� �w��]�w�Y�'��iOr�Cӊ�2�H��9[ x��������I��<MX���j���_n8�=��~�z���P]7�_Y��8K5��,����k�GY�qw/���/UB֡�.�}�]��3��`"t%dA����4���P$-Ryd,��e%�Y8��(�Yս�@VwN�b��7�1���p�E�:N�q�m-�;6��1�%-x9ŷϩe�xe�n���:
�(�L�t���������	L �2�>y�#U�����9��ÿ�&(-��h��t���29)����[��tt��[��J/'0'E����j���9���l��W�K��Q�
�<���]&�U�� n�(;T��#9�[���Ƃ�)�z��Ǥ���O�s:q�<9�^���#��Z���9�m`pI�8��%]_nP�'�j�_; v^�X�+d{S$'/�κ��+��ǭW~(m-Ğ���Cm��e�����8��q@�����u�n�ɤm���c]c�p�U�P�s�`��3#��Ěw�y�z���v���㜎���<?m9�ϒK��FL�Y(�ԗ6���)}-l�i��5��KXr�^eA�v��5�8��v�ơ�u���WwC�qY���QQ1.�zȏ�eEx�TQY�A1�9Q%5S==�?_��wb*(�ȣ�d�^�E�TFf`�As�}��o�^?46����f8U�i��E1UŖݔD�3�On�뮆�ɕ�����
(��.fS�a-�(:��2��{{{x���]����
������(��	'^�u�]}6�+�$�h����NE�UiTQC�E���믮�l�Gy�1]�N���JD�M[`�������~�x�u<����B�`Ș��$�z�i��h��e�8��뮾��m4�U�SE5E/�d��a}��aU���i��:��h�)b=�ɠ�=T(�,�R��dJ5�}�]�v����}Y/2�u�©�������7��;�κ�{���13131�c���Sַ��r?Y�j6�iixu^+%�!���0:=-Y�$oG�ï��XX���!n{u~�_���{�����J�[�'��%��I���u8��T�f��GMs���.{ü�C� �M2n7٩e
�uVC�PaK�]�X܉�.)8L�kQ���T���^c&-m�_�����-��b����V�� cڭݎ�G��5��%���ie��A�`��U����5��(Z��� ��*r���?��ߥ哇�M<�P���d����>�.!ñ��<�m�Mk�&b�ӆ��9o�߶L�~��ŎjXr�mr:*���繅(C 0���ћ��P�Ѕ@醤�1;��V��~��Nݜ��[��Vl����j�G�`3��>���q�cl��D�\���+��a#�y���GU^,~�m���X��}�����!���� =�E<�򇛼,5_JCI����+=���d�B{9���mR/�i4x#�U�&p8(k�^*rȻ=i���w��lZ����Y�v��_C�o#��0�v�Es�,]�7�̽�{.�S�miY;���|)�J� j��3����c~�<{�v��R[�.��ֺm��tt�a��d�2U�H�j{ۋ��j�+tJ�̾�M�^E@xQu�G�1,KHĆ %��z�=}���:���LI�Zm�k��fX9�L�S�d6�^كk`wf����ĥ�B��iWk�&�Og�&e�8]Kf�s����=r�j�������f����9&�'��B}D�
�;�y�}���b�����͎\"�yW�@\}��;���W@��l?��q����槇DT�],R�f_�y���j[%XGPx]�:,���TE��_��4w���^����ڙ�g/��1�M��z&3jG)�M:�Ls������c#�SB�BMJ��R�(�����}w��Y3r�.�wJ�Ú���Gz)!�J׋X�����USTa�	yƽ�hF�[�r���y򸶆ĽJk��U��񻮄���$��ú��D�CH2�	����$�g�ns'���7'oB3kqe!ω�d�.>��-��~Ŵ6���q��.����Ԝ���Ȭ�z�rXZ�Q��o�z���)�-�F�����*<�,�X����>�<}Z[�u4�^������h���j�:`;�d�'�h��yۢ
y�{Afzì�{s+bz������'M�50�����%�V��@z���::������i{-����ea"�mc)09!����Y�O�0�ة#n��s�W�{��跕f�bU�zdJ�n����΄��J����͗��U�W�v�mP�i2L�tS�!:�0�a� �s|X�ĳȱI���=�k��ìN��]�Ga�Y��6�[꡴*H֕��(F(gT\K�u�T�s��Mɐ�N)췋u��*����"`�uIcφ*Su�L���+�x�?�@�Ў���$<�hko?b��Jʹ)3��p"���\
��p��\��FHQh��)�֯��1�燲y-]ă��f��vra�_l@�F�6�3��4�4*�U��lbr��V���tI2�8*��N��ߴ�����˭��b�����{U��KU󷓌�OTc߬��&��A�����.�a�뗕����׾
�S�1�� 8Xkd5@x��$~j1�Bs_ƞX eA
����en�ZEM��zr%�-����'<�І�E>��*7�U��IVE9Tv۞�Fu�D�پμuѨ��xr���Z�Y ;{f}�T�0Rv���dy���5�m��OSw�=62�yO�ڪ�zt�>�&�M�-9����>���������hI��`���>�X�$��},;{�TN�߸�{��x�\Ǔ�����E�*M\�i�m�j�U��g����p�Ի��i�b*W���.�2 ���6��Ǵ�,��r�FtZ�ٕz��9�;���-��=%�DOP�cV�a���V�bx�]v%YfG7Ecr�ٗX->�w���P2�.`ƶ���Ym�/o�%�������C�,V�3�p�ųמ8�X��ymijy�K��O,Nyez�.�@M��(V=�Z�"�;Q�O��Z_vwn��Y��Tu�����w�=����%J�mN��Q�e�D�k�3eI�\�����I<�W�.�*<�&���4]�g*�9��fj�Xd�)����
�*�=XGj�6�ƀ�\���6��\�
O[8^C����P.�@L���6%�+���ja-D<�r6=������م8�nZg��F�G���n����^� f�����_�[zB3s��kH��%��7ʁ����Tsg�c��0����Ykî�Hu��n^z���P�q|�iZ�S����n�Jy�>�F����(�e�`m�Om�0ٵ��*F��ɬ���m�󉃎|�I�1�h~>��"GY"Mz�g�� (QeG4ڈ�K�(�qv��
:a��Ah�	�C�3a��m��?<�p�}�B)��QC�<�F����M�{=��r.�Q�Uq9�Z;�&v��.)�I"}�A���,���a��l�(���^�LS?Sf{�����ž*����Q�J���Bp��
�'����/%�n|rX�.^���6A {�"w���� ���Т�4�]��]�魧�|�%.��:;�t�N���T��������4�wǊ�X���1E�12dbň,F1r%�vg�w
��O��;ef����lCcf�XgB6�&l�v���a��J����?��|���._�-�����rz�&��ʯ�ͰY�7��'5�,��_A^���~��Ɛ�{��5�4�&[@�r2�lƸ��6xT)���j;�����[���v�`:�|b�a�8�$�h`��w�\6�j�X�_���o��'�KϠ1��$��m]O�g�ٰ�)"�R���R�G�9��X�)
�QV���G��Xm�>����#m�p:c���\��Z�v�Z�ۄG��;鄧� uD�}_璏�t#�,0A�7���2���e/m�Һ�rގO;'<k;�d��vH�k�N�4�Z��xKN�>��Fsp�	|N_�f�I�U��oS��%���ݎ�<I��	����'��>cGK8�T���[8�x���v���7���z�2�ˋ���)�b�L��v@�ZJ�1���q]*V��T&��M�T�Q4H�;�[���g���gW�ګ�|V��]�м��&���|�s�	}��3��-)�4���oz�n�T�X��2�ɰH�Jm��|�~$n9�2����)����+�Ԉ=��������w�ٖ:Fۊ�ߵn����rD�+��(��*<�{��s�n��ӝ.Rn'�Ku�_7՝��h��oe�J�e��E��P�[Pp:�����Ű0d���ȱ,X]�-ȉ�>~�~ϜV�{"<�U�^<�<guѝ����zj�L0~5t.;��UG8N�w!0��uH�Cp�ȳ��l�'�R!q�[���� ν߇�m9ʲ���% ��. +H�OzW7mF�5��x�[��<��״�6	�e�3��f�	Q匌^��.F*:}z)f�K�XʕȪ����ѿ-솫�C���M�hD���*�I��{����߁
�z1�ң"tС�S���=���f���y�Mx׵�B���б}]�L��5��<S�F��0 8[K%��ޫ���S>��"@���? G��~�x�4T�UՖ`s���O��qH���֠%�.�]-nM��������8�|���j�û#Y�=U�Fz����Z��S:s�0�w<ē�g��;=��gꦉ|=P�UP���p���2z�"٥+����ƚ�����G�^U�o�Nb�ڙ�ڑʊ~�ެު�;R�^�.�5��<�� �7�&>��plͻ�쩈sC#��&�g\�I��	C�6��1��f�f��]U�'WީQ�NX7���(��]�a������T��ܲQ[^DM
lS6�ree,£[��W��|��+Ȧ����We7ٳ�r���s9�V�<�r�{�(ò�bM�#e@XM���L� �O%�e���i-ŀ!ɁgSD%�N�z���'bJ���¥ꔊ�z"LSH��Cׯ����
����Չ�%J��پ��y8~���롕���+�1^q�yE����M�!}�j����T]��F;��k�	̾DM$r�Yh���/y>'�cH8����R}§ˉw��,A���c"e�<��N�5�b��8����e�ܸb��؜�Myj����ӓ�\��g8b�e��T��+7q�ۣ5���4���,������s�Om�f+j�t� ۊu���/�u[(���<v��]�����~|.a���R�	��A���SG�T�o]���s�P�1��aC�<�JDڎ.(j��d3�a`���"Ϭ��Ƣ��!�3(v1��#I�č�X�yQnܧ���
�S�� sf���-(�EF7iKL��p*�擝�_���w� �������9�]��,=�*L\T�*\m�����Ynd)��݉y�k��΁�#�N4���)����P�����?�>�{N�:��Ö��ҧ�\W�d��G�'��s�aC�i��Y��n�d��.+����ږ�y(;zd��G"�M���v��ٕ�����d8lb��b&�P���ռ9Y�2ӧZ�ei�1�|ΩkD��p_�)Q��R����Q`��nL�L�$g�r7�ľw����:d�RѮ7�Ζ�@��D��=�)�ryQ�>{��x�ܼ2�[�o/óFK���q��3�Jk�$��gܭ<�KJ*�[�X�8w� ���U擙Y[��ޫ�����.����������X����W'@�{X�KK�*=����)���9��z�j̀�K׭�0窀��^(���>��άN�����T'���cA��~�k1z�y�'�PV0���GI<h��T}}-tD��`&��
ǚ�K�
������G���\Ma�Y����B?y�D38�q��XB�o_��CI�\����Ô�)�ڵ�5��w0�'r#WF������̕&~�ESD� o��!">�
k[ �[8��w]�SWo��3��nL�;��S.|O-�YX�ȁK�r�H���l�(d�,5���r�Pn[�#��ɗ��)��v�4�n���\G�Ơ6({�0_��ԷϚcqW��`z7#����f�!M�ye��3�V��ü��wGZ�]=��z�;Ġ�bN����Q�9v��i5����C�ҩ]����Q�h.�ۗ$�j���)A��\�uN*ٴ�=$o�A;m��ܖB�o�=��ˆ�јެ=� �q�W`�$+駺�i�kVLh&2�l�3e������1��L��8,K'L�38��oݲx,��K�;�R�]��H�5���z�#"$qo*�r�̷���r���s��ʯtnt�i<(�g�?<j=ca^�<��!�ǫ�Hv�B����n`�@,n�u�m�-�t����q��O!�P��5�a�ϾN_��t�|�i���e�K���ӻ�y9dC����0��f�l+�S�ƍr ��ZށC���~�|s���|'_��y*h���\� ���b���I�~S`n�m)�F̳�ق�L��	U��<*R�7g��P.�����پޔ�`!#`��8�qHѯMm������^�7�<^$�!WZ��3�u>�r���L�4�v����%����d�B��Ty�G\A�3K�����A�2�W����·��BV`wsI�4^��S�H�dc�>-� v��X]2Yf��r�0Y��;%�	d4��{Ʌ��Q9МF(T�L=>�i�0�$j1�L�ɜA�˴�8u�/(%%#�Ǿp�m�>���9RW�W��yM+�w�^kl�����֕� �T����]��
m�^�Q��ۺܤ��ޑͳ�%����Gh�bW&��#�ccs���O�Q��A�M�1Φm�ʫ\ ")r����\�x��%��S�����<��� :�aی�`��*���i�ڦ������'i廯_|X���Ř�HN�{/�?
���f���{2j�ɶ�)�ݱ\��[EC�ш��Tj�C��i`�5ó�J�=Y ǵ�K��厽�/�`Kl�*�>f:��/!��8��t�����@! ��m�t�	i)�:#��^Κ,țp85'����tJ�����+`D����E��;pc�6�zf�se����6�:��_z�n|��ཀK��f�LqzO�t�n���Tt�D_&���a�!,�ۡ�=u���1�*=E�x�L�ewE��@�ۙ=�O�g]���#��ʝ�{�<������͜�����N�!��c`��ʄ_��s듖v0��&U�`%��ЖB���^S��ױ��|킸<���i��!N0�B�� �.���ݥ�OU\vދ�t�k�V����v�0h���'�^;<�e�_��p7������
��v�o���֭A�L���i�Ǥ�r�M�)����U�=��Kc��}���M���K����p�~ ޯ:&\����8v~���G��#u��>������| �����J���v�<MW2�PO��kr͍w�S�(Ai��u��"�oo�R���ܛ���5��|���QU�p,�n�B�#�V��\�M,h�����:/CҫU��v��c3l�E�͘9�S�	b�����s�I�����Iy�*�[�%�~��{)�rQ"��o�Q�'P}�-�Q���Cs��͝�&�� *������#].�W�d[�st����	@�8̰f�q�.5�i.�����7� �Lnttz�+���+!�0����t�L�����RU&��J�&�ר�<�l�:�MQ�=��3"�a�)w��l�n��,*W]b��Q� �W��V�cpyԐI�}��	Ѽ6E��Ց�-WL�=��C|�^%r�toa,���+'�� �֛��"�]�˳7�s�ns�����vcw4*��/����J�2W`7{�pf)]��c6���yS�Ҷ�^���� �V���b_MR��ɒ
KZ��=�!T���Z�oy�7��r�V�i/rm���k����lv7W[)��pܢ��;�֕Z�%�������uh�Ǻ���׮�	&du&f���0)_nQF�Z�V��7u`���g11^��M��Y�+���[DlP�vkf��ŗ�Ƅn�\��hnĭGI[:�@s3GMHԚ�F�aX+�v��]dnj�N
PgW���lY�n༩��'�)�_õX����t�<���`F��D�`9f�
�[J�5ͻ���,�쿩<2���9ho�W-I�_��kN�X�����/�c�i��}v�+l� [���v�I����3��b��^-v����N�Ŧ� �}����
}�w��鷐v�Z�i�m����@�
�;�vnch.���%��`�I�]5��ْvծ�zl<��-�j��_d��>��^S�O:�(��u�%d����d$!���G�=U�nbǃ��S/�N[2�Ɨd򮾋wc
���Ó��wh�YS���%�N1��ݳ���{NiYFQ躄<�m79�U$9��q�Wf���x6_Z�Cm�pL:u��l
>����u:�r�Q�om�h��N�9A��\�c���;�v���8g����XA�!��#�5�Ѻu0��U��0����ڥE-	g'˯rLb`;S�[�-��Í�T%�2�;�øM�$�Q;�y�k�]hMW:-���/:D��M~�9I�&��`!�m�~2)�G�]�:����нڝL?w[h�n(�&ZN�ֲ��v>۶�8շ��+qՊJ�~a�ȮWeGK��11�T/�S��A�*�J�&�6/�Y&��xȉ��V��)�4�؍�x�x��6��*7��Mq���e�kA�N��]��O\�]����g����o;rpn٨���lF�"j��Ru �R�
�D��J��QSPU0�N5��4
H�h�����r!Q�$?��b&���PK [�E[i�Q�\ �i��BE��?(�	�i���g�e����Ku�I�5����QITQE-fn9Ub��UA==?�����QAL�EE4�W��4P�T��MR�m�N=:뮺��!*��DGiMPS��c�;"��aU@AU�$���?<t6N��uIT$@U%$A�S hI��Ǐx鑰�A�TTPS5Q�LMD�RӲd�Ӯ��믱�5��H|�!z�h�9As�����PQ�aA8����M�>��5MRnORQOQ�-�VE-_Ŋ��$ɟ�Ǐx�l�P��z�)��7X�v4QSJ�s"�����Jg������u�6��f���?n�#�&�����{Hr���J��(j��ʞ_H:�"B�����Ơ���5�إ���_�I��&��e*����@����#PEΆ���v����\w�^��-ɈH��h�6&��ԝ���"$��\�,[t�`�
fA��y�V772�t���ı,�����>�4�Ċ4����|�9�1Z��.���y���z�94v+��-�xo[���<惪�(�;���1�]a���͘�璹it��}�Q)�l�B:0��xz>�W]��r���r���͍��Y����b��)]��5n�G�TL<��ّ>���r���M��c���3�/9p�����./�H��,`�P�*dKe.�وF-�`3k%��޳6c���񖈝���Wc��Y�*Y�o�C���P�/�xo4���[�H�C;���m�����f�ʄw!Ui���5�m�(���S��.n+*�`��VW{j���L]�P��.p���J:�z*��[n���ͼ��r�HM;���d�Z�Mf:��)=�`���3��ۘzux�\�=W�n@��r�p�M��ź��-��R�0�@Cq��'�'3J�[�/�3����C<�d�X�U�ڃW:� jq��7��6-��fE���������q�^VP���
xf8�)�w)�9�P�����61}a�j�<�Q�]N�\"G8j���pȕ�v�s��]�0='Yr�S�6��b�]6ĩ��4A�$ܻ�.�O{.U��;A@c���ar��W:�Ǫ�\�XQy�/�5���o9�p�O���b������Ub��S�>m!�!������/�k>�Q�J������E��
v��ނͭs�7K�NU.�v!��/ʡ�p���d��V�9���wV_�-x�X7Oien�	���/��{�L�h��R��8��'��&�>�\T�[����i$�n�T��$7�؋���T����f�/2 tq�y��#���kQ�z\_�LV���=��o���LB��,��2��fMOb)OXU��wޞ�� �2�m���[��a�z��GC��~�A���enok�8�e�]��I�j������tЄi ��i�;oC�uFR�d�%n����~k=��\�qs9�ݛ���=���va�帰���ё���e���DwT�U��J�{�+w�ܛ�W�⯬�_h���V��e�)�d��#Z��W�
����y����h�*�g�lPV�w򊵲(��h�5o�K#%��ⴄ��:�u��^����H�Ox[y�:«*��Z\�O������er�}���͎�	F���Wa4�\�i��m���6u*;p�MT-�id}�lr����x�T[�y��H�:�1hn�ќ�-ͭ�ݙmv�x��S��95������d���j������de�U�g�m)J�jrJ�4���2�ff����6oEN�;Fx>��J<*��V8�*�0��K��*���m��^��Q�����G��_uP+̷�E�4K�7����tR�ev�J��Ҥ�u;Q=�¦h{�;=׍1��R�(�'xz�7l�p�iT�ٵ'{��ʂ}��l�7͓51C�/����59ܰ�1������8dz�DBޡ1��ЪY�OR��va��{y��Vu(�,�&�S_�t�u��K0�#Ude�O~�3��A��>��:�]]]�]?=������~����)<�+���{�^�,��R/({�RZ'䤜�zZ��f�[��C�E�����ͽY�xEO�А��罆����^SaԺpğ�7�X�h�u(�=��ӱ`�]V����7.�Խ)�?��2�@֧��?�w}&D:�����U��.�\6�33�G����ۦh=Q��_�� ����֗�o}:��?a�Gz
~<�L��ݒJl��#�f�t�$���]D$)��\�~h-�Y1`	�;��l_n�&,�Y9�/v5Ĳ�M�ǨU�_y�Y��TM��cd����5*
>�lR��]��X��T2I��$�e����M�(�)g�/0�noӢn��s`�(�[2��F�c����U>�CNK󆶝8�_c���P	����.}��J0\*��B�~����X�,(ǥq���}
��ɽ�R�'���'=+�r�ɜ�n��FEe[�ީܤ��8c�כ`�[���@N�;B���J���2��x��]��<�Z�Mw4�d��]z����A��]��	e���x�X�g��}�EgH�����jQC�O�����G��g�jЅg1{~�7�z�&g��uUc8�1/��}�z��
ԢF�
�uʄ���ǆ�5?<;�*JG�3r����f.#N���:H��}�H���uE �Џ�}ޯ��H��7B��e����{$�X�x�u��jgK�s�N���
��!x�A,�:uZ���n&P�kUD&�˛������5���}��͚q�hg������)�ȃ=U.�sWRA�`b�I�ݒ�\�/{j��5�&�M)�����;����Χ����?.C��C�=��X�f��3����L~+����W����lk�P���B�n��N_�������M4Lx�f������Y]���ަuLˆw{���9+ٵ�{g"�c�6���Y�Zn�;��@��q��әk�c�d �a�]Ũ";��p0n�bN�^Je��l{O�S]mhX/���r3����m������dƪP�YÞ,��vE�2�`r��>���T [v9�m���qC�.�x;����R�0iba�7O�6���z#�=��u��-_��F�PY�ɮ��|��Z2��ZZS>ךʇ���eA�W_Nb���;�zϢq]]�Ym�+|7���F}��q�?��5�.�l�T��c����@������۞�f]��i�7�q��=C*v[��u�"�f��^�U�^�4�HJ\�t�0��cCP�tV_{Og���|�m�K�Y,�N�&�8�����6�\����`���u��vC�0��Q�w�%�ss���t�W��c�"��=�Z;�&cC˺��CFU�\�G6������{s�4$z��Us�V�)�b8�7vۥf���@������i�3gqS�D}�UU�c7�zC]�ڏ\��
΍��d�KESe��j���2L�[$v��F�ݝ���ec���i�M��5M�\ݴE�m�Sۺ7�m��!��2�gͱƏJ�ⷂ�w�W1��C�rV�S2b��]Fj�A.q�w4g�&�ǁ~��˳�J�\�=��UYS��Gse44Y�WP�=m��3��Z��^K<c��8�1�L��q炩GK��4�R!���	���D $Г��,n.5yjx��c��z�z	h{xyyFɆ�YI'{�J�����V���>�N[9.�z����3��%Q�Y]���J��`_���!��^��u��� / �zez+�k_��B��\�0�����LE������	�ق�`?o6�	O�l�ב�&q�?�"����C�u�6������
G��Cu�	m�|~�T~��t$r|ꇈUd�݃ �������O�>Fe�r��s�؝�{��Ŕ&B|��k�슣5�h��sb`�{�O���/���`��g�	�Z�AG�:�Ȯ`Ƌ��جs�e�͉�-����pާn��9����A�zٱ5�b��Hg%�������<P�.3s���^*��*�X��i3�(Lj/2�2V�2i�3I��j�ՙ���Қ�fOj��qTե��*���O���Onv�㼢_�Λ�f�C�]�C@�y�vb}ă}""+�wz��� ����ZۥۄB�;q�oa�B����;�}P,�>�:���5�QL��h��ǟ��g}��F�sXM��z~'��	u�~�fbo��=]�Z�WE����'H�����	aP�Z��\���rU��)�07��O��.�J� �y�U�z�L2v	��|pg����3��a����u���3yd�\��h��C�i��mK������o.�]����u�Ꙋ�܃��8�O wWO��٦Z�7i̭�2��`�P'�����\�0�#z�1���m��?s߉g���Xbx	z�6)B[��n��P�R�빷����abW]�v��+������s�G��dh�CԮ�^���2�VA^5㎧l�Y��4R��%���qg����B�����pBE��ۚ��0��$��hG�A�ޓ�z�A{��� c.U�]���S|�����줋"��'v}��J,$���rpTN4�l�������{{��wu��8��)�Q��'����b�Z�kb���"������@�a��<a�D�I��cH�W�{��mo�:زH�#J4I&�^�F���~�[�Y�;���
l���T,L��u*�rM�Y�a��QiH�pϮқƶ�zy��'L��>�-7+�4s�N
STj����-�d,qp�vDr*��/�Fc�5�ۥˌ�tTԶU�zr�&�g9h׸'�hV�s��w�Vk����rt��+�f��)W�f���U�J޼�Lz�/��Ѽ���/17YT�|)dT�l�J�F�68��@��S^�5'�����g���Y��b��f.曶��������J��/9U4ϓw���ĸgy���L&�m�KjY2,Ӽ{Sj���!�%��&��H���5~g��"�u��n7I��hY�ZU�]�=_��}�&�y���(��v
�;y�'	Z�'����� ݬ�/8u1w����u�(��j��&�t��}kd({�I���S��]��Z[˅v��\��n��F��ut�7�}�5'�!�B������Mm�N����o֫:c��Q�������������� ���Zq�{�=�hi�N����;�Vf�m�]������z�	.�Z�1��]73yy�Pf��M"M=�����U�rר_��9�e,~���
�Y��捍��k��wv:���Ԣ���B[0���69�z9�"ec[�#�vi��x�c�z/yŞ%�gk�ԃ�Md�o_���Ί�M>*��m����Üf+�K�T�AK���8�`Z�_3G�)�Y��NIn��]���v���UBy���Z��YW��V=D�JEuT���x���7C�v&K��4;����.9�};��Jq��we�y~QyR<��+��iy
�^��8�84�M��:��7~��v;���ݥ�5���$�mg�3=��L�	���g��Y��(-��vW�bc֜=֡��$��������x�qm�H�������.T�ӤXC�`}`�T�t#s�4�F-��MתW���W�m��N���}����"POV��"��Y�JZ~��AX	lm_R�=�]�9��+�#3�	���~��y]���,y��83n�����
+]�3�FP��ϩp�Kp%hq�B��gz6�!��� |�I�i����8��o�n-�w��	P��Z�S>^s���u�*V���//)����(�̺��m��ԁ�Qxc�#L�I�m�5�z}�V���ϗ��R�����v J��zշ;�9�éeޛ;:������_Y��6�7j/��ӡ/��?!"����&�ʞ�c��0*��5����1�Y;n���^�R�{m���U ��ݼ�&� �k�u�Ck��U��\��xG[F�0{;�.+g *��UqV�s�q�9gP���Ύ��&�8�m����/=q��/2��=���i�{-���Y�8��f�W���������(�{�:OT��Z[�b�qH�令�����j��$�kЫ�.p�����
�׷:a~ɗ}��.޿l����<L.��]�1�*8u�V��������9�0v�e~��%�ݞ��X&�ы���A�t|��3� ��
r�rį��FN��puk��W>�~�ތlS�.�Kt��PaE�Qs�;�ƞ����ZJSL��=w�����x��y�j��Mk��}JN=���P���XX��.���H|��ﳏ�.�:����c%*x��4q�u��l�ZJ�"�*�l�f���l�m�������o��C,�j� Lzzk ���ø�^��r��l�fԭF�m��[�ݸ���T�>*g��iZkK�oA��^� c�b�c��t.�]��A��]v�r0���#�N��p\�nOxG�5�X��e��V�+[��1&wh[z�sBs7�ѭ�pX�!��-�YN=�с5u7Z���,�b=Ӕ&nӃ��}Q�@GgBn�_�Y�>��TO��=��B�[{��ӓ6����@+5��a����_"�tu'X
�Ѡj���5�\��o*Y�}gKV�YM*��@��܍l�8��\;&�l�]���D7;�i����V�ǹ��G���@��V/.lT�mv�{Wn �ǳZ�B�\b�p���8|5�)��C�(3#��܌5����v������[+u��r��OL��ul��!֬Q��w@�o�� 
��ux�ޣ��DW���Z
bwi��n*W̸��t:�-Z�8v�Z v��68��T�P��'x2�2�xsPk��;�k�5�^YX�%��ڴ�R'5��m���*k��e ��x5�Z0�z�)F�b΍]�\�Wv*˥�Y�(�d_j��2-����<W��}���=o!ܷ��C�,���
����U���B0	���Ń��oׄ��B̐$G81;w�Y������*�X;)#1��n%����iS��NL�t]�[G!d��jܙ9z�[s�5�o+�)�m�A���޻y��tj�{��!��J��Y��0y�Է[���:��N������<�]�kr����Qm<G�ZN����u[2�N��;�� =y�y5ڛu*n���E[�T�!\)����[S�8�GKw��Θ�Ҏ���]�n˷�oJ}P/��`U;�lh�ݘԺ�.u�Н���8��c��U�rʆ"�
jU��<��%�H4e'1�H��2E}����@�S��6 ��I��B�\��g=3,Ji��u˻�>Qӱ��!����&�
< ���O���ݣ�O5"��z���6cQf�6';A���N��"��'�7Y�pa���w��O]Hi9��^��c/�L-���o��v�j�{�Kk����<uV�O��y���I�p1�+��O;*�g������ᦈ���1��:�u2����$�V^�^�Q��1#2���h3�ђ��N�zm(0�َ��=/�v ��2�kA�%*Y���#V�t�;,�Y��̳AL8�t��:U �"-
B!1�ї�T획KQ���4�
͐�����J>F���"���e�X��FI@�3����_���X�wU<�
e�����$�j�J(<�:���g�����׎��T`1��cUQR�T�xu!@=C�T���{~�_��며y�Q�KM$�$�eJ�g
��{z~��_��O�<����Ji��ɦ����I��Q�f_p29�}�L�ޞ߯����ؠ)�d=���(sq��;��4��g]t,�����ǎ�����%+M&�rN���*�@���*�$��><x�׻a�2{9 P��@]�E���~�y*tJU	BO���������ȣez��ʑ���
\�-�(��r*�U�����W%�i3�|��S�1�i(:�>��;.U���~Q��!�ZΉ���:��p���\��-̙ٔE��s�� %(��1s��Qs#n6���LAș���^ߺ�_�+g�f�{Ey�-"D�L����_I���'��(�"`���
Z&vH���m1ܽ�8͚>�l��@hlFD�{�
��Y��e�Di9BW�ʆ\w�N�=�0_L�-��ht��]�a|L2P�������76,��Y�r�s)�(������_ſ0�]5��.�ݗ7u}A�l"ۤ�������S�b�Xk���t��	T�+5#t"�!R���j'���ݨ�� j*@�iTԛ�v���V���.Rib�N�[�`wa=��F���f�)-��+̧�>��>��@Weo��H�Fn;U��%�۷�l�%����m r�g�>�+/ѭm���6����i�������>CV��M��+PeQzB�Fב���eV+�DH��d3���̾y�C���#/9���H�UnO[=	���d�z.3��ԍ~��Ae+~�{85� �W����W;���";�yu��v].����q� Ԣ-�b5�=BwNXn���G`;��K%-��q���/���Mڲ#�@�fn��)V��7P�.���KNS�3o�\ie�ھ7���5f�����׏�¯�|�y���ZV<*޾���oC�&>V���rʨ�-i��%]d�-m���x��|-�-���Ⱥ�c��dր����:�Pc���tR�[�}/��D����٬�a�@|$P�h�{�������ߚǳ�=��6��&�w<�R�Wy�67\y�����l��u�/�^��<�?8�V8�������A3���~�O��]
�e!7:�c5����ec�&��\������o�L�H���5���}\Z���"{Ս�Dm��<� �F*�]-7�CUl���Y)�2�9a=|(�cX�a��m*.��A����]��ˡY�:-d6We6�q��d���37W�U^�-�.�gvwY��޿=W��LZ*�0a���x���D�#4x��-�%cѽc���G;��`?|�u�U�s�ch30�r��S�g���~�\9���.���v�$��cq���˖��E�>�43����:.���pT?:ui����4\�z)&2Lq���]z��s�˙ƺ�Z�c�mc��KJYȹQ 
;:�n'
����p��p�5h����D�t:��!�*^Z��Ar ���� ��h8��4� ƀ��PW3��ķ�v�G�'�Ŀj�X6	`���>R��x�\�+v�i�X�n�Ϥ*�TC��s�/J����]M}[��j��#��K�G��3�KY��pgKY�V����I������u=�*\�j��^em%s�,��j�w�˓�-a��:�=���eX �H��<��T^�nB�������mv�I��|��j�wOE�<U��u�3��q�y�P'�¾���ss:Yޓ��2b���0%ixyf�Fy^�[<lć,7_�O��+%�ݛ��Ö�6<?]�'7t���㩶I6^V킲ueGR��6<%�w��v�ب�v�����s�U;Y�7���<�iC�rBFض��,V���nR�z��Vn�a�?���Kz詛�ޫ���n���Ь�v42��l���7�{�U���(�@�D$hOV��%�l�׮���׸׸�36�2�Q�]���5��α�=�j�ۖKZ �qTkE����f!���P�Ж�F�c��ePK[D':�T�N�,�5>��v�:��9%��̈֕F�Pu9.��[��xP���Jά�^�݊�7B�0e��ww��������A�k=��M�u���>���_��td����fT;��uE^��[2o�xOV�Fm6�rĊ�`�o�|�7�C��W&�Z�ny!o;Cw-m���3D��;V96,ć�a���x�'�}P�F�<�ا��ֶh�����EjU���n<x_��Q�*�롵H����VNn����f�OI��x��{k��v�$W=:=|$< ݼ�A���ۜ�ژ�.NȕxE����\Z6�W�j殻�-��MH�`�ҧ)v;U��2e���/rЅ�c���`�6�[�5�<��U~��:�+��y�oN.�OsOo�_�k����3��ޱS�"���=s�X"�!���	烽��G*4�FVե��afL�����Z�j�?�PPư�.�hUuB���8�gyH�IZU���+��g�^D��Č��zRm����>���6]��))�cU@���N��u֒��[��H�y|�+%��{R�c�Ҩ$�̫��C0�c��bJ����D�Zp���j<���c3� �f�Њv9^���][Vn�����ߥ�|Z�(��5�N%-Ѿ<��Dp�n!���?���З�"�5�3����lq]4��9qU7�od�B=u�d�>�5��M�-�N(�Z#9*�z�y[�oQ6�秜%���T�����<\�J5m���j~ֆ�y���R�>�)�\^؃V^0�o*:��i�Hj�F�b��t�?@w��=��FoT��C�����
Pמ��^�G�	v��� J����]��ю'</-y�Cqh�v�!�^�	�9E@g��\v؞"�^��rU�sєD8&�	��o6Hn,1-�5�..A�k1���h��.n�?=��q-�K���׌v�Ĩ>+���q�]u��:��m��Z���3^M�1k!�}WX��٠`�� 1��\��U[�e��C`��e�W��!a������qd���w�C"��z�l��cǾ��U>?}�d#9�����byɟr�~�o^0���m^���"2�C�j��3��ԅZ��v�5asw���YR94?ȝ��z�/����!���ix����ʗCT�_CAO"���z �{y4���'sz��c��������Tv4��2��h�,P3�hj�߄%���u���Ը?
�?�͈��G��{y&���'�)}q�\��H��"�.b����݅����/��"8�O^�GoI�X� -�x�k�S��U��ܽ�h�]b��'����v�-���>�Ġs�H�@�VM,(�V*�Do`FC]��{4�[�:yf�trͧ9kL��܎<�dJ������J�ʹ�<oLU���a��C]�S����$�Go�g��;�m.��[��I	�>���]n���T�[M�҃+��O�,���ڗ`m;ó�`Ǉȑ���ٷ	�
W΋�u����-�**=���r�N���r�.ֈ���#����ܺÝ�t�:�3��Xg���"���k^In7�\��uI5������QG����HEz�ly;���s��gw=U̝\f\�M2�w�Je@zΪ*�v�O[�'cĊ��}�RP斴`�u��Ϣ��F���n�M*j�Y���DLȪ��G�[��	,�F���HG��e�D�K��um9�v�2�¾�>��Qt� ҝ�:���eu:��֡�3� �)������Z��G{��;×s�h,����",�R{P�mt�<-��"��?�E/�!�t�����|�������Ν���M����:DٹY",�g,�;��+������};?��5#Ō;��/��an�S�5�`��ɼOq����lS������u�ޫ|�:'g^���w����y;+�EV�3}`s�N���_`誱��/���%$)�!^��X�c���>�x��Y�D�P�gt�e������_�m�Tg��c34�Q܂���wJ5ޜ]/d��Ĝ�Lblzt�-�%i��A��#�ʪ+���_�Y�/I��M6�l���a4�Bt�j�a�誛O�C�{�u(���f��E�[I\� �Mv��.�'I���o�2�}��S[ߤ�������~��ӻB��.j0 � >7��f�nbA�7%ك�"y��Ic@�n��5v�C���z�H��8�tk�MCJuXfo'�o_Q��x�o���\U\,��]�@}OrB���W(�(iӃ��2��Y�Z�����×���{y+� ^��QZoV^����ӎe]
�{V5�y�=˓��J�2L�x��|_f���eH[���tV@�./rV�#���<��ηRrȪ�4�T�qlk*b��"��:��f���=o� 2�Oow�}#�W�-����o�D�znghą���Ǆ����n́{:EwJ��@ �g����Eb��[ӽs^)�Љ��À��^�����|�����5��j�c�Tߨ���]$T�w`�!T��56�p���O�x��>�7��	�o"�:cqi���Eە�fM�V-�&��̴ӥ�T�}���#]�~`Qy�ngfsj�6�s;�;��qק���]���v �O�����\������Q�R�]�Y��U���F^��D=0r�nt�v��K����+��p�p�Z ����q����MWU�y��z�h����O}4"�z6B���c��黂�pj1�;��ȑo�{W�T^.nh���-b�L�����@��@='ν|����ɭ������v&�mA���&�m���d���S}��B�w�3���� ������3�<-V��i��2c���5�M�V�7r�G�+s�r�@Fr�X��u_S��y4Oe����K��ri�2qs����h�ՙ6���4��\�m%�7mne�Ѿ.�sZ�n��~��,�в,�Χ������d�Isnz�th/f���v�
��xE> �"2��˜����+�ظ�G�0.�Tzp�ꟹ�}��uj8�:e��95G}Y��X�#�f!6�'
q�V�u��l{�>�[q����Z�|s����vN�q����t��NP%$mmb���O�ʼc2�[]����yHB�nR}���!���b�y;"�=W+����B}gmu��*r�%�[��I����j�?C��]��g}^�;�%4�_�Ģf���aŸ�w�a��*��5�G*n�������%��j>�cbc.Q����ұYΤ"t�B^+՞�蕫j����A��M
�g;l�sH�p��A��PCf7V[f�K��i��8�,D��������0n�K8���Mt�M#�j���6޼�z�1��r�x�nF�u��kp೿V���E��ױv�~_�h��*�	]+�F����x$��N�ְ6+��J��T�O�Q-����v�K��ԯ�+ݾ�SޢUmp�f�ƙ{�(�:��)ku���%xcMI����|���[|�۾8���ￏ���y�z7��,�K_@��r�:��YF��7\y��q�����R�I�D�z�˫�=t94\="�Fs�1�&��� ��#����v{�kg�4Lz^.��2�3i�)�/Gz(��|�g�9!����n��T�ᅺ���8�� x_��(�O@ms�U9�ӎ�0��j����w�}�ʳ�4�ʝЛy�U�����6���1�����Y�b� ��ͯ�,ڎ̀8�/�4aoM��.����m���RS��f�U#����[��n�#[8�)���ȫ1Ϊo�2(쬳kRV�Dk{�cѾm�ƍu]��Kdq�|&�eX˲���5��Ǥʽ�$i~�uBd��o��n�[x��Ý�YU��dӸΫ�|�W���Z�	-�6�%iR�w���qUgluT��.��	���T7�5�'��R��^ 0��s�=�l�XAq�f����7�b� ��i��ch
�f�ו!f��>�2) �ҳpo8��㧵��B�������|�3 ��W�VF\K3.�&
}�+�2UǄ���p>��%8TZj^`G cv
�.�2{b�}-Z�Vd�P�*���7Ct��
���q���ۏ��&Iw˒K*����.箸�yr�fcv�Vo`�(�a�W=�{:n���vDR�#���F�k꼛#�fL�8���U�t{9�}����.�[�\����E��uc�ۛd�Tl֭Ĉ�U�|��Mҩ��t'*�Au�Y���kް����#N'Y/Th8�ʵbc2G0��Vu�6��e(�xrBnm���P�֜�: ����4���(�����ۺU>��cz�srԒ�J��@*���%���4Ѿ�1�����}��kJ���=��q���Ln��O�(���
ZwwJ>G�Y���y�}��E����'{�i�;�Z�J�EiD���n�a���	�]�f��v�Zw+��/b����P�ˇB�[;2q��1��1
���яx}���CT��X�qv+��:V�d��Z�J�㊰��b⦁�t�����G7qwfc��J����b�r�M�B���`��J�'C���L|�y7�4������Y���O�*x�{q�Z2=�*��l#10*�$����
ľ�)'_,�������z�:2��!2����Q�%:,�U+]MKa2����sh<�5"��Y�uIt�+ҩZj%��en- [�R{��ӳO���t�����L��o֑wDg����
z� �c�ա��'�@^���jܾBĔ��O�"l�(c��(�~�­�m�)R���3�|6�/'3��j,�]��V��H$�����K	�P���J��Ӳ{I��ܓ�M��݅��n�u��D���v�b���q��� �p�:���}�Nr��%ܹyI��!p߬�oJ�ʐH��ł��2�7n�3NH�G��H؝b×;.�B��v�瀝o�5�%�<)�Y��-���bj�4P2���־C���dȟ-�K�)j�.���PZ��X�u{��*�uV�)��~���`|8Ů��"������xm�g;\�0{r�g&M�4=��ۜQF��/��_MYp*��CZ�Ln��+�C^�D���3z����GL�.�H��7W�]� S����z`���+z�*��;�
n�(2v�W)jr� :R��:��]�,�������%(u����K1Y��L��Z�V�����c�e��|e� �F�pr�Jԓ�n�D�$���]���e��v�"�8�	X�pq�.���Y}\�[��f����f�]�tN=£�E��j�sw��G� ����/�73�K��$��,!�"M�h�!.2ف�d B-�a���T-�b�H��.
Uv1�d�)Yh;�T���9�u]dy��]=��G�������(��(�O��/Il(d��H��������]Gd��'R��$H�E)�HUP�b�P|��h�x�����㼇���+�H�ug0L�����Ru&}��Od�g�����~���"��H�Pd5��pe��OqFAJ�I�2c�Ƿ�<}�k�'��O�?d�@���{�{����%����~�]�`9�_;�&���*��9}�2
�	�������uM��)iC���A���\���(h����	�?�>�x�Ԕ? 0����:�6ʁ�G�7�%׷���׎��a�\���	��%�$��%))�ZS�T�a��<��D�iB���N���]O�܍�3:�u�uv	$#6�2���5sSjv�8_ql_V:v��N�A:ӳR�u�_wS�A/�^����K��ve��N�*�q��4�%��"���p��߸����f�d�x˽'J�)����|��i����tY�7�OW��1.�Dpث��x�u+y�D�`:H��ąf��r��Ɵ�䕝R����qߛ^��45O_k7He�S��E�����aQ]�嬴EZ;[#k�/����*#b�]��[�6�y��40oGs;�3�\��e=e�I�$R�q�֦^i�q����b`�L �웏>�SꛯwO���Y���KQ���#md:����3�f�sZ�iM�����B��*�������q>��T��¶�qV�'��=�o��U�)t�S�{���IͿf�0�XQ�z�K6S�����2k��X϶����xs�(<�Cm+tb���m�s�}���g�.!f�V�:�*���!��o��G�[���Oo30(y�QKf&�]O�8��cV������#L����v*s��~����/xKwr�ޯY|�L���>]tw���M�V�ݗ�[ͼVo&�z�s��yB�̧p��pd�j�0�/,~�������}ٍ=�2��y�F>c��%Yn.َz���Y��*���Apd����7t*�`�l,X�C|X㽻�}�nk|2e�U�ϖ�	L4����J�s�x�$}�L��?wa�͙���O�`�$�Vy�Mf^l�ss��4Ҭ���Ɇ�Bb*�Iw~��>ҫhs*���#2�(i��(�z�����z�.$���V&� ��OYg���:NMg�ҏo+�T�;U!�
�r��=�lC����1/d� F�����5�m�,������v�=�S��3i�S-�բL��J}p�RG�eg��7���m���7�b���ћ�SM'�9i�\�n��OJ1k���3���t�]ǣϪ���.�J�}���{y�V�{#m��� � ��t��\U�Ŧ�ݚ���ʓ��pi��ZE�N��E�;���@6��C�p���{��SZ�0�5����V��m���N|O�^v-���4lɈ����nm^_R<{q�]
x�$�<Y�w2�X�X�圔�:(L�T�|1�Y�/�!���Хy�v���:@j�|.�+��O:qw\�k�"� 辙��7��'��N��xa߳v�;�T6S�9�.nd=W/�\�2���j�wV�y��kxڸ��Koٚ�r��ӕ��!3	X&��Q��ua�g�A�j'֚��k��B�(�Zst��d_���ک��6�nѳ[����'A�
�}�+���߆��S�9�n�<�y�+;���5K��TҜ˻ �A�O�O��� ���-s�l�,��^1 ��wՂ���v�*��$�7ۏ��{�_\�@^����������k������ǟXre�����W9��tO�c����j�˛��X���w)N"�N��m�U���ĳոoґ�͒��e��xˀ��ڽt��l�5��Z�Z����O��{6
��+�ٹ5��t>�i㧊�0�꤃�Y�ler�smxF�l�;"�W&�1oH}�]�&�t㶗^�.����8�U����{��o�U�F�>��z$��i�}�Ns�i��׾�!�\w�镻��w9׌��,v����d�#"�;�:�V&�1�Cȍ�#!���}y�]��#�D���[�J��b����6n��4��9P���&��w^��e�]*z�Y۽�N�l�����T��d����0fs�˧z�P�?;W����ֻ�	u�"y7��
����ٕ���t�Ǭ8+��rtub]�n��O�� �t�[���ZvH�wP��I�E\<���w=ڽ�\����V��NCΧ�۪,$c؅l�3`>�D~�2���n=���JoWs�wE�"3�>Ҥa4��M=ɶ�7���u�y���1FxwM/���3Y��Q���1�:�*8�K�%�ݧ��A}02ᶺĪ��U���Ռ%	v�9Θ
̋��>X��W@4zw�z���nT�V%\�'�7�5�.�^��#��N��p��T+l)"�|]O�M�_���cMߗ����*ʯR��Ϲ�'܂Ⱥ�gv�qx�M���D|e�&���ͬ@H���\E�}H��j�59P����
���'�;��W}ydEuG�V�G��}6����''+V4[l���[u�D���xh޺VB~>����8���nuMH�#����<_<͊N3c�B�,`¢�Ϋ�p�05M�E6½H�>u��
N�SkeZPg�Ҽ2�$}[K�F�<��w��N�rk��|�AO��8^�}hb-m��c�u��I�[d I-8�h5#��� ~���]�}2�ԭ�ζ5��C�Cc(?qث�N��B�"�o�X
V.��3j��y75���d�Vj���3�$��Uw l�D��Դ��9#�R�JWZ�Nam���mn�o��멤�/��0��ސ�/EI�	��zZj���5B��qELNeZ�%��KM�ݼ}�	�
�`��c���u�[��d��2L�^Cn���J�ga��m%�RX��� C��t�{2�f�6�~9�#�F�z�=q&�����	\'�4ݖJ��{��v���2�{�����PO�4o1���u������o_��ה�|��Z��ۍţr�2�2Z�fݴ�7q�}7zC�R&v��U��=tk�� 4ǉ�3P��WsU���i�:spp��e�i���X�=�*�:�ܨ�%����������1|���U2�^�Nd����͑�3�1+�vb�6��k��oT�^�o��u�����̤�(�/��L2����VY`*�)ep��x1֬L2�J]�u�*�[��P�=%��"��x��c橘F]�'K��\���1r±�.:���e<��A��NR��}0�XP4�UN|+j�����\ۭ��Ӗ�_7���� Ğioa�ˌv��:�~\ڍz7Qufr�GX�@O9�S\��dw
�:����u� k�΋f!�Z�C,��ܐz�:�g��������\B�7���T털�]�j�l�����[
�-*��`��&j�����b�B�?X��{&���d"�u�\���D3���)�4�g�U"�2,ʛ�u߶��Epk�E�|1*��ܒ��c~?t7l��<���QY���6����Sm�2NW����LJ(�xfE�oE��g���{!���k�MH^�j֢"�d�'��S�ۺ������<�=�]W!]v�r�\�eTW�����Uz�^wNȈ>��E����f���s��D�`��D�;z�QjuW��{]4�oMlCxV{!@��\�aosytnHH�Z[Ds�灇A<���UU@�����y�EM�o��НM���S�7g9v�U�Ց��iU���Y���a�,i�5v����i�dkl[lv�An���V��ͳ��o�!�f�
W9=�)Q�͔t�K^��u����$�x{��k-l3|[rꬥ
(Ϯ>}��*u��Ƽ��֤��ާ���xк����l�{O�:]�|xJ�p�~��otGȼu�a��Z���F&�#��h�Nw6U����tL��YRc���2#��]uA���@u�oU^?.S�gI^�㵔,�i��4�Z�aC�-��RQ1�2�:�L�M�o����e"]"�Ð���x\{�*�e?ܧ�S���;���hH���e�v����O�^�<	�cӨ	E
 �-�7���t����S�����u=�/��v^�j����SY����]�i߻ ��x��0(�ϟq�W@��w
8뚘�P=��ў�guT�6�[=��t[T�g���ϔ���|�#,.�N���E�(�����`�GCY��!���ٗ�%e O���5��Q�=���)Mu9��|1��uM�@Ub�x�Kl4��c�{ú9�,C�a��bU+j����l�#�,�Ǘ�E��+�8�A��ou�5���ʺ�PFt���!�r-�*�}Z>�+���.1>Z���'����3�[��\�<Z32i�Q��%�|�/�9q�7�N���"�rMr�����vӞ�HqZ7��0���+>�����~���4���9���Hk��QY��`��|�T���9�9��=�u��#z�r�mSzk�+��Ǫ�M�{�AD�9sY��^˦"αp��$K��y���'�}��[c�ҷo�G2���=�h~���6�-���jP�O��d al�d�4@��H�V�tuhڜZ:���ὲ8�q^X� ��>�K�u����A�a@���)�9 ���Nu�x�5o�<[کb���&�r�����:a����ە��܉����+�s]q]�֑�b�FtxB�vm�$�#P��\w�(�+h�x���U�<��O=Μ�}Ց�h���FEN4��)l�S������nR��X��l�u�`�ݾQ�1��*]��ct��É��q���<Ѻ\*�,Y�YSm;����*aQ�:��ݗ��,�}A/����Ɣ�I�������2j�MV M^z9�,������
/�C B#<�%[�Z�h|�:|-�q)�v�1/JXK��Y��=mgT&J�sN^�A�"+r*0^T��;"{�wm�T��Vv$-@�I")�M��Q$D$_��f��i�Q�|�{r�����q�A�����g��dy�x���Y"�.�_S�n
U ��:�'�����q�(@&�I4�za�ђ��B*}f�$*���+�דSk�����Z�=ޑ�<���J.�FA�KHx���i�u�\f��n�����������W��t���t}/qU�W�L|a���~�*+�X���\�MW�L�tf�dQ�t�M�%wR���c1���W}љNu�;���<�Pʭ;*)M�7#�t%�
����x4o�������ә3�T�-�:��~'�F���3�������;�r0����g�Y���{h�%9UW;�yL5/Jq�]�΁l3K��&C�<��a.��$�x�K2���ogV�ڢc۔	;��<�z=]A�����r��D8g�w�a��*���粨0}p0��oP�v���}��n�hy�����k�JrI�MҖ���$j��(U��|n��+��g���3�V��I}�5u�P�]!K�ɺ�j�3�-ћՉ��!��"�o]9+n�u�KY�&1�ǒ�^�Fm�h��Ѻ���u��_����z���	����<�r�&6(�4����t�J�8�r���56Ϙ��Ðy���n��q��	��J����L��+��˨�o5����zT�+v;�Ӑ6�er����wr��l�d��m���s_�(�n�uȝl���G��?w��1=1���O�ұCU����^A�0��f���l�~G�x�D��m���d[����܊�����h^'}�o7yg���T]�U�loj��b5�\�F�a����K2V^L��}��=��z��N4�<(��>����/�;�}�wx�C�����4�%66.Y�*�n��]�o�q��~�/�n�Zǳ��GP�I\2I���~�F{���{��l�蘆K��lǞ���H]]��mq앻-�hqg��Q	����Y͎��|{M>-%�@g�ݏm5G�6��݃A�.���ltt®��`�)u�ь�"�t�M������׭�z�ɝ/��9��[�д1�3.:�1�c��[y���6�g]n�<�d��'�TxY��j3�ڟ ��G�N��+3�(8c	�b�1�y�NN�9����}�Q���4�>3��
��5��IՍl��uqAte^l��k�}K"�"v��u۹�/JyQ�'�b���z�M��P�,�%X?CM��K����1��e.y#���l�G
O
�$�����
���`����]�#.\�0b�R9�w���ʐ#�<��+c�=�o�ɲnP�!,�w�D> C��x����b��ݎ��+���a��Ac��[{�k�˵�3V*^��K������R4"�xZ����U���\�B�s9�;�D��M��mq��V�$o�r�����1Z��J�K��،�y��Q{��v7#�+RݣڣԂ��(��	�]�'E�%�+|��-ld��7dG JcN���fS�Ԭ����N���v�R�}�nJ��F
:�{FE�*[݆̽`�0u�'�C��x���ʙ��܅���%�H��c��}��4�J�w�pPI-n/���p��hV�餭�N&�+*U�Qj�fWp;�,&�0�p���Wś����8�[;�����'��V�\"A�1K�� ���՘�V60�G�\e�W�nq���hv
���w�(ek��I���v�S{��绗6Ӯ�Z�G�3%����xE��3��l櫶rk�.�Ȉ�`�l�d.���y�9�Y��̬�v��ZЌAu�:śPu�	��'h��qk:�G9`@��Qє�ۥL���-�(���N��1��\Р���.
���gq���ڝvWh�d�l6�l�bb�|�mhg���-�h��T"� �x$�j���i9���Z��#Z%�ێ����s�]�V������p.T�u�x$�Kr�=w �G�b����XHL��Vͪ�sh�سe��7��F[ސ�il9�
�]���k)�#m\��s�o;�*(y�u�V���Z <u������5��U-0W[S�:Rob7j��E���^m��vi� ��̝�w���%1Ԣ�l쫿���c�d��t%L��,��7EǶ����gG�D����.�?`ܳj�ٱ�&�R,��t-�Na�寠R��F��(�|�e��=D�gJN$`���4���G�Vd��[Dɶ�u9��j���\��k=�5�<%X�^�Z�Ln��O\V� �4��m'K�6��%����<���돈ݡ��߯���'�]����
D� 2�\�
�9�t/PPD��	?�_^?�M�(y'p�B%r@�^@�f`-��C=��x�׎�yVY�5��܍~3�'w��dw�D�@d�Ò3�ۯ���Eڃ�!
������;���@d	ԇV]e�t�������sph��c!�-D�f+�e�gH)��E4=<x��We9	�=T���dK��]X%U'rd-'�e���O�����t>���B��f�d�M
p� t��0Y�����~�]O#�\�6�=���r+��C�N�_!�gx��oo�^<t���3��d eK��@����p+�!�uQ�%30J�f��O��u�u=u�d�ԟTFW��޿z�:�;�75�z���\�F�eu�M�E���U���P`ޒ�������۱e_n��PbN'PsI�-�2ȮJ��T���ە��ё��|Z�WYqT]��g��2�Ah����ս;4V�p��:�Nj�'�s�Y~Io��m[mr���ݙk���=�9���}[-ӭI���c��x!��-�[�:q�V����uc���іck��![�o���;஋&c���Ewg�}�Ҩt�41�+�mJ������ӽ�j&�7LH��i��=��[ڮ.���O)�0�ޮ�J�̩X���y7ۥ�����Y~Q|+'���}���>����Vƚ��ʺS��{G�K�~*A?o���^��G �����k\es#Y�9�����[�Y�zI���{у^/'�C>�;!i�i���F���̵�_�V�
Hϱh�9�;��^=՘�f�$�7?3ۻ��T�1�v�qhN�����	',�/j,d��Կx���;2k1N6!��Tb��&�ǜ�T�Յ3ҝ[8*�m��kׂw+#��4m^�ttaU
�^u tP���*�3�Y��㎥F"��ʡ�޷�6��+��҅�u��w"�;�X�7s����!��$q1>ӛ~��(��`�-Lo���3z�7��^�4z���o����!
�j��ѵ*�p���/�6��+$׍{���o��e�U햷/<���1���᦯~��o4�΄����'�s[y�#M��*��ӷ�=L���u�2׵+e4����Lu��X���٢�<���v�Lp�����xE�@�otz\̌H�fV՛�	]�9�e�n���%Nh�ݭ�~�}�����p���t��ێ�Q�|R�qQ�����F�,μȉ�\l��DV2�u�G�/�_����s^��r�y֎2�t]ޥ�`�W�{= ��u��Y��nA�	W�J��U����&z��Ow<���<����D��5	Z�U8u5�@���^����澒_�vwNi/�u�y:��[�Y��0�3���~�s�R��������2��Ǆ��)�4�e���:��g�5V�U!��#�� �{WeZ�Bj�ˡ��:NQ����n�����D�É)��ˌ�V�z
������"�	,�:��-�9�v-�d�oN���3��f��I���e9cVmi��uMK�|�i:ě{�4X�Str}{B�[F�����Q��T�O��Cߘ%�CNV�y�h�o3��]�}_]3���oO�5�VN��T�İ��x�;4m��Zl�z�i��k��f��^�L핔$�@i���=l�\ߩߢhA��g�g�d<�`- T
�����<]]�"hw����|S��GefM��9]�0gSb��n5��d@Vl_e��ʳ�7%��=·Um}���aoQ����vXd]�eX��j��a7mO��Rび�舼��#I���,�m޹j�EL��ۈ��P�Ɵ��}�z=�p�)%7�h��@ײQ���SP�9О�}��'�H*����t����u�`Ut:Od'�ⶼ	��Ռ�s��N���Q�7yk/v��&��[�مQ0=�*�Ӭ����0�m���NĻ�z�=���?�^�	~�	N�Pm�Y���)lN���KD�x~i/U1�v"ڻz�[r�#�gG�H��!��-�#K��'�r���Duz�<�G�����0-�u�s������
<@e��k�+���1�d\�w*O#�M0�oU#зώk1��eG�ݫ�Î���g#����L=_�m������ܥzl^ߺ�<�,��h8��~Y"�?��y�7\4�Q"��[v��=d6A�rK����	Vm�guX�56�뒇�GqG_S���[�dWoC՞�HW^��q&Cr�C���0I!bΡ����ӫ|~�W���ҭ#��|�\��T=��G}⊛w�0��$���:z��L�j�o��8�ӹ"f
�w��`�3�1V��l�Ew+eL�ͺ����[�M�~#S(��h��F�����W5�yU޻���SdVNf:"v� ���C�8zq��]��ݖ��2{�C���P<9��ͼj���_ L3��¬���uO�w�Z:=���1�c��e/����;�<7�U�_[��.$����� 2am-E`�1�e���-F��b�|�d�)�pf����Xn
;=J`��.��5pD
�If%ʳe�Ⱥw[)��/���[��d�6fZ^�b�U�b3b�מʑ�3���c^e�G]	ޭ�~Q�Q����=ѢXafj(�nJ�$^Θ�ٸqss?�z�@.��o��,��{r3��On�Kݧ�i8�������3_k٫�ָ�����w��"��nڎ�v�eq� �V�
�F�s9�a��Ǉ��|ς�ʮg���MV¥�|�$2X��n��}�I�w���B��=�E>ԥ��)��gV��v�S�����9���u,9ۯcR�mK+]^K	T�"-����\��lw<��О���w�kkCC� ����w�,����[EfU�y�u�,얻Ү�ۦj�l�އ�<��[`�����iG�^x��C��z�]-���$��\��!�j��w[^�R�,��>��Ca�A�����]YQ�u?k�i'�v;2�c�Xo'bl�@���W�KEj��[��j�L\ի;�:��Ew���'���n��ta�z�.>��n;�ّ~��	�*Uϙ������;U�縘���d��=�e{!Kog�
3%��3��F�8��뻁�r���՝�B`� �A�Cjѳ2#LQӴ0�6�u��0:�]����ì)��ѥ<�ճ,�Hє��"�Cpt���ήH� �M���;����6�MϾ'uW�y{l�8��;��	��5�3m�swbl���~�x�������M�Z�כ�g�!R9t��M�Wnq����H0�«;��z�6���O�޿agmS��!=[Em��ZWЃ�����γ��e�pk��[:h�gݠuO���&x��s�H�����x���.(jyw�
�ԍ�(���7鐙��e5[o��9[�N	�� �W8��z/����d�Φ��L�;���ݍ'*�v�h{\z]�F
�5��3ɏK��k-iX�V�݌�D����J��Cjɧ��[n �4��X�U!��j�lz�x	4ʉ:n�/���})j������7����Z�;�6�X{�[X��װ����;ў1��驽1I�d��u�J�\cwG-�^��ma7l ��ZTF�WsML�a��,"V���t�Y�
(�ٳl�����5c��x-��I�܏KT�Z�fD6��Gd�]�N����x�x�E�T�q×�ק��JC�"�!q��"7��i����}�:/os6�bް��8o���}3?c�|_`��\
eY'��T�d��]���IX��\�Uv�ā~p@�d�-&YD�!�Q���l*��g��X% �m�$�����M��_z�`�l܇�qlGF�*L/ga�gky��ęy��ʾի�K^Гw:*�*X/y}e'V�+�c��$��ݣy�z�#��z�^V�-��U�\��;-�����әX���Y�{tz�P����}�|WrV˺q^�:�� Y�Rfi��[A5[�w��Q�VMR�5n��۫-#y��T��凷+<f6'#b��:�`�[��LAوV���J��ٶ�73Κ��"	i�{��!�Uw���y϶$�r�zD�p���	��0��w��Ү�FH���uy���ϙ�v���r^��P�O�bD�fF�Yz�Ҏ+���5P^��=/����i�g5��\Z�X�mf�~~���,3S��bD[f��U�È���qVÖ�Nx���΋��:��u��L�T�~F��|/�^��S&��9��Y�ou��&0 �5�N���Up�yYf���2�н�X�di�}t���3�6�k��0�����4�d�n�Ͳ%�N����d��N�����{�'��_ ���iQƷ��V!�7^���酯_��]uq�*�9�K0\E�u; '���u6���lB�:�8��-3���SRJ�6By�+k�Nj�{�7��r��4�Wx�FKZ��tZk�5��_&S^Y�.�;Y��`r��xyy�a?�ߚ[��n�(-�h���r)Xu���PU�T\*�)���[+k 1�E��n�
	8UY�Y��f��`�g{���z��=<CE�?����~���VT���n �Q���LpD>���� �7�����V��J�ӽ\�KV*픺�f��������W��d^tf�T�z�ꞶD���J޾E�J#H��J��j��Ѹ��b�ou,ާ�bd_�*b�zccԢVnm�Wu!��~yޝ�Gw���`�"�]ٔ*����b#R�3��ޑ8��g�����Տ����yό�����Gf���P�fs8Q��pj�Z���U�M{�A��k�j��6���f{ta��t� h�@����^���h�	���.|�7Q�j�N:�Q�&�!-�ֶ�f����,VPV��#�]��.�GhY��;��D�����OR{`D�@ַu-�4��XDmz�Gm�6�����"M���mv�OG���3z��{-��ψۻZNM��=�Xm�4�6������l���br�I99�9�9���e�I��9J���u���Ռ3��NV��j�W��#�W@zU:��o������o�"� u���1d� �3}�m��<b��[�V���w�:����D#
z���=��U��!&&n�]�k�@��<P�䌀oZ�H�3����=�gv�H&��2���TϞ���L\���{"�7]F�d]����a�x��u��v��&@�N�52�wa�@n�!�wTH�ӽ3(��z8��P܊�Nm)&��[@��t���u��P�}��TVjZxtsL3{���ŀ.�焎�@�h����ͱ׏��I��U}䶔�)֕�øc7�Ze}��v�d��1��L�Q��yHh˳�4�O.�ʱDj���/��U���ͫMN��:ޫd�7遉�u3�ʂ+���yDt��rm�ɛv"ۢ���}��&?,9����۾�Fǻ\
��ˈn?��~�����h��9��d{�{=���}-�V؂4�§�k�Z�:&�s5��O<s���V�vf����v��t����� ��Kׯ]:����n ���߈�*^=.�9���$�?�5�}!��{3�w�W	�l� lAU��\�Qj򞢧C9a��_/�&��f��R_��O�;�TWVҟ]
�N���|���ܷ._6؇�׻XRn7��Uw�'*�6���O�����Ш6��G_�Z�8���y.�ƧOT��v�x`#���r�Lf�3�C��(=��h�De�(��^{�ز=�y:�zC6�����X(
��f����*�B~g�r�0��'~�'���1L��s�x��VʬV�[�9o
�hG���!���}��:ߟ���_�s1�* *��Q�k��@�ʈW��0�L�����b)���! �(�! Ȩ(! Ȣ�! ��������B� �QC `THED�`AHDD�a@H�e��D�d@�`TE@�`@�d�@��� � �P Q� � �@pA�P hQ�� E�P � D� κ zUBV��`Q�`F�XT`Q�`��^��V�Q`Q�eFD�`G���eB����Q�eF�@`Q�aR�Xa�	D�`� pq�p  ��Ώ�A�a��� ���"� �1$?��/7������Q� ?O� �����/���������A���?����w�_�����]�� ���������;�??�T
 *��{�����q�PDE���N*� �"'���������I���؇��
����z�~�����t���rz���'� ����?]�~� #�"�b�H,BD+,@��-"%% ģH�,J3"�- �,ȱ(�,@���H� ģ�@H�#,@�*�"Ҍ�,�"��H��1У@��,H� �+2- ���(ЌH��0,�,���Ҍ2
P�@3�-�0,H�2�H�ʳă,��,J0B��,��
�J�@�,@�$0,,��-�!*��,Ȳ�3�0��+*��,2,�$�$�$� ,�,�,Ȳ���"�� ��*ċ0,��2H�(�$� H�(�ċ�Ȱ���̂�,0,@Ҍ,´H1�+�,H,´�,@� ����,��
�#- @�"��,��Ă�(�-*�@��,�*"�R"
x�(* P��(�#B��
%�B�4 � �Ă�(�-
���c�����@E��
 @)���� �����_�P}���?�)����W����D\0?�����x'?��a�����?���Ϗ�QW����?���6@P~~�QW���?�?W_�����"(�������
� ���R`���=�������;�=�@vb���?��~����D_�~��P�~?x{����Г��?�?A�QW���@(�����o�`P���o��?p��ރ������;�t$���� *�̢`��i��5��!�������O���Ȉ�/�?�|`�<�E�/�~�~K'�@L�a_�������e5��*�@1A]�!�?���}�������P�(�B�J�DP�"*�*� ��B�
�R��	)(��UR�*��$��J%H����ڎ�{�$��*% ����AAP�AU*R�D������W  m�
�ҨR�Ҙ�m�E
�kV�d�TMi)Tn5N�����h�K`hZ�ؠ�U(i��T�@*ۀ.�A�H	 ��T@T�XE*+k�	S�����vْl�����ڰQ
 ��%� ��
c�P� �͂�ZԦl�m�j$��F�B5ن����!��%ke��kkfV��i�%b�V��b���̚RQE*�&��Y����ƔmA@�` Dd�Z����h-`
! 	�T�
p]���PM��f�4,��EhU
6�X��fR�M� %`�(T�9�9j�B��҅ i��R"�H�l�Ġ��`�T� (�F�7g �D�6�A�Ql��,� �X����I�lh�@  P �� RA ����R�4�`��р� 4)�IIUC@  �   H�4����i'�M�6Q��&�ځ�~%*��I&��h��c�2b`b0#L1&L0I�I����    h׳N����B"[�-k�Ҷ��TAw��M&sPQ�~�2�� �t"��Z2>�4�A,�~�&����T�����I�k[��Umer�}W��kZ���y���j��jͶ���((� ��v�cZ�?n�=\��F��)3v���&r	�%b:�e�&�K��q�m%�x�l�Lm($��� $DKl&	��J��E
1��@�SAD�K�' P�$H��
 ҌFሠE�LI�ۂ'�!��L�L�I	m�d)2B(B�d"IFYq���H��4S}J7-�!4�F0�����b*b!36\PH?�,��@�5-����m|�sS,�fhۆ�cv�s{�aX ݧ-9��̑���`����)��F��e�
�l-v�/!�%�w �1���h��O�	�߆�lf<ܳ�Re��eضmn*� �[Rm]�S�r�{�������j�]��)�
�� �iܠjVL�4�Vó�/kp��^�|�� a<=������s�)TMK�i,c�Y۹�E����'	�f�lA}���B2�U��p��U���UF�.�Cʗy'�H�����-�#��0�\��ʦ�7 ݴ�N���k5��[�1�qd�՗5k�8�V�n�Ծ�)jk �2�!�Ǔ1S�{(J?f�໊R*�I<�UB[*�wb��T�h7���Bj��˛��N[�d�6�R�L�ͧ��q�R�DT�f������:I^e�ޠd�����`'���.j��̙�/a�w3	�w�7���L�i�����LX�kwq��&�u���T�$�	����+^�d�����u�bZ��K&�t)����f���NO��5A�t��f�/&�X\I�fdэ:)]���!zs3&��
YIШ�C5V�S�hU!+Y�4�t0J����:�"�YC��T�Đ�2�L��/�w5UʨA��u�Э�j|�E1w�u�%�H+�����eU��J�q���9F�_e;5�����`2LNd����ַg�"������bK���6Q�8��Uj�Cl'1��Ʀ����a5Wp�[�f8+-�I+��j�$Cw���/NmM�f���HV$pϕKj�f�.�;�I6��ԋ�Sn��#*8EZ���;����*]�:��
�T��kt�Oko+��Q!c��-����qkR�ЫW2���If����L�fƝcv�3,1P�3m�������m2�L�����s\N*͹�����)N23���Fv�,��D�*�L�bS��n+��Ir�ը*f���_n�j�)YT�)�k1SsE�A�3��ꬼ˚�d��!�����dz��CB�Ğ����D*ݡ��`�CU�3	1� ����`��p�+az幺ld��/-z]`&��5�U�Ʒ)4�Ad��V�2��sے�TEGp���[,�U�ѻrL@��L�%m���kv�OU��a�6ەpJ��:��I۸���ʼ8/w'$�4-��r�6����Y &˱�[�f�2��+V��Qҥ�Z�J>L�6_ԖA��#k���#;��<d�vZ�ԛJa�[����y�Jݤ���p$X腕cVLdVT��vr��=X��
YXB�{�Yɶ%���4�i��c4��v��Y�����*�,�sph��T�um�� h���j3v��i��T��K5`�ݗ�0�k!lGИZ���ղ�����2�a����+�)+�g>�9�ӫ!�@L��l�lf`wJ
���@N*Շ�VĹ3kAjE��Z�8اF�Fmm��1Z6\���ktc7�0t�� ۟fUۂ�<��S4*��d�hwD�GJ�a��u��r�X�"��i�,0}<:]��HY��ǔ6��b%y���-�Y��#��D�74V��T�#Ad'F�c�QN�"�Mn��x�+;+spܳ���1����Q�=˘�Ɏ��r��d�J�����F�se��	����=�6��ڙ�����L�:���Kr�@��PU�%�laB�n�#Jj'Dvn��C�vV�I�cD�@��M*�Y��f�q�w�S�LJcjO���MklB31���V b`��rC6]IOh�FB袆8�����!��B�mU�$X�F��!l:��+��b�r]��G(U��!�����xe#��K�T2\��%�,7NeC�T_'-��eլ�5��q�֝o,T��[�
xM�[�������꽢l�����n��1�r���h�5U(^G+u4��n�ʹh��щ�����䙈xD��-epeUd&;��AyRG0���U�֔KS�d]��J�^ِ�N���b%*U�bSdRC2��U��lFv���7F��J�ۓ�DZ[����Qr��9��	Ɍf7v�d�[��/�ܺ$6����v�U�A}a:ז�e��IC�S��Em
�oLV�"�ѳyּje%S�Ɨ���,�1b{��[�)Z��ֽ�e��6GK�]����"�r6���qg�;�����.�3jm�=�`n�Ê�c/^l?-"���hY ���`X@z�#���c�O����U��4[����T�Y��q���D�Ʋ�ު`�����4%Q3��:ȳ�?M݅��9GI�B,�sl\�[�cX5�HC5�ы\ dDm�Gw|���&�����t��!\w��;W(8M�&��ȍc�Ѣ]
�3U�:-x�x�ь ���t�m;؋^�MӸn">[��8�����;A��cQ�����UoC�̼s��r�nI��w]JKw�(^ m�ͫ���8^�A���7�����G��)�>���63WSe�W�Ҽղ�M����d����E�����A��X�6�m桤�
�T�JXz���O5˧�����;u�(*LT�t\t>�5іt�@�\ȉM�h�ƫ�I�c�*aoDY>��t,�Y(�s%)V=4�!�GǷ(��9/m[2c�f:���ՠ�:ȬKr���K��eܬ�6Z�MV��C8�wM�Ãs$Iś�R�;�V��Qd'TkBu��)ނ�u�P潪��Z\SP�\ �{�L�ݛ&�ّV�ջ�M�Km�n/�,֫6�,�y�_�[����2�(�DQ�F��Xӈ��'76^�;���V=98�{"W{NVۚ�=��b�e��:���xL�4\�v�yOi�,�r�@i�N<���ku�t�9TXbR��/[ӕlY��չ�nA�]���.�J�j�P������	*�l3:�h�rL�t��[7ٴ����{�ÁI�T5�P3WJ���s��ʖ۫r� �˷��6�B�.�䔲���q��Y(�E7�(�:�E1-՚H�M0�d��!���1bؚ��KKƞ��e�h�-��(�N-��R��W�IUѸ�[�$.��0Buf[!�uU켼���%�j�KJۖ1��s>̺JI��""��Z����N\��f�l��L�V��jm
�H��*�Sl��:ʗ�\���dDK�	�o��K$[�đ���6LD3�q @MD�M� ���a$d$�A����2�4�IFa���R"q�gђĊ2J��K� 	)#���g�FBh6��$�B!1����!L!	J} l��ɴSF_4�i"�d$�e�X���&�)�>P�L�>?6��\%��L�?I��`8 �!�5\F�n�V�a��lc=�CU�b`퉮�6t�\6wMaP�ݱ����달C�j�%J@륛n�낊uO��P��NҝEVJ�i��´h�;E�;�nQ��k���1d*໡o�˱�� �U2�^�V��o
9M7}��L��}M���U��bӪ��BR��,���ҬS����FgZ�1kO)E_]�x�.�K5�6Ů�ni�5b�;�m�;�̧J��Y6�3�p;��Fh)7z�ݼ�m����۽��Y��>��%��w���~zYyN��Wҝ�$Gr���X���C3KiǤff������d���c�B�vද��F�)�e��pY�s�Kb_S��w�Xˇ���`4�j]p�����IAh8¶�R�aܬ�4To���@[�y"ˌ���;^��.�|p��[W�M�ʝ��Ypp��\��(4x��̡�o>o<h��ݶ��Ȇ�hj�l(�np�ށvT�8����ڏ$�:��ϳ2��A��,蕹#��.��m�t�m��ѽb�� (�=�}QG��<#��=�blu\B��sX�leԭ�G��췯��r�$�'S]ƺ�g[å����Ȳ��N�qJ<��V��l�I8\�r ݓƱLdQ^�kMF��	�z�wddp����aokrs��%\�u̠��e�u��d���C�azzlUb�d+J�2yE�2^�mF�DTT7��Q�������SN-��!��F�TBt	��ܾؓx�c���	�����L���M��Z9���[�6��Xn�j���Mh�;H�9�Ԗ�cC~/ܗ��K���A��gm���4�}�ʏjgo�a'*����Q�FkԦ���ؙ��+e��q�m���O/YTS^��_�����"��Wp��I�¬�\��6�GQWn���=J�Ɲ�UB�͆����Z�u}{�R�E�{v��ǿd]��s2��(���^�gE�^m��.qmT��ӷNw{�,.Z� �Bq�¯0��`��d����N>ެ�U��*.����.�ev�t���*�u��O^�n�۪�E�dg��[E�C`�bP�vz>h(����.p m@�ui��6Ga��VM��ĸ����CgZ��f,�2�9	��Kgg�6s�+ۨw)�ː�v��H�<_Xz��(L�/ 8�r�7V�P���KZ�4�K�.0gP���:ʮ\�d�:�"��̃�0S���'r�m��Ӓ�N�;�{�כ'P�W�`����J�f��n� X�*�s	ڮޔ��Dt{�κw��f���zz��9jD��~������=t��|���=���\i�U��j��a�{��	V3+�V���1>L��T��S��J�ZU��q쨎_�K6��A�x��9�Rޮ����켩9�{�WXYÛ����x�Hm���5՝����7Ij�"��1!tXչ�Y�Z��qu-�u-3+o%$[��7Vd�:rYW]ú\й.mé��V�2
IBq71
���n���8��*�qc��*�T*v�pR�f�j�z�4Ņ�*�P��B�k��v�:RX�,�^Fk����#.�:+^7��eյ�v���;�렁��C���T�nbή��	2�<P�isK�՘��U�	�$�]:i��w!0��,.�2`ߦ�/�gp>�%��8�Up�����:�$��jɖ	*��6�Ÿ�^v�/�5gN�;������2�B�Ի�c��g�\v��B_]�=��s �ֶ#{è�Q�9ή"��d��
0eh��F�=	���ո�u�r��"��E�D�U�]�bĈq�l��-���E�:s��T���޻J;q^�R8�E��.˷ϱi�/3p�дqӼD@�L�Υ:����n�6���ֶƙ�Z5�[�{�\{��jY��9*![V�P���9��C9�8��aI��f=kמu��æ��a�m�٫���&���0�ܼ�glv y��ɫ�v!-�ݒޚr�V�Ps��ʞH*�0�ى�n��za�i�ɺ0�#�w9[C��KGi"�k����(nwj���+H��n�cY�9�>�J�W,꿬w�@�����_+/z���3G<ۂ?�� V�`;c���~��h�O6��
�%�TH5*���S����La��xf�Ԓ�v�W�g�����f#E��ps�Xzu�#�j���y��y��<ǒ�x�[����=[��1�ۤ-����m�r�I;7����̦���ç���ïCӗ!��\_@�1ԍ������jN̂�ޫW�]�Y�K�s���.:-Dh�X|M�D(��/Ř��mV�ݾHt�u��1h�U٣�J=���we^�m��ծ�;�(:*�-�$`�v�ȏz�$ǥ{����y׆�0ʸ��3�V�a�.v9��S��\�n�����2���'HN��"�Y���5�ܖ���9����Ge�+�����7��p�+�L��k�m�١`�X�[��Ǒ�8櫌M�W`�5��\6�%�C�n>��T�V���3 I�{gQ�����$�T3|fd��-}/;2F��m�g���%�'
���X̉��T���j��<&���̉'>x^�R�Ga難T��G
�ɘ��f%�͇|���sz�eY7������@�wG�NLE5v��ʴ��r[�'�b	��f����w�4u��!>�.I�
��0�]�w˻[�1�#J��ضsz�ƅ�|����s�`Ǧ� r��k���+'W^��& <&���6��b�Ʉ2��Ǵ��.��mhnJC9>ʘ��0�"��=���s�KVEwL�-�oGu79�F�o��C]��˚��P�}Y�]В�ڠ+i�,:IF����o^����0���@E�y�K�o���������|M����O1*骳���,uǂ��a�n��L�I+�I$�I$�I$�I$�wwp�W)U��Þt&�����tm�R����_նQ�{}ӗ�d�"��Cv��Çn�P���P�U�\�;1�ք�3�{|a��.���_ڵRNs�(lV�y|[����7���ͅO�ft<�U�ֻ�O���
�qq(5g�6*{DԴ�톪NxR�9~�g�H��1ˌչ�y��?�*��ϖ-�Pl�0��O�K��vZF��B�J�s�Ѵ�m�9�e�5X X6�s�ì�x�X��huf�u�
�ܻ�B9��&ե�3�^2r�&��KZBCl-MkD���GKr���m��jm^B8�Ͳ%d�
��%u�s+ՋެEP��S�ky$��0j�����Ro��?q�����?{�����}_��ߝ��~~����p�[Y�f����D�Um�l
&��ך��[
�x�����6�p���2�̰'F.��t5WujG|���4���/�W+55K.�:���Ôu�����9��Ar2�_e@#X�c��4;�Aw�rZ�̥�>,���ocd�滑9k�
}!��ˎ�Z�9>�Ta�j�t�Zܭxy�$��o�Z�n���Y�F�'I:��]{�Z�%��X&�:�J�.���r$c���^LC��vwɼ.�vE�VoacS5��0�
��.���|L��h5�\z���dli��I�qt�G��֔M�3F�����*��Z��k]�[��"r�3/`Q��κ�5y4���G5mr��j=yI�ɢj�d��ݛ�&<��
��Ӛ��"��B�!Vy���j�6꩑��^jJ�qY̬����*�V�:&���U����o�ռg[�;r>u݊,��6q$�X=,̬y���vHnnÔ������݄[\w,r�@����e��z3�wW:�LWC.��E:�FK��xL]Pq�H��NΓD#���=���$|/{�[�Ci�D��lE�dW�L��$�|"ƾ�f��ݣ��Sv
�(L�ۺ$�v@�[{�N\�'%֠�2��R�1|�S����\/K��v�C�C.e�Aj��SЪ[ݰ����tdoD�s�V��[l.���6������s����ϐ�y�Ο:.��,�x8;�W;�F�r���>J� #��*Oqp�f ����G�]�
ߓ�'u��\ƹ��u�*S��UyO]�\��Ź@�"��7��k�J��:�V��NR�ЏEƲ��k�u�k�7����W8ե�E��a��7.tW8�]+��z�ae�	hn��͞�;�em���ͽ'��;���g�G>"ES��s��]wc���9H�V�M2�,0�h�����*�]`��A��}oe�K��/�;erz7�R�L���j���z�(��{N���r��{	��wtݚ.^)���ެ0X�5�T�v*�X��6q���¶6:�b�O��P��o�`����W�PF��vku��֪Xʄ�[��i�4rxs�Ag!�3��N�܂�i8��J�IQ6�VGN��a��ZoNn�yl�Z8�k6>�^b���VWS��f���'����f=<��c����S�#[W�^SH�D�ا۔fkkq�o2h����{���b�	�.7���8��K����)�CM90�3	ǰ�rՙ�*����M�n�u�r&=�I
�N���.���h	��C�WvC��C�K[�Ax����+[��a@NK%�9�f�����w�㴾5���幒n���˱�~�Lų�*k�t��2~�B����Uu�L��2�}}˝����.Hdzfm1�u�H�<�e�=�uۤ�!�U��- �3����|���[J��?[����\���te��z��$?+�>����i_�Kۦ�7�L�"����rƍ�"���:e�櫈���P]؆�c����}O5�YZ���"���r�=̟���:еG���P��]���]K=;0Y�}0��1w'n��9��ʼ!e�̆��2������'�ۋ{xm|$P�N�l],7�7 ��:&�u}9�ߦ�fL��nf*j�d�]$�
f�êo-7��_2s~��X��j�uҬ6 WtK_;
�R٢�����Z���w>~�ūU�\y6% �����Wc14��9QS�}�`�|ᨫ���gkX��s��_	�|W��1`�U�O?��{W��v_a����n�ۣ8%�
����v��t�ڤ�s���f��]Go��](�g=��)�Wc�h'r��}�5����<3u�%=�O�J���,��ԩ �X�F!�ӈt� N7���:� �pVJ�p>/T�m�M��ݷ.sx��u���sx�h[�x��}yE�N�N��2k���B���
`���*`�C\�yQ p�\���U,�ay_L��4}�
��J�����_/�����������m�s�h�v}@�b�UJ�.�^h�0�E�paw@�N��r�v��E���M���Ld���҃��5s}��n* �o����r��^a�8�+��ͱU�6�7.f�v�_}RE2κLN��΢D�r봾�ՠh�*��vRS[��V�Ue�wf�t����xv��c�f��2B���ŕX�	*�k�7V���XQ�%U��hŷ�t��s	x��@����5�w��,�U�f��'5����	�f����׽�zb����]+��l�5K��Ֆ|M���>ϐ:�n�����w���v�����k�q鿞��aa�����1Ҳ�7��*�EbtǉC;�˘�^SXx��^<̿����Qr�̛1�Vħ}%����)Z�i4���me|	[�N���6*h}�"&����sI�1^��u�b�{U���R�7�_;�is5��7YB�WÉ�`e�I��7���T�:p}z��ॢ<Z̖f�T��p���weYfvf�"��L=�ф�*޸om���e��v��w��V�d	[�W[ι�J�hEE�I����9|2�W����LUc��Jz�a4,eN5"18w5fu�e7.�r�y3n�{�ǔ8��A�\���k��b���	u5D��|5�	�X�Z��wu��W.{b;� Z��_@����� �o���:�U�^��]B%��i���$��ֈ�8IE�_U��Y�CU֎d��Z�� V��^��}��[��2j�w�SM�!�AFv9�fZ�I�7u����H�����V�ߦ��k�/�Y�-��8�ȸEbd�n�M����-����c5+c6��r�$jCX�6.S*�Oꝰ��pS����ߥ���K�%���Z���u�7�%"�DM���ܗ�sb�+�����-�se\��K���U�N��@��!̍r尣m+)�{�>R�a8;Ejh�&�� �۳&V��GpP�ܣ̭{wY��8�VE�H�sR �׋���j����Ȳ<�}�d
��?j5����Tz�A��tVH��i�I-ƭc=�E"�ᙻڔ�n��V��̨�QfV��׆ni��+��ʣ!ؘ��^;H]�L��2�W��Z�J�˷��ݕs��{ΰ�oM�vX�8nt�1YxKr�p����SY��5N�	�[��m��y� �P�}]�)nT�55O���F�T#IOk7�0oh�A��tm�;ΗH���jo�	�TV�*��o�n�T�'�4Fݚs
I�ڰ��ɪ�����Ѫz� ~��� �����[_z��>_^g�~n�����|RL�2Fc���!#l�r�H"CF'@~a G�ȱb�`��E��)8��1CB�8AM&b`O�mY�k��S���3P*&�!��1-�Ƞ�q�{e�gi�iJ��ؼwf]��A�Z%��(���t���ƕX����.�L���\����,U`����,0�&}�� íVM�
�u�s�	��w2V>%f�n�e�H��-�{rqF�,F�5�I����&�(c�P�η;����ĖX�S^�?d�JΪ{�� �S�Sn�l�Y{:u1�lԬ�δ�i:h��Y�"㼉<�Sw�d�6WGj>X 'v���;�o��z�6�[x��o�j�-���W�U�k�oZ�[�;^�E�h�>����.J�M�M$�zܘ��q۱T[$�i|�vܼ����sU$d��Jm�	7������S2)�F󮵋Q�h�`���ve�6(�2�Q�\�D�m&�*��P�)1TZ5ɥ�e�V�b�Uʍ�]���Q�V5�4VR�a)�v��o�ח�F��ܢ4QfJk	��QL�bL��;���7���[��^+�b���:|������"ݘɑ��23��&�c�ܢ�
u�W�gv�����u��:�e���r�����,�J\��%��
7f�� �h���ӡ�N�Zc��=sF�7�=ZǓ�[3�������o��I�1y��ӄ�{�����kK�����4�x��&7�����Ap�F��>rP=�)������)�"n��P����sڳ����-?I�u<�t����J���ͻsa��S�?L�
��;�*�[� |N�ׇ���G�q+��ұU��/�[tvd��Ʋ���=��U�4Nת{E�g���+���Vѡ�P�X�^�Te�ܔ��<>�+y=���5�T͜�ة&�uʈ���U�¿'�#F��b�j&��ۍR���'<wv��q��3���r���]��7�z�n�����j��g���i�Ǔ���.�T�����l���,���M=����v����;�v&���_�>�^��+�|�V���_�[籮��}T�E{\��)nG=�]��w�T^�eUȤ<قF�����}��'B�����l�Uwz&��;-��n<۫"CR���t�p�4v�[��`������1����� յ�Goi@�J�6�\�mKCE��f��ʪn�L��G}3�X�iBix�wF�\��Q�K��8�}||�e�~�4��y����X��&���7����y=��i@=�;�7Ǜoژ+�Ng�l�Sg��鍃�o����<�����v�t&
������;��"z=��R9+�ym�:�gl���j������7�۝}C�MN�(5�=���o`uٹ�.����`��{k{D��>`e���6Z�����'�*U��櫽��v��9�t�[�k��͹�[|�vm���'�V����MJ�>�[kg��\%��՝���_:^�z����ߚt�}�-]/Vk�j���MN󯻘lu�]N��s����62��h�c�f����7a�S�K���H�TN�S�{U�ۓV!*b-���é��A��^�5���p�н��/1O�Jx���ѭx��jk��[��Cyz��a���*)�S���?zC�}v�E����v���cױ"����}�'�ڙ��ë�N�s>�#���s����`�{q�I�*��6r���P�v-e�}�|�.��&�=sb������/�>��pQ�6�D��)j��L55'�J��d�{�'/z�8�싸���h����O9�ߛ�I�k�V��WCw�~�������P�t�wo1OV{(�|��o�:�i�ϞUS��o³�|䋶�z��~�)��&D�l�/O>[��~5ew��u���jy/��%���}�w�|�7l�d�_��H�@�y�U��>2A�k"є�����Nɼ-/���6�z����X���Uٹ�fy?E���>�Y#G���'P#�'�GR�6'`���ŭwu�奇z;՗�񐇧�ڿ`�b�+�9b��5�i����3�{�; �g-�o#�g������H��C��f��};^���KPӽ̜7J�s����'�L��)��)&�^i%2ϧ�&�y�����|�4����]��^��F�9����y�|���{&�%�����9H�|sQ��!yS�I�'�t�?-j�G���Y<�f�rq���,�t��;�`��A-W
9t����MS���s�mԤ�k<�j��yY�R�̹g�g�ck��.�n;M��E��{2�Wx�o�J�>��A���Cw<J�=Cw�=�`|�4���Z��Uҧ�a��|���vf#�LTq�w<���>[<D�^���BS��P�����몞�T�%!�sɘv������㆐�ɐ�]<*�<^�m�(����Z�����)Ը��=���flfv�5n�o�]ѡ�{�r[���U�9���l'7\���P����R�9�kMg���w���{�^Fւ:D6�1wC�q���6kw���O�ㆰ�oA}�8c襷�3l��':��Z�j���ڞI��׹c��]�ojJ;�rX�3]�V�r���P1{�>��b��V�_�����fY��]Vytƚ��ꈌe��
����_I��#<(���s6L��.��u� �~g޺���=��S���Wv�љ��'�c�{|(���Jr������uUm���Onb���EM�6=�y�}���gA��~��^�tʝ2��I���7���o8N<�%f�`�E����U�k�.�t�H;�+��߳��}΂�ӥ�#CkX˗���DG�:���B��ᣫS��:Z\u_!�k{5	Kt���gm��|tٱA"�*:���n�o*،�x�{E�b.��������ю��gsnC�l���Vͅ����Qe��gO�۝��z#��|~)�UG�;�{��[�ws���ۉR0s��m�������<�~�ձ�f����͝�����_��W9���b�Rd�A=�f�����Q�K3&0�E�ar��R}��Mv4�Ӻ�k����S�I�_$��W��;��-�o�{
�ރU�zR�'.�Qh<�_s�K��Wg�9b��3�"��I�]*���P�s|�

����R�MK�=��M���`�VQA��Z��#�u��)��=cL�g5ۺ�M���OT��tt�Yo"��]��(8�y���gPV���LN�M�!����w0�2���g��>�Z�>�.ך~�1b�P�67,�u�Wz��O����y��Q{��4�b��;޾��Ǿ�
w��gJ���L\���N^�V>p̅n͏��g���Y��R�|/z��d�,���ƹ~���Sqy�~��^Ͷ��_����l����>�]>�^��!��O��o����BD����y�2 <o��𳑖���5{�GK��$����w7�j��g�mm��$w6���Y�ra����m����+d�ك�0�o͊��e�*P�yaa�v�����Jo�,mG�JVնw�#j�_.	7&����׌��]\�͹b�p-��x��̐�`�M��Ȭ�w�t�7w;y�Q�s���J�+8d�yxFGdH5�!6T��Ld�;����ќç�:��p]���IV���uܾ�p�]��K0"-��3k���kh	p��ݐn#�c��$��	J���Y�.�Wu��֚���/Reȴ�Z'L�����f��:����U\t�p�A���Ɉ�������M�9��-��2���:��WY���1�v
ƫ�A�ǋo��3�H����BnkyZ`W#Θ�f�t�*ŷ9����ڈ�lO���0I�F*���l,)�E��r�j�[�R�h����8��,Z�ز�A�������	kd��7��<��f�$��wI�D�L\�t�*Sv8�C!���Q�9��צU�p�;RK��vR�8�5D�ʐ��R֎���>�d]gM�[�����{�Ƴ;�v�X��Q�����"��G{���]6���R�^BI��C�����R���}4��;��o�=��I�+�\zې�|V�J�p�t��cx�������p�;IS���<[3^*|�Jx�����;2]\���<�����|�y���]��ߚɵ���/U�o��׍\��F����ܽz�K���i5�^-��rK4-C�w����Twu���t�\�c^�b�:��[�r�]v�l��3Y/^+�n\����x�ʻ���r<��|	 W�Vj�қc*cG{�����Ūg'�Z�%��Vj/'��ڃLe��b�ut�8V1���soÓt].)�w�m�a���b��k�����;Y5t����u΂�\onlʇ�}�����Ĵ����Q����w���罵fY�ө�s0X�ED�P�α�
Esoj�ƌ�Ka���8z[slE
9�� ��ʹ�����]���KZe�c�T��*,^�wQ�Tzy8x�,ϳv�.�VB�Fٝ��֍�z����z��P���N��V^��vV������%>K�bws'���I���@��8���-r�Z^�ޝ�0��6;R�m���[ħ����B��A�x5ϕq��8�����W�F}��;���A����hޤ�y�`�K��c���[�o�{�������j�T�@̽>�l��GO�u���1�7�M/���w:E^��9�'�V��).L�G���R��]j{k
ia�mjr보�`N<����kw����)%�����LtOc���/�-���V*��׋����.j49�N.�<1K7{�����#&f���h��DTh3��LP�ޠ��v^���������`��ݚ�� W�
�6�~��/)�von�ɘ͉�c���5wFm��C����o޾Ol����{�b�{̧F~�A@X���v+��6m��̍�hH5��7�+�n4����~���y�����B�t��&'{k�:�-�!���]�#d�ɕ%��a��ɽÖoߟ���kl�8��هU}]u���qt#_�ᥖ���e)�X�:����xK��x�ɮ������y��vq���n�֪�eۏ6��i����4��gVd��R|1��u�}�"���-�"�z��h��޹�u�΋�;r(�k7�s��ˆv��K�ؤ�
;�R��ez���<���λ�TDDE��h)�^�����=xx{�6��jx@��O�1zzG=�����7���c�6":���k�v�z"���L^g�D�5��g�y��l�J�	���&U�����۷b�%Ou�L��\nYW7�G��a���q�̋�wL)��|�%�����b��U����4��xE��~	[C�ڈ�}Ȝ!�}���XG'��&+��;5;δ�.��]j���J�K���L�QQ<�d���Y@WJz�g���믖� ��}�GѮr5~��I��י����S����V^/ �S���G���E��z��P����~
x\<9ܱǐZ�s-�J��"Sx~�{ި��U�ɔz��3-U;�%�o�,Y�3�k�����ʦ��`�hZ�%3���}Q�O�y�y�D,�����32y����ʙZ �o�S���\O�=���fM��3׏��v��s���؂��"oT�˚�����q)6^?���Q������y���nd��:�]M`g�ny��t��*���=>�H��m�ƞ'�c�n���g�2s�c�QYN��=&^(��_�?��
a�K�H����sSn~z���!"�y��~�bŞ��rH�<��f�k�Y>���yW�h�u|�;c�E1���O�dTT�lK��x��k�����
L>��
����A���U��']�,�y��Y�/,l�0�Ɂ��$G@����.����������h�dZ��ܱ��)�lGdY��Uŋ��7S��yUU�!����q�.2E�XU�-~��ۦ��>�'od��)i�u�Ǩ�9�M��;�G�1,n��v�O�n�-��K�Ψ��YsN?UHxz�8�Y�����T%��蜚4�5Oʯ_�_V<gH�����W�7���h��t����#-YAůn��W��E�0[^Y]I�'��n�ې���	��h�g����ݿ&�>��7�%�i���e<��]�_}�W�b�-5g{{���N5���Ffέ\����d�52�^F�K���Es�kɢ��"�=����'tL���5S����9�ӽ��=�k�V~�}h�*��_���BmsX�.��_vO4[�ts�v���ZA�_([�[�����mE�.�lDeћ������F<��s���Z�'��]���(��O_Lչn,�3���%���aǄ=���3M7�=���EoC3�c����b�9j�x�_�T̲�Z���R����:d���OT�a8%zq��KdGU�S�qf�JR,��h��r�B��|< �h�Wo�.k���3*!L)�h����g����̶K�\�����j�y�*C��q��E:l)�0U�(����Z!KB�̼׮��p�m���XګO�ٌК0�m�;��(s>��[j^7�Ouػ�xw˝�V�f�ǆ�T�ʇ����<;d9��n��=��Uea����e�ڃ����1�͊��B�za�,����Cv�3���b�C�޾�ctD�nK���:�י���<5��P3���������GP�����T>�{[��U3y�z|�����Y�$L����[ڄ��qlv�q&�G�_��vum��N�����"V'�����W=�}/�n9��h>|JJ�8B��x��p��ي���DvV;.S�.C�u��ɦ�j�q�Q�:�O���}a]n�~��=sҿGV!�b����׻^�{U�&S#F��|�R='Y���n	[���K�lS��@�W��a.R�,�+*Z�]�u1P�U�K">��G�6�/{���u� =LT*0�:۝�46[b�;-��Rח2[|��i�n�'��$�T��8$�	Iٿ��-`��č<f�����ҔM4Ї�he\�P������>��
O����xo�uZl���}Օz���Uu���͞��sS�7b�N��'��U�" M���ɨ˥���]0}���=
圝2gQ��1�v������/A�}%��U>F��7��+M�� ;����7?Lઋ�z�^��
��5�Iy������A��@���uC%�v21t3�u�M[@��c���@B��⳺0cS�^)�n��5��7m:���o�g���Q�A��mHb0&X��>���N0�и���Q���E�����@��I��85^ɮQ�-mpH�m�B��xդ��ŭ�+�v��Č*���]���gk��[�4�����N%��ԭ}�,�v7N�f��/��]5�k]j���\�W��|�L���u!$1a�8��Z�aN����.��:]Nl뵥�n�N�\AҮ�5�SP�Y)���˦b4v<+�y�^��o�]$�g�T�tM䉳]awm�
�\L��zڛ��V����4���wKJ�	n�k�ҝ�	Ԅ1�R�Xv�����L瀛sAz�p����B�d2+[IWZM��X��l�VWe�G�m�X�'mBu���"p aoV��YG�n��j�>���A�c)���(��W^��A3�azF�,I�bDSM�Z,��"�)|� ����C�w��~v�'��}Y��cr��ҥ0�:����oUä�ZJ����Y�H�������] ����G^�A㏚�V��H�݋��T���Ȓ��x��Yw���uQ��u�^�aܗ.iB�z&��e�[�E݂.4��L�rV��Co_t��ЛL�Mu�-f�w�)��(�e�l��D�'*8U�Y�B"���k�m�1����b-l`W�T��*q��NC�BeJh����f�ծu+Zh�m�-n�W��m�S��k�V���#��a"���4��g˴�dZ���l͊p5�\7�dh�C�w�:�p?��5mFP�-}w,����K}6�$��_���7$�W��|�U�Dl&�wb�<k�	,c<�\�ۚ��qF���)�F䗋F�|�+׾:�K�)�/�u�=Q�W6�	�\�^(�'��'�����;�	��"�A\����Cu挙$�:��;s�"�O��m+Q�4"�1�����D��g��t�s�����do�f�K�=�x��3R����ɟ��Ņ�}	�zr��w�]�OѲ�L�\6��퇆���M���v��F�B�|��@�}���}3L�9�y[�-�^�<(�$wk�U����W�\�-���k�k�ك��W����g����}��zXO'�m���Q�w�"�}v��\k��q��z�ߤ�ث�2�O����~{����aI��G,�a��5�0;��և=�;�C<�,����S���n��]�l��o ׾s㾢�i2]F7���.D�64	���6duV�Ӝx�kQ��]>�i�b�����Õ��̧��O�JJ4�d��� {��Ws�ܕ���_�0������͏9��������? �9�W�{º��ܛ�!��3�՛��b*bqm�Y-�V�Y�]h�6t<�T7]�[������nzǁQ�o�13���ݧ�SQ�M�ݱ�*��Bþ�΅ �D���*ꋌ��S1���H	�g�٬#��vb�cb��v��~�l�7���'�b�w��^@/uQ�.��⫆ЩP�aq�C����j-����
�J���׳��Ú&��v��ڠc7���I�[7��L:���GYbra=��+���xxxd�%p�ͽ#9�-�ճ��P���T9��;'#-�N�����{�Y!�6�h�����@�ra��M�יR�7[/y�xL8�	�z�E`��)����	��ݭB�r�ڜ&��ʨ�I�I|�R�WP���qP��e��*��GOR�����廰�
��+�Ũ=��U���k~5�R7' ���&ʻC������nu�Όkhw��i��畲W[h���Y13�3�~uءjy�_�nzQ8�;��{{/��ycX�
��s�v���w�-�!���i�������K%��9�\z�UK�5]ZX��xx{��r�[`[4��}8շ�q�_f3�q��\��圚Ly,u����?�����@h�O�J�c�Av�]�d
6�Ԏ���̖�T�(�ޘ;F~>��E�� ��o��0�=\�\�lfG����q�FLF��ave!$=�8a��s�E[N�ƕzI��2�oq9f�<���*�8��u��mJ���̯O4[0L�F�
�"Q5����8���J�٘��z^��&Y��-@���1������o�k��iH�p�~&�:/x=�3�(#w	i�/�nQy�n�ܯ���;�!D[��ݺ]b�4|�J,�"���ΐXt5�����z���"]��!C�FϾ�h��jh��o=2{�Y�d+A徜rv7**3�JiC�x�mQq�:IcT\N�*yl���Vt���G2��vܲp���[�4���m{���ds�B�����QWt���Lm�YxB�ܹ܌����D(��}�S�O���������՗Oj%�$Z��騽�P(UԊ�W8����u����a�|��SE4�܁/;r�\ ������:�Ɏ�������y�v�<�m��NDu��2�/1SWh��Sm�|70��nW0�tR��ˤ�)��n;�L3V�tHo�x2�-����兀�l�����Bm��M�Ch6���2��v�i�g��11�'��]����A���V���޶8�o�,�"�G�eR��W#��V��q�"��0&�e��]�U<ź��R��nM����΢�k+&9Kt6L�ȋ�h
XWjy2���fW�U.�6��˨�q�|>��u�k��;Uξ���mo�M6���q ���Ҏy3��P6f�)����ݔ
��V��P����
#rGD>������h���n�n)a�x��%��}�^Y�o�-��������̴��Te���
(1��?��t�^�|��U��_0��k5"9�N�*U�mY���p:���鼠����ȧ!�`�Tc��><������B)o��qvF���@K�[�됉������Gb;`�P*E���[��|�^q���=����j�{+q�\��m����w�ɎP|'X8���=��;���v�=�8�93��Z����c�ץ��^nd���e�s���\�'r�Z�o0^t];50?���R*���{��w���������v�E�.���roY2����d+�@��ܬ}h�=WWu��}��҆��������`�ho���m5�W��'7�7ڥ�"��~_����� g�����w�}V>k�/���i���Ա�S)��hy<�c!��_n�"3�m��I�_��~��ra��ߘ��y�1MW;;�wh>�2�ɠ��]m쾢�j�X�H�s�S�4c1.�����+������Ȑ!6�3$��ڴ��b�3C���*s�^�9&3��L�W�^Etu1�ΛU4t�vb_���,h�v�͡��g8]��~�3O!�4���koK�4E`��s�e��v�T�*b�'}\W��.'�b��O�����UV[횱�g��=&����_i�������3���G.[,D�.d��sF�y�x�\y�S'wE��a[R��g��l����ŬK�u���9;���If�_�Dٿؑ���zk�5�|d"��N0�j8e�����|�%X���(t�����Vޫ� b�����-���(���4��7O�e��'�bJ<�d����F�[�#��q0�����W	�]V+3Z���ϖ,@'=BkI�e�ƥ�sԂZ�����yt�J$�:�X1��:�	�w�tr���^��w�eݏ�Z�+f� C����e����?6����t�9��k�v�̟M=M���M��dnۗl
{qZ/Y|ا�4P��mY{w]=9B#3zsq���`�Z1��>���Og�������zatpx<I�cd�?�w������~U{��g�!��B֚뱇#��ga�0�n�s�E��j���P��Ϟ�²�y]()+��:aKN�g��s��Zw��L׆e��T��5��:Ά��EM����o�#0�O�葂xX�r��S:эA�(�6weѸ��f�w1���e�"Rp�mK�v������X�:��!��-�
��4��i�AdÌ�䥓���\���%fJ��8*���z�t������*Rr��N,�O� ��ּ���+<0��{}%���!
��S�M�R�p��z]e]�J{_h'N���1ui]������n��c�w�뻫b�'�j)�\�O�Q��?+m+���Eav�ޣ�MNG0��:��@P�%�\�{�����% ���u�]��t�����B�唃�d�+Z�RՓo~%���tM�x������{�5WӚz&k�NKɄ�;��Aay�g�z�K���D0��Zc]��0�wS���n��˵����۵�����VȷPEv.��ǖ��@���9��4⦣�	"-U㷸��
��ܩ�Y,=�N5ֺ�f|��Ъ���:������SyZ�J�MPs3�^ң�K�w�)�us7'T)��%�N�'���}�zv����ki0t���A)�xIi�(,U��صv֭p��@chM����e��f�*q1p�ww�f��\�: �Q�V_=\:�����wo�+ӷ(�U&(���Q�X'�|��n��G.TY��#E"�W+���e�`����D��4V"#\�g���2ČMx�%(I��I�x�v�__͊�q�5�K�䌤�3�21$����u��A�-&�p�	$���ukXѹ��w:��R�G�\z'>����vn/�>.]���_�s��U�щ ���mŀ��}Y}�՝�����,r�m�~�?8�exJ��ߩ ����zk����*��f�nV�wքI��ߕJ�W���\Gx�8��x̄��8}N�<m�V��C�U��so˶���2ƅ죂��>�=��C��ED?~��g�w����k>ґ+;{��s��T����D�����tOB�*x���k����:��sGn���s�b��?�wUЭ4<׏l7̣
H�{+Z�[���!�qJ��dY*R�>�nix4���n��:��3��Q�`�Yڦg��g.�����L�齼�,�[&��ݪvJ��[w�"����p=<��"��O��j᭥���F�0yUsGM�s��s(mY�\�a��aR��WqU�G.�����.���bq����xR�ޙ�����Y���G���m~z�Vޡ��/�=\���iS\����4N��V��[��6zqY'����ޕɂ9��ͪ��yH��?�Ғ�ɐ�9��_e���1��ϙ�Z����~9���Y�=t��]�{A;���E)��OLT�tr[��L6��?8FzA�%���6U�Głַ��N�C�Jk&��tQ#&�G�M��%7i�eq�n�3�/�p	����7?���3>��N�,BC̵7[�x�9��g�wx���[pi�-�c	����ö:{�ތ���Ҧ�5�M>oNTm� 7hW=QM=�>�GUM�v���W!ȓ0�Cz�{�ku�c��ŏ����a�0}��A\	.��6��K�~*K�b�\�O"�Q���r�Y���tR����ڣ���ߣ&�
��~�����QN���o��	�S�ĩ�wn̸�n�B3m��K�<䬆F�OLʡ2����<퉣*g�	{�P�Ɵ%������J����3I5\;�� k�[y�(ؗ��ze�+��j�̥��2���P�rjS�n5R���T�ڭԲ��=!E�-��ޙ��JAT�Ȏ޹��2$j��Av�zx�6S�V�;����,Q���o%�wSl�WGn#oe֎���pc'%��R��a�չ/s�@�Yf�HzB�����9�T�|����م7���שf���/���?;��qN��Gs��n�B���y����J{����2���Ǫ�K��e�_���Cz�ۚ��wt�������Yo������%��W��U������kU(�2Y�˱����^�/��}���Ub{׮�X��5"�ZF(�T�2�Z�w�ES�{(��ffLYis�N	��vέ���h[&u�?e7m�S�%0i��@�v��Eu��v�Ph%�J��n�m���5-WhZb��l����%'�$�ޏ�_���<�[F�.-j]�wS���m1R+�����䚋q�~UЩ�i��"��/[f�n���5�Gw����H)��9�f���#o|����}Oߋ�'6k�?o�DH��>�Y�c�����]�淴�6�
�����vn�-����von��Vļ�(�w�����¿�=�΅`����Zޘ�\���˶���)Sݼc�Ƽy�K�tDw�����of��*�]+=��瘫�k�F�"��Q��g�k���s�)����G����������@���C«���^�vAw/YV�<�o2D��m�s�M{�#wm�GG4�6\i;�����;�d�/6`׳5�bo���������{�,�Na�Of���j��!Ⱎ��q�p�*��,U=��%����d=z�·*ի$��in�ޥ����|2��xY�Ʀ�.�%�vollK"�}'JZ�"�$�M��\�Yof`㸺��p.Ve(�F�[���4K�}[#6��˺�����'9uO����E�T�(1�JO�<���7�� T�D+�-]e'�����{�ݴ�
qa��TVڭ�G߰����V#s�=v���y��_��\���xg��B����3�մ�[�Rx�3[�j�0Q�+-�[�L'T���Үm�*�M'�{����CӪPd�`���ץswqC��n��/��v����_��";��7[��|�	F��*�lل�GU�W^��8���c������2�N��n�}��
?�U�L}�=Xb�*��UB$>�������?-��P�y9}pr/'��HU�Ψt̺-�J92K��V�#���0�51���t�ϳ0�t)o���C^o<��*����z���Gd�gFr�S��-f:����I@�qԌ[U���i�mv����W�-U���n��7���z����ȼ떔9_Ӳ�)G��W~�*�~�7�~�wl��J��uT���;"YWCN�ɭ��=�){o���)�՜�m�!��Xu���];���밽yL_L���]�pۢ���{�u�ul�L�۽�GG#�ފ���޻�����?�:�s�1�d��cM��-{ݩ�⢳����#�7�UQ��[5n��ѵS��|�*u�"m��WD�������Ům���jC���*2�;О���Xvب4L0[�4f)p��;�wz�т����9qw��'�������f-�]�G�9�;9Wl�qb2�Vnn!�,���,�h�V�`����zPU|�za^���a�ʷ>�f^��D�4;ړn����!�uW��*�x��n��s/H=��O���u��۷�3��RgtT��M���"d^z�U@�;9�KxL�`n��h����s�seƘ��ڒ��D�e�.�mo�wPa��Y����8��a���<B�78�R`_��Jn��㲧�y'�S����c���{�O4v�l!Q6q�1P�Ս�ǻ�+u�3��F��kg��b�':V�U������l�\�̢�Ƕ�V�$c�Y޾;�E��zt�n�g_�	�μ�mV�>�͆kE΀�Q���k�{��ڟ
8�os���/��r������C�	Ą`�ۄ�2#XK�r(�X*��𿇨o�_m���S��)&#�"��m��^h�Wl�v�M�H�GT�qK�Y�[4�i��\H�"��t;lb�[IyX8gSE@ʝ�F���"���uZs���8�Ýs�e�����U�(��f�(��tTAi��tˏ8�o2�t:��/z���mv�A�1�a�YW]���G;���:᜖���]�^�P+�zۖ4h�XL��S���W�}N��o{�8IC9���u	�ͫ�q�t(���(��I�Yʸ�Al�6��-�Tj�vy��+��w�5��.:*s��(.��ͨ���T1�]������Tw�q�f}���Yךf��W�x�]l�ga�U�X|�[��.�(�9�=�������-�O̤�lJR3�����_4q�:~���')e#Q|a��:)vUe��wKǶ�+c?nh�C��D�FX���.CP��X�W]`+l6���k�|���ckwqңN�3�9�=���ƙrSݮS�q���!�7��]�,U��.*B� z�В�/���6E�[�F�2J,��}���SN��)r���"��n>}�ɠ�[�@*j�T�s�����"qŎ�5u��Gp� �ݏ4�]֔�W6�;�S����%"sK<�j_+0I��>ޫ���*=αu��V ��F4;�ϰk,v`݀�/���ΝԤ�#�;�{�������m���<��ps���6�S�sP�r���̣�mwp�p�9sooH6(QEDj�Q�H���������μ��ϗ��>�w:`�i�R	}��(�}u�iB|뻵���$�:�]݁�Is���Lu�a�f�褂F#BL���L�c'9��^Re����Da������d`�vlb( �	$�Fb4B�iQL��ŔV~�鵮����ie�,�I�8��=��M��f~{�LN��P����!)�nD9i�;H�8�q��2��k,CJ�%?SS�J��
d�73]O]�U/{�+J��ݰRí��D�}�9�dLPh��ɻ��-u�֛n�Wds���kk��
f�V��|edu�Or��ژ�k�}��ϣ!N���n:l)�x�N�������Ī�
�Iy���zx���'{ycٜSe��L'��mr1�vjo:�边`5�`�g}�������/�Q`։��KW]��|.um��mn���)q�c��-�D�
�Y|�	�޲�c����&!>C�ĮCa/T����K�D�le�?���4����G���2.8ԅ+�3K�=�bC���E�3M]#���lDYݝ��h�,�x��ꞣ,�1����,�9ۀ����j��y�Z����ǃ�<m��Ϭ#�ʘ����w��Ãx��N�T̙��9�^����öZp`�~��&�d_�0O��c�=_N�쾜��u,�%@�k!�2_����	�QSʲvs�3���sQwq���2"�ヨ��N�Q�(�st�^k.m��} ��R{�;�
)QA�z��Sl���+�RG8p��WG��Z���O6��3w��_9ٖ�]�����(������O�ߞ��_)x�N*�Y�����݉䰓���k�e���|��y��{;�6�Q�T��d%�b��,қ�������{����F�Mv��.��>pZ5�[������i�Z��k���Dg
��&x��i�a{��'6v�Lc�釭�e]���W�.�0��S-r��N��뵺���+o:�~c�|6�ý��c���>}����~>�
����;��M�-�v��~F׈d_�noJ�}~�Y���KOζ�ǩP�>1n��]o���T˥6��Dv�������j�E���d�D��:�mT~7X��ƫ�$]|V���_.�:Yk�g3�}����.��З���V�1
�["�:4t�+���(�G/��j��d��z٫��<�1I�gf��խ3.�ΆO ���";�I�!��h"m4Ȫ0����SwC�&m�c������'8��\�ؖ,������*v�*떖���j��@�ɀ}�˵����#ى�\�*��ʶ�'3`H�TS\.v�l���["r=�����C�B����;Ce�P4Ӂ|���Sϟ�?g9y]�l�j�Uu��C�YV��W��d���F��AX�6�u�O����v��b�h���<#�f*�#��!����/��j7���ڻ���ӱ�W��b'��UR���uх�T���h�����������d���G<��%�l�!���oS�?Q��a�u5�v{��n4�F��omF`�*3��x��o"z���vh�_�po�J�ly�Ւ�9\�
��t=�1��+ۼk��C��ʝ�t����hն8Ұ��؏�?H+�/�T3�WTz�̋�N<�a�Q��Q����A>�~a��vٻ9Y�N)�x�$�~����t��zt�v�bĪ���u�;����hJt�5�L��V��U[n���N\����ܺP��ٖ�A-�]��o�I�M~����P�W�1������u�}=���)��9�r޺�BVT3������3!n	��@-P������-�g-���3�k0.�q����������k�C|k�U;cqD��ƞ%������Q���x�L�(���*�ۙåح@���
��A�J|��w#g��d�/�t��k��n����%nwNYvǿnl�_�]c�)��x(&��ՌSͱ:���Abh_��ߢ��͔��J�@�[��*ڥ�θ��a�W��<u�e�f���Ӑ�v{Z������W�2^���ꢝ����y��f�S����7¤D0��j����/zVyŅ��S�
g|݊f/Ъ���u�mV��i�Cac�v��n�9��/��nH�ז�?m\H>��g�6����Zx,I��n��#{-Bia�{�5�	ڨ`!n6�̳�$���m9����>��}u�yvq��c�Wsj��S��h���YU��9���?y��s6�D>�ED5��Imu����B~X&�s�h'�dҍ�:^6���Tk�Nfm�|���Czxr��m�{.Z̸[1�-��}H�gs�����ӹT�կ�Q���2v�:3/>���|���I����8��|w��՜X����'�H��;�g�����I|mގ;9s��Z��n��@N�Y�	�Z��]Pz��9���Ҝ�T�����zt�N���ެ�����\\DM\��9,����N�}�
�n��l����p�meHX[��UY�E�o�#^��z��{�R���T�:z��ȷ�V� X9n�#�̦�1}®i�Jy��z:Ȱ�Y��T�kt�90�!�
����j���>�_s�#�3�qQ�j��9MN�[(�� �MY��s7U���톒���6�swϡ]�{��{���b7�f��^}C��ֹ���ؖA���7��f����/��O0e��JҁAϷ�ڑR��;���oeX�Q���4쩳�P�w��l�uΙ�T*ԬS�f��qw�䞄:0���ebs0?^@{{6�ۼ�}���۹X���6Nk9i����9�M>A[�������h��ot�:|X�UUR���ʩ%�����/���:Ȯ�~9#~�Sf7����N��b�t�YS��uT�Yn�Q�p�Aϸ�K2�Y�����d�B,y/�sTe�
�X�r�7���U�������`��i�gCH!�y9׾��-�+q�;Z2*�t�lc���[�(���*�|�l�и���t����}�G���{rşQ2�
c�/�C������A��{�``{2b�{��n-���L���Rў�.�������c�NW���O*����)���lyTQ��ʪf�~:I�m��}���W��j���z�i_�+���'�zf�d4^[�Ǻ�/��y^��CG�<.����Y?e-�׬���@��s������Aw�-�z�ҙ�����B֑r"������x:g^C�-P����MΆ�سKޯ���i�!3��:�耪\�w�����*L��t��kv�6n���q:/hc�Ë�v|�@;R��:��s��$�C��6⫮�]�x4jX��K8�9	��̶�y:Xtw�.����k^ジ�c�y�lݱǝ>����7ɇ��Ccx&�3h_a���q�twpFOm��!ݾZj�'���l�j9�1_e�<�C|�Ω�n�ř��M2�YuN����Gh��i�F����:�&&�-�E3 距e,�
U�H�&v��$h#4Y}������&9![���H������/�V1ٶ�)�#d3�j�c:�+�2����Q*��2r�0�9����pb1'C2�0���뎯56�R^Q�M�Yw{���hU�JZY����S���Q���C>=CY�=}#r�=8��h^%`���;�SQ�>M��:���b���M��o�'^�ʆ.NKF��v��"�e3W�ek�2��U7�s 7q�ak��}&&Q����	ٙ�Q��T���Rc� �2$����,�u�8���B�`�k��&ʩ��%�nd	�}��طٹ�a��c��#Cb4U��B�EA&ɣ%�5cHj1�-sn�`׭�h�X�cEx���hة4U	X�H� ?�ě=]<��/_�{)h��_��Ptݍ�Tzv?�>� ګ�lo��'�(���� ]^���)z�w\���J`�V��UxZ�0�pcb��;���[���T��e<v�|�d�������X@��Z�=��UX)�^�z��kk��_�3<����}"w��a���}8)Q��[���A��%ڸ/"�oJ8���(�TG�������;9.���m:��O{%������y���_m�_����5��M���+� �ک]�'��>�ˣ����*�q��DF2�N��������˗-�-n�-t.wk{G��-TziA`Ԯ+�-Ŝ:��ˆ�SD���M�g��y�������͋N��������K���
�'P��[�h�v�y3ŪڷI�\l銶ʼ�E����e�_B�Y��$�w�Z�fW�62NH���%-�V��,�{���������}]mC�V2�}�\�s]�mefL������l�D�Us���A؉���nV{���G�L^�ݮ��e,�(����?[�^�8�����b�����\���Ź})}���d���o����)U�Zt.�Y�����2H/I����*����׶��3D�����}�?[�<���=���ˤ�n��z��c~d����(�y�h�xO��3k�w1���b�M���f�wp�����{]w��l��7c�-��.z��Ƶ�S6d>��h
X��gzy�r�vV�g���A�^�3[)�g��T5����`9�3Z�.q,�E��c}�%^�!��?T��ծ`"���!�VC�m2���iM�g��M^�2��vg�h��ϖ��d&��o����4��>�g�/�zǻ�n�IOd�uokX�d@]���]�V��6��)m=)Z���\�Թ��0͛Z9Ɇ���������᪎�s�Cfu�{� @uc3��ʦ3r_F�ғv��b��@&� ���jO=����֡��6�g�/��^�@I���(<��<�VbX���߾��\l�bO�'^@y��y7=�[�z4Y�AJ����t��L����gk����E}Y~!㊤e�s�OY�S&�#5��5y1tA�Z�K6ִFҠ�eu��1{��yyz.ʘ|��H���V�
 B����,	xZY�2�eH�_�e�d%��5aњ�]\>�NL������1(��`�|�u��f*�mb�?{bb�ZaC�coET�ͪ�sAmN!�ŝ,���>����)���tL4��$\7�_��{*y�{����i8.Z�V���z����,�<K�>��.�նa���vW����{�qzP�*�p����:������u��Ϻ�����V��S˵��X#����p`�"m�����@V��{f+���/��.�9wg���<���
~��ޛ��1��T>J���;���mn�L�f�ЋR�н�6��.��u������Q]���O9;���J�������z̢:h"e�;���*j�ǜy`����ڋ?���_�	W*q6�i�?#���c�T�qyy�P1�*�s�g]��F�0�ox/[p5�r���pѵ\�T�{b:��U��=O/�,���~���*����K����{Kͼ��4HYo��F��2��N�	��K!�8��Y���mnê�����������x��Gs<LF�~�a�]�����y�&��1Ҟ�I[�|.-Bw��=F�9���~��|M��_np��u������f���ngM֙�y�w��=u;J̍h�������Fc���G'6>{N�����_�oE��M	��a��K1�����͉�ֺ��;��f*9Ϳ�P��'���s���N�mܼiyn��+fa�v坘���{��§��y:�C�o2���J��ȴw)�ee�ƃ,!�7kO:c@#˲�!YP��-\��&�1��q�qYkչo�n����}�..vda��;���R��zO�7Oa�e�|����ͷ���狇;b�e��z]���=�*�E��Я.i<3����� P�
����9y��5�Ws�6�M��Q����p�8<��ޝ�fQ�����|︳3�L��w-�	u���g�JF�nn����{�����#:�u���:a�����r�u�9�0S��h�sL�qdOodbSѳѹOmx�Tl���������ֱ��!��jЮ#[O��_e�v���5�թw���Ok��׽����+Wn?����v-�77p��O���[S��@/�,��k0j�~�s�,3�tpO+��=�3w�>R3��e�JVɾC�Pb����f�7=#��~��T��}+0g����C���ߚ�I6�kсWRJ��ڙ¬#D%�Z�����Z�����*n�7� lڬSS��G"e�&���>|2����J���.��Dv� �w~���ʽ]�?��xu�Im�q�kpEq����VJ����Q�*vgK���������g��޷���/�s�����DFݡY��u� �<����5�@�p�4GJ0v�>��e}M���~�S��[���$��я��،�oй�e���f�kک�ܕD�i�܈�����c"��y�y{x!Re �FٓfH��xڥ`�{�����&���>mᗼd��(՛pr �̹O9u!�(�6����1tJ}���(,\�d;Yp�;���l)�$��(���wm�+����X��,q���id�V�l�8���(��i��ꊝ.����<����w��(á/33|߳}���Z0M�	��S��pi��k�V[�����pt��!�
6�Z�!���o����ڗR|�^gy�(�	�ȸ�{����7*��������2��c��q�XR�����9�^�=���D�r=���ͧ�+��z��%^g6�M�:��f3n}�)�W��,��:"P��MD��DA�c��ЍFa�'�
��`?����4�C>��X1�S�VW�6��2<溫#�b��a�i'�Ƶ)];��glC�K:�n��ز���&'}�*Zn�Wv��.�Ģ!�ohG�� � Y�x'.�}-���Ε�%��yq���ؒfv<Y��ӖI7:N9+2V�6(�;@���u\��z�tl�znf
]������?�iξnS��۞8�M�����4�p-�z ����J���]��P}���)e�9�l9oZ�g.l@�0ը7����n�R�B�'�5s����h;zxꕺS76�"�V��3�_l���o��ɱ���Yԁ��'���u7���ؼ�1�2����K���ws��gj�o^:<���D�Bd� 9q9�HRP�X���3�_(�	#CP��}���z�}T��\P�v�c4[hvk��\���u@��7m��Nsmc�A:��#���T{��eE�K����C��I�wA����9�SI�U�z�\�F�Vm�,Ѩ���[�$t��8�/�et��/!��mܫqY�Q<��t3 w���E�ޞ�.ڏ'7(ۧ׎�����|e�[n��V���%�.س%������"3&��R�F�ik����@���U��c8q%��H�k�Gz�!��q��#v?L;>m�zqlI�.�=v� ���u!՚d�U]3I��R��s�+�:*`ԓsk:h᭺�Gt�������8&uM�MJ�9�o�S�{���x�uEH�^d�����	b�j�N��*66�����f�J�QA�g����Fѭ�Z�Q�RcQ�U���-��h�b�5�5y�n��64m�����^4V�	���nssWwF�«����E�x�梈�m������wx��!�8��A/a�U{�]֗�>��}jb�Z��r{�j�Oo�w�����J�*w�;~�+2��]���ΐ!KC�CǾ}2�{i�ۗ���ک֞L��
*�`��;!�ĉv9[f.��˷�Y8�Jp�������q�E�E6�g5]�܆o!gHp!�����h�}���E���8����=��ic�mO�Ԭyf��my����CQ9l9��5��f����>�L���Ow
	Ӎ� $?W}@@"}
,�QY/jQF_><A8����im�NfXh�6�������.1-����_����v\�l�٭ʀ���HMY��KZ�����ٱ*+}�!>'w��G*�n7�Õ]2���0�TAfؘ��F&�d�1n"[��ݻ2/S�?� ;_��hFZ�1?����%�C��p��M�<��?J��kj![A�mЙ�-e@a$a$e�o2��؛��6�l���`�����y�ɂc"]��𺶇���!�q빧Mjty�Q#� �#���J�ܥ׬&]���}q2Ȍ�m�ǒ�0�"2�������͢�<8mx�9�1}g.D���T�{�n~/�5ǋ�>��ݫ�<qc���0ׇs�Ra'�jư��./F-���=|�Uhsy��-@8���D[ؑ���t��d�9��[y:��|�T1Q��}l!s��X�}r�Asټ�'wH��alz׈�˵@�y���	3�c}Dx����W��&��/Y�>�"?�7r�$j�}�Wx��x�w/������Ͻ����0`�5�$V0�:�bQ�g��m|���n��9M�6��|��m4G�d�����g��:p�N�I���C�|�B5��k;N�M���tX��s�<Rl8\�C"�/֙h�hQ���J�,�L���ex����}V�7S�Ƴ�������yd�W��I%;
�
���5�,+qE��Ⴚ:zgsv�iy�ɀl��p>sz.�J�}9�Gt�0�Y�6�U1���S6���k�6�����f͔n�y5�$y���6P�)��"��P>ll0�'��4�#�7�����Z�"�n,�5��qǊ5�d�!����o-��>>���?�-��Ex@29Ĝ�o}�{�rœ�#�W�k�ws(�U�Ķ2x���j�1�e+��Q5+g������?�)C�!�7���Ãiဳy���C�mT��;��zPsIF2M0��D�p�oe5iuM�[�/{�4L�GO��$i�Ǹ5`��tp�|�-�ݩ[/�"� �`C{A`�z���N�(��dK�� �o;��}�c l F6�K,�;"��b��j&us4�aD�#�{Z��q�(��sy�Qa<։�	ʇ������X�㠎��vXU18bZS	,�gt�2Q�S`[?��b��Ka�v����23�g���u�[�(��
 s��p�T��g<�s� ��s�L���լ	O��?y9�x��e�N�j)	Y��P����}�X�N�c׹V��ȺnB�K�wi���-�Ngh�[ͮ��tɐp	iGo����Q��e2�X�X�"=�<2�L�i�sg^�a6�U.E��_ �8���rXJh��oN=�� ���rh�N��z�Ku4k/r��&�P+�L0��'q��՝���n؜m�$��ۑ�\�� Cz��T�ܰ��=�5;�-dC�Ʀ_�{���(�g�i�q�$,�='F���_tL?]�	�8x���:�C���>�0��E�v4��m���<��׷�a��2X�5cq�$;s��}��͗f�.�!.,�;�m��a儝.ఞn �'#�c�ڊ�Md�=�D����"��4lǹ�i�������:���pEBL��0L�0�E���>ƍ$�2�C��#�/ӥ:��a9)i3�F�uf��2 ����QL���V����n�%�"��%��W86����.�6��3�(]��V�r �5P�Q�a�����g�g�*��B�gi"��p���p�38Ʋ����/K��8�$�EO��l�2%h�V���w�-k�2��[ҿy��|��C���C>f4���1����N`�Xg���g0�oFU.jE����8`J�p%��l�ץ�C�Ʊ3"�k�5i�g-�G����j�����;���xn:lٛaE��`q�����v5=���mBD���4I�eΛ�~8us�Ӕ�FCi�5e�"��i���m/:���"���Z�{5\��3W	j�����*��d�f�K�qSa��Fō L�z�����cv��s�	�|���t�L�S]�V��ⴃ�`�m��u`�u�hvIç$P�b}c_Rt��j�e��Oi�i(���u�T��E%c�,���qM�˻�a�j���FwEO�wP�v-�����.j�&Ak�+4�_P�̈́H�~<���+�pΜ(�ð	�$F��T��O!�2 ⎐���t��D&��:�.����hTB,����"��c����;�}i�{��/G�����}�2�B"	����8�,r���2Ew����j���j���F�#�����,��4t�����$�'غU�Ɠ��E�"'SF�8T�k���:q���ff����/�1�,����� �+�"˙�{8
1���oVQӄq%ð���&���[\
7G�����
��}��H�k�ś� ��9�Pb�u�
�+�=dj�u:K��|;3����v��T-N���My9E�r4�4�Ǚ���M�z9��f\�;�᝵�j���"1��odah�7�y�ٳwܔ��z7UMlɿ���w����!W[�db�:t��ĺ7�mΧ9U!&�J"��(�i8{�	!��0��y�}S5+%հ�i����FkL+����DIu���݆n�y�Ì�4�������%8��",�]
}����5٭	��AF�OE�y�����27�c�/K#�����Y�����C_1X����s�˓חAV����_ͩ�d0�2]���y0sL�@S^�]��by�n8�O3&���e;�ϯ�z옏J8V��̄��e	kj*Bp��+��wN��W�v�C}N���0��� Ecz���d����:k��"��B�7]��7)�쟇�����$g2"���"�c2�qDaxh���R�{w7L�����X~xE�"ӱ�#��t�����k�lr�1'���M8l,t��i��d7�u@|`Xuǘ-��Ԝ�:ȇ6_O���1�a��@���8���/�c����h�7M�Q�4��2�h�f|e�����כrzXj`�-z1mE���/N!�oY�)Moj�t'8����J36�F��y�b{\T~+e0rB\�~�'��<D"�K��^0�+�?!R��6�}�ccE q��UoWz���j,�����������U��iocVƁ��Q���`�J�A�<6g+,D0������U5�d��.�����GD���^K�5;hms�q�]��c~΋EΊ�+'�P�ܞ��S�����r�V�	���c�W���zk=5�d�y ���F�Y�w8�XM��Ok��x�n��(��t�"u�m�!L�Uo��q�l.��"�g���5��b���T��o?N�S����2�Mk�r�Z���$�3�"u�,\�\V��r���;Y#3�½m~q��!�æ�g���[]���-��.GE�qɆ�(l��ә��(D� �����vA��$Է�ɣ�<�.{Yv�}��;��| ���sq4�r��ߜ527,0�^Ng�U��z����n4���;a�aYs솏yӷeK����5�
��!'������CT6z��n֭&�ʅY&����S�1'Y���9]]��N캇���Xv�L����7����k���*���tl!}N5p�t�ؖ���v��h-�^r�,|��>Jv\,w҄����O;�c�b�yV�>��(����*��ֻ-]�k![��Ro;v�B(�R�����$v�2�e�H�v1�3�_WI�������B�봒'OT��N�^$��x�����1����3�ZW:��@��î�f-S�����m��pW�;g[`�EÚ��"�uk1q�θ��D�L��O��ѽ6�$�i�.�m��}Q�w���!�˦��U�T�9�VֺA�ʾv�ECs2�w#�.	� (�]�kE�/I��̠��YGm*��20L5O����a�L*�2��u-�mӈd�c���X��YZ��T��ڒ�Ҭ�FD� L��O���ͰMg����P�$������)�/T�j� b{z��r������nb����$��c������K�eY�7���[�EI���v�ݝ܅m tU<n�˷$oE�?�	bC��̊Vݜ���z^㨢�)%��E��@�5�"7�]+�ȔrJ+��i���T�+�^"�%|�b�W�&�J�2�+Xq+�ٷk0�1�b�0u��f����>� {�+F�6���j�lm�-^*�n\�Z�^-��m��z�1�U�ƫ�Ʒ,V�V��\ޭ�wUWƵ�1b�^�_���Z�վ-oU|mπc���'�h�g�}���j��.�g.*�kJ���ʻ;�L�8Ú�~��!�Pٲ.�Z޸/���Cċ�I��]a8��`x���T6�7|�5�@�f�73��>��$�f@q͇ 0�a��19���u��n1;5s����p�㋎J:h1������*��{$6=[�(��B2�\ᓰ�Q\�����dE&�g�Agu�N�;���*��X��+>�ǋ���zy.#uY�:�4V=F�b⹈�A�5k�tIZ6��p���4Ī��\㶃4��d�x�� ��N1ź!s61("�hlu�x���Dpmp��K	 �4:d�Vč��7\�}a�̈́���Ф0��a�afE��gc�Ӈ�N>�خIuf���|��=~��yV�h��ϼ3�W�i/�)���|��8%G]����k�vN�Ԍ5�����.__si��;�L�k8F�p�p��\޵d���CJ�}z!��Tb~~(�C�ȣeh�3"�-�W�}ɜ�:��x8}5�i����5L�(F�XU����#I,Fd��^�� >2"����5�w͸ݶ
�A�"afi#�6��,��?�f���l1���K�櫇�i"M��G��䷦'b�W4ntNf���F�������CN�B�#��}���vEuW!�[�ư�Z�^�Σ���`;Y�h��3�����kP�a)�XV��m|�\��q>L�xw6p�ݎj�I\�kz���c���L���{D�x�O�m��<^C�s�*nb�*]1��Q̄v���A�/�M�����6�E)�\�q�4�W|s	�M(�,���NRgV@vnt�[wÆ�v_N`X#)U�h�O�e����湫��梊<c<����j|���SǟY�EC<\�
7\�pRL���L^�����I�3"ݽň�h!�
����'.� hS�)�@f�#��"�Z�h�$1�*�[�A�b#
>F+V���S��g�kq�Ǭ�Ӆo[@����Y-U�i�
:^����3����oa�f�p�õ�v� �(���Ľ�i�l&�{������|�[ ש����L<�t���A[��cL��f�8�$˰�aF���pW�^@����~���wS����ƴ�-��\0�aE@����z���ܲGzǹ�c0z6h�cɳ�qNXO!`�P�n8.����YS�)J��pnkK�M��4/�|��9�n){��jV�*�"���0��j��xt���[�U��n�G3�i�D#p��	��>E�����i`Cy�\�؞�q�:g[�ڗG���3Ն6�^-�d9{���ɨú�D�Y�������{x���~1�g�����P:_�Uq����V��|]Nbbi�Oc{yl����QT�>�m#�s�5N�g!u�ǵ��L�5�28@�"����?����P��N�'|*/v0�qiq{l$ְU3[�a�j5����C�.t�+ iӆ��O;m��&%.����J�e�7�G]��Y�A�S�Rt�"�+裭{]t�8�����Q�@�b�Sǘ���rS����z�n�k��O�{ۚI��ÀV�,���]�V����E�T.��h�ǝ�i���ھ�U.���K{��Բ;���!��<�ς�ʧ�j�<u�Y=o(۽Q�Of�p[O��w9���9_"�c��7;Wl��X�3�W��98GmE��HX�[�(�3��fHvî�{ĝ�ɵ�6�¦m��|���[f20p����r7���%�1{e��%��Q�]/F(��R6��w*�!�(�rL��M�<� ܅t�t��
��������+2��B:�9L"-O�G��?Z߯V~�Opױ�L�Ř�q�-��|�
W@��X�=���O���Y�����ϥ6E���d�u5f���\t:���2�C�c�KO�p����Wn��O*��*�#��*�<�W$'>��aꞞ��8 �«(�cF�g����S7��ɕ��b]��yJ��5�u�͝<���f�{!�������_sk�s��u�w\��1�ic720�L+�rtq`L�'A/��>��O�;�=:.��$v�ȇ.\�G��0"�����wץ�Q2D�..�ڙSy�$��\�4���[�;�jeVi�wb��m�OSq42;�\����k3���;*��(t8�a��X��}0���������<�/Ʉ�󿬅�堲�3����z]~5���q�Y����KQ��"K�q�ax��N�b��8�VYv������O64�f� 郅s6.ߌ�˗��A�P_�N�x���>ci���VD6C�����)�@G����oN��,�i�����2��(5;�`�:�u}c	�$�SukG=cq���}X��fF���p�h�{u!e�f�Ֆ3d�Ӧ�~�dm�+�N�l@i��%:_Ӭ�����Rz뾞��=�3��<l�sO���K!��`��X3PDtZG�[o�xQCo��O�e2�=l��ʌlOKu��x����0Y}�%Ɣ�C��F�{���`��-��(�\��i&�i#���a��M]sqX;��'�>�B�5!��""_�X��,��lƸޅgY���koXR��9	��,D� ׳��fƈ.�a��M�0�Ebx1��F��v���U���q�����+�܎#o64�S��N�
.5�ph���8��"/P�y��c�+�x���?&Ҡ(��<�;.Ș�Ǆ.1C;����[[/�ӻZ5�G�^Iţ�xq��[ys����WS��8u��->�vn�����-q�8��zp����`�6��c
�K����5�)�θ�	�7���S.!��=1��ٹ�4�$	%��k��(�4�v�)�̙2r(�Y��2l0��XB���s1���va���
~ܡy�g�������c�4p�q���w0�l;���UunF�1���i<D�
�q#Y���k����6#�c�,U�MG+��GD94C�Fȧj=-gy��@U��2{��a�F�+,ٍa���k:�.�y���v�mg�sn���:t�(��ݻo�A���!������ZhM����55�H����Y6�V'}r��rT��B�I�g�޿\W<�<C���T�v�Y)�����\��si˝]M
���X,�/ߐC)�'���jp�
���/J�)�U=+D���A�EH��#�	(�q7�90_t-𛫑�u
#b�`��Y���i�bAŔR�/~��8���-���D?xzߎS��w���;����1��j6~�-�5Qb!u��`�痲]�.��d*a��ǈ&;v	�� ���r�������"�`��6���A͇x�i�y(����:���g�A�f~�~�V6+?X!�=�Q���� ���8(U�Ko3���91��ODl3�q��Rމk6ې�:�LV�-��|ւ��fya�^C�^.,D2��<���=E�tΛ�	_��vغ|+X�#yr�fdB͍Q_�����{�l�a�[�^��0��OM
*�T�I"�%��q7>���/dNc�L��EK5���=P���Iu��u��n�y	�Y��?˶��?#�
���#lz��갷�����������kZ�3�@����aG9�{����0�E�40�}���'"2[���fy�+C�]���t�-���$C^2"�����ٰ���)�u�Q{�u�-��7:��&�/%��	xx��L�Wt8�̽W�uۀA!o!�8\����zؑщG(麷�l���7���4�.�⭨3,Q�����i��|���0r�܋2���O���]7��`��Z���,(�C��q�ɨ���?8x�e|(�	���Q3H6��G���
�DL(�J"&I�D��'�u�!� ��P��E��K�����C���bo����So+���K�&���rX�C�������5��<�s"�%�=�����w�f�i��0�P7�����s�b:������kՁ���qY��F�)R��XMq�K3��Ĩ_^[�Fº�:�ö���{�Ӥ�f�N[e �wD���3sCwt�\�v2i,�V�9���x>�p
�p�(���dq=g������b�n�p?����_�,]��c���Q�,T깚h�X󲱲�p�K*�\[�-ԛ�j�>�v����X_ķ*l�tz"t�Fr��p��!(K}���u��+Q� .�0�ۧ�T��=*��O�'k,f�9��1ޕ.��
������5܁* �)�B4�hK�&����ȡ��٬���+�ȑ���w�x2�Mǚ\�@e	m�u4���\�_U4�I]��r�n es�:�U<Ӯ�ʣ7���1V��p+�K�M@�S�h�=��R�����oV�!��D%��o7v+�'[�v��U�z~�(S]�����t��ύ2��h�&���إ8��+�6�rFn���$ӼL�������m�Xn��3*&ƍ��;n�۱��H�h��+�ZUY;�h��I�|k�u�xbL�3��.�8��+���w%ҝ�_Twx��"�@��+ﯥ�5�U}��ߪ�����b��.V�5�k�ޫ|V�m�k\��ݶ�X6�|j�����حͯ�U�z��V�z�\�x�W��6�z��Wů����V6�ܯ�x��o��ǭ���kz֯���ߥ�w�^}��y{�=��u�NB~�R����1a��g�
A4D&�H�I h�����mF��N�h��p������z���?|���ݲ�(�a��X�$��D@��N��L�!u�u�f<�cXW���oC0�bh�\��a~1F�;?tEw6caC���?�Z�� ͷ�Q�Yé16̲ym�W��Y�(�FSg5�#%�Z|.-��q �#-2{|�מ�`���>��b9�/���'��k$��	:Z6'n�������sY�|��v�Z�	����M�Ƀ'
�ޢ���\�y���9R���Q�#����j�=�ψ����B�r����I�$=Y����M��"�r<3���D�Q�L���8^UQ7�������wpZ�=eV��J~N�*�':�����*G&��/!��tξ����J�{�+Wtta�m$����4�@j�������}��Gʕ��t�L$��&>󓀄gY��ˎEƎ`��/� Y����i���/[N�Xs룭��۹FۡOਠaFψ�W[���h��oi~�ָ#�F��f�FF2&p�ŝ&С-p�ڒ�9�U��s�����<���*�/Jb���D�H�q��˟��Mh�v������O���	�N8�7kM�4a�r������l����#�^��~֣�މ���z�����w��h#�xق.���a����?´�an�]�!��-<ER�������?ޟ0�-�	3h����ƙU�ƛ]f�t�!}$�h-�
��if���X��a��Ӳ�L9�.wMJ*���6�G�i�6�kx��Vuڬ�Y�a>-q����Å�[|8���G�z0�7��6B�5������P�͑ɽsΌs�a�m�����5��?]�=A�5�<j��!�,�5��d�V� �cP�m���k�F����42���G�8�3�ͦE$`��]��~����p�
��\Xq-$<zI����_=cT�=�һB=�fϫX9s`��q)�r0��ҙ6⌎��$�u0�ZXU!
��O0�jA�9j2�=��m� ��pĻ��#:o�8�a�F�f1��0�!m��̈́
�㌜-.��l�68�ê.g�XJ�,#m���CX��B��I���V'-�MCz_�G?Yׂ��nv�Z2Y�F��9���UIS8wʚ�ޓ<!�L�n!x���7׹��ư��d*��4�aG�,"������FG8�k"sMV��S�Z8;��#`�sǸ0�a��e��3��i�%�i�s�)磤Q�v��!���]��Cו%0���H��-���2��ƛZl8|�aE#D�Iz#;;l��:�h�7X��6c#`��c ^�'�z����=���F�y��Lkqxk(�녬2(��E&�jO&<jb�$���9,-��*ۊ;,�f��#�vħ;Y���������U��'����I��c#cvn���uN����<D3QC�q�,!��Si
x��qx~��&ͫ#�U�4�4Uh��.
J7iM����y�u#�u��t_����4��n��|N�geZȺ���_��a����2�2s���Lh*��y��ժi2�5�'�S�`�0���	0�m#��6`٨��n
"h�U���I3m��+m���,�_0��L���V��ӎ<m5d;<p�Ӝ��kH ��=�1l���E:s[)��q|�,}.hF�E;��B��]u8M���F���R��h^&V��P^���4�s-�E�Y�<`�(�Ĺi���0���O3�9�u���Ԙ_�=�D����Egs����~�]��kΏsw7����(��~j!��YX��>�~�������)�V�;��f3�a�dM�y-ϣl[�Qt����v6M��
n�<��P�-��>��ӝ�;:�#����;�}�4��ۡ�]�,��3�x�ʳm�ݚ�9D�	�yɹ~�O�CB1D4�E��^���_#_��>��6�Ю�s��DM��&�M�І
��^��*\�FOV���2��7'DF�Q�i:;T�l����n����X˖��y��Fb��Cs�r�<~�d\_qmC�[�<C�;͇��W>Q�֭ǣ��HΈ�`ͫ�M�5U׬xĳ�6�N;�`2��0�F��-1�ͳP"oc.�|��b�U��ӵ)��'�����1��O��=Hx�,�BGH�hk�A�b=�~�o*ȯ�4��~k���"�t��`�-��v�Ty��e0�a<��\y��co1�!0�L��y<�<čR�$�lc���M
���.�V�%��_��lY���N��zR�9�1Ǔ�AԳT^h��$�%�:b^@r�3���&)v��y�x̅w�a�k惱��y:q�Φ,�G�[H��]t�Xn��JϏW������cX���g-�=݆/w��q���1�8��4�E�,>�+�������v��,������
ie�_��(��s���@�p�6��!Ⱥ�D45���]�舩��Y��/�(��a]���|(�#�-F-��m��Rb���K	�(�s��(�]spM��:���El�d�ڌ��M�&&�^�~;!8�`��q����bh�M�nP�����Ɂ � �L��KaqN�`�&�`����N�ᵱ�+*:O��ú��a�l7|�9��N��4��}�q*�T��Q�2���ych�C������3�Ws�S!ԝ��;���?"p��(��Y�TT}<ǭ�0���h�F�v�����^a���D#��M��L:_Z�K"s�*����F�ybO����a�Y�d��j̛,���gU���z^�o'܎>cCuѲ1k����v�UOa�?��a����y:GV>��p��M��tZ4t2�0�7L��Z�00�g�
뽐T��݌���x��ad�����aDͽ �*���v��1	���G�XB$!G�8���4�V:3g#h��!���yt�\%��S��p����b�u��;���b0`��Nb��������R�1h�K���n���f�\���}�6��÷�U�F�zg;E1ŔA����&�v����×��<����[�Yn�̂1G)lo!ޚ�d�,,s2��/Xltǭ4��Eᬣ�H�N��b��s@Gm���w6�#M����`#����EM���#���F��z�ECa�9�Ur�Mc	�#g�l�"�pK�&e{ӿD�U,��4b��%��f�F4 >,���ۺ�nQ�D�Ѿa�̗m�t0�A0jl.C�Q�ϡv�c6�x����^��3�X:z��g*Ds,m� ����#0��3,̓��m9�;�Mi�p��vY����DO�a�af�TEbg��x%�ߧ~/�,�t�6�#�4�]d�"��3�#G��	�����I�*���\m����{���wR�-�IC�_\�*5��J�E�=Ƌ����|��2�s�T�w�4�{�g��+Z�N0��C80���i!���!)��9*<�N�U2����d��֛o<5���K��E����j�ӆ�;��C�8���F]P[���fib�����j�i���a�'�]���u6Y��:C��8�[H�h<o�)h;�Y~.�t�~�8�q�N�kQ\�4x�k�`���tz�;VB\���u�v�'[-������q	��`N�.`��˪��5[u�IDrj:5�6k�d�Ǜ8���C\8�(�nj�����c�1�qn�B&@��8H8�w���R������h�<�C�4��rna���J�quE��'����UՇeC�kH�����\+{ra/i�/�,Z�W6�.;ΡCk��z1����UJKq�Ֆ�{�4!��z����J=�K�4-�9��f��a�*\P�:��	�v[����������-QЎ��`�29&ɷٷ���}���=^.P8�����BniX����L7Zʾ�ㅳ�1{���#R	do(�A;��'s����v>�C�M�.�S|����Ͷ����ecb=�ǀ���魴�=�Re�k;��P�zg�C��:k]G��C���ٙw��LWk�D+����B��\��*5�C�}��-: h's7��Gz��^tj�KV%݄b]��_l�8�Z]���T��ه��c�r:�z�=W�ݶ����f&�|�V$�9�"�k�I������\4�4@EV>p]_M)��4"��<r��NL�N��֦���gq�6�\�b��iΧ�Up[�'&���O&�2�/���Y�E�ü�V����	��:�#D5��ܜĖz�6�P0���oZy���w3�X�m'Uf��\�rp\ؚ��EW$�5\/�X��:!®e����H�d���a�tA��x��ֱYh᮶��.3 ��8&,{Ң�2>�ٵ5�Æ]�����v�!6�]:�k<�={%���	�\l�IR��ݱ͑$T���ɥ��+�[��V��v�v�:�JS���A�;+yu9ܳ.Ք�-BU��^0�MH�&�@��l?�}��~�����-%o��V��k��]�F�ݶ�F�+w�sE�X�.���U�nm[�z��h��oZض�V��5�mm�mꯂ�-��zۛj-��[o���ޯ\���Uʍg~��]�xy��mJ���=\����1о�f�V��sI�Yo���f����\�0�j��[no��y���w��3m7Ty*P�8�
aF����Y_�H~�V�mX���d{���q
~ve!tك��d�Y�V���	8�+z���}���g�l�#EF�?>[��i*���m;�擑���i㋞4rYL�tTB�Q���a�m-��v�u�*�78�52�Y3ݼnPg0��8^���j�_�Ñ�WIy�E՜�,�����>&���%�ӌ��yaQlW��>V�����,"��m�k�C��"ڎ�k3���_X�T��u7Y�1S��+rE�6Ǎ�BF�2kv?U��UPtaL~�`ʲ�}�c^K�6H'=y蘽H�����
mՎ̒-�F��Y�Q���?�bˍÚ��Y���0��xh�oV,a�w���1�L�ئε,P13��Ť��`ߧ��C!+d'|���Jٻ��f7�*}}y��a�C:k�U{ۆ�c���c�X�V���a��s��v�u�כ�A��Y��ޜ��o���5�����'���]Hi~�%=�f\!Sޕ��Ot]W��͇�|�hl[��jnx�TxF��-��n�j���yRe&��y|���qR�`�����r Jl-i�L������u{)��kz�Xs����
�_U�3.��T4�Zw��N��J���`�@,��_r���]�{��jt����]w8���l'��ۅ+�u��wk?[�ѳ�/�=�x�{�V��͂�x�	�cu�|v>k��̋g�C�A{xN��r��t���$����e�@�����Wg�;��/|gD0Nּ:w�����=�|�)+%��ݹ����j�h"�ܽ(��̀d���RL��K^Wf�r��w���[�����'�Y����Y�{<��tP&�Ñg��/*Q�x�����:�d�*���8�n:1i��f�]3oiu�+�VaE�{�юz���R��^��mO\��X����nu��P���:q��s�䆥.�)=f�G{�At?nS��jb�꣯mW�7���;@X�_�;oY���e
(gk�:+ΖzL^�o&ά���93�AքA*+�H��K�#$�wko�T2��k�������P�2�>��·�c<�M^�$�*� 4��[;:e�G6��u�`�Wl�Ћu�O%���ȟ����M�=���ʼE���m�N�����KS�|�j�wH�ubV�˚xS哯7:mh�&��a>z���gG^�����c�t@G��+����=+2��m�C尞����үC���upg��2]f/�}�Jr���q��/l��
dĻfV�ٖ�Z�f����ٺ���t�;�c7,hL=U��sSľ��MI�*�x��1{냰^����yZ"�}��U	k��*S���{o�n��t�zX��k/�Q�=��\�x�q���#{���th�����[�p�����fm9H���{Y�|lC�X�pt������5}��5b�$�8c���<���^%ɞ���pe��}y���4����\Ӥ�w�&�]���R��y�qyn�·y@��*�qH�#�g=�N*Al��+o�\�=at������	2)��ԞOf{��֕l��i��s�5�RE�P�k�Յe�N�x�4f�{�����}7��>`��	�g�5��ߦ#]o�TA�����\ڜ��Ǻ}� {3��{ �>gא6����,�ݘ�')�řz�<	���r����\�5 ���Jd;s���J�3��Z����"0� �(����5�PR�A�q�xwU�ESkN�����m��	 \-����� �)��K�%��Gr�׾;�8t`���@�!:��A��v��i���ͩ�!E��>͛�p�����_�;l�T5��kw-V���wO=�|�J����u&���l}��3c*H|��vΜ�3�q�s�|��=��evCM3���Gئ�������_��_u���D���z|�u9��F�	����ΜN��#������#��{D/��k�n����{t��L�o{���U�VqCUA����8�_-�eW:���Y��*���%s�K�ɸ�"����^�Oz�g��W���#�@/�����a�)�Xԣ�r�ԮJ}_K������͝�o�dӹ(��'R�~���U����{Uv�(����`'|�B��˳�Ͽ<x�MϣN\/-W�{g'�g��@ְmh�VGkW�&�gR������Fl/��J`��➓�vzh:���è���tyU77�y=GӪ[�4x��bcf
��~u�G�*�1�c �iu�K�Ŝj�˕���{�
S~�����=݊G�ku��mi����Tل�B���vg6�z��g�Hg/i���׷�"��nQ�v%���i��ؠ�������=ֳ���q����>�A|�g,a�D��G��*����`w���1E
���#�ZX���Y/U��XJ�"/}<\Y�3ء�"ǅdW��N��ˍi�]�Wbr_���<)ܘ6����Z�S��n�N�n����F���ݲܦ�0��]|�ڛv��ּ��������B�b�z+/�_t��P��7,po��uY���ʂ���J�P[�S�Q�N��o��vNǸR��ގ5�̫��;�[�We����;�A�4D�i�޺��
�l��C���ε*֒uTʙ�-]���8&Od�tC���f�;p�-|����dr���kHx����"�����~�Y)��j<��ouÌ�c�D�/��Z�ve�{�ޕ�w�V�袤r����e��������ޫ�x;��i���rz�Y�z��4�"Bq6�r��� �ztG����}�ߏ����߿����ѿ�j�?�\���g9� ||I���mo�{��f>���vn���n���o�U[_�y_ۿ�~�o���}W���&�+]-�T����˯n��V�Z���>�V�^1Z�_.�Z�Z��&���}����Ƶ��SU��i����ڿ�7������j�-�v������omU���X�_g����{��������������M�o�~�!$B�H�"#2BD)L��@������DH�)��3 �I&i �	)�D�d�SB���H` �0FP����H�A$�H��K2a��$	&H$!L̒�20! Lș��� L�@  7�|����ټ�~���ߚ��b�^Cu���w�$��\D���HD�+������30I0fdM �i�S%���f�h�*E,Y,�Ke0�K#MK,ٴ�%H�L��f��)dؙ�(�S%$SLL���B��I�d��J1)�&e&a��L�JY��f2I�(Ȓ�$A&b����R��K4�1�F ����๶@
?��w���)p$	r�~aaA_�:D"K3�1�b�b�n����=C�PE��<���3�S�����8 
7�`|��&��a"j�"��^��k������j�v�nZ������|�K�J��;#vm9�xs6��(r��f2gȀ?�X��`V5@S	�fș�X^�Zֽ�Z���W��^Ҷֶ�ֵ���U~>Uחo���e6oePP},\&�ɯ�м� @Q�,��� ����(<�D8�(:�Po�n-r��@�KhG��Y�%�G�����4h��q)���	>G���]���F\ (׭$��44Z����9i�(����m%4Ԅ��r�s�ȷGRp"*�-D��;����$y��x���a�TG4�@����~���R�ڷ�"z�uX{Hw�u��(Չ�`
>i�@�H�����H���f4��	9PO[���W[o��������mV��_-����08ّ�BC�.��QtAA�4&�$6�6���Q��Q<:o�9���,�m���6Z�������kɮ��o�/~����W�VÀ*ëq�v�PڧB��Q�8��a�^`�0�����&��������3����$��t�����N/�1	ڞ
�ɰI��2�������A�һ#@#�e&@<���/H��EOϸVQUh��4m���cUEmQ�UF6�cj�V6ն5�mQ�Z*ص�F��-�U�kcZص�صj�klmlkV6��b��ŵF�mElkUF��V���b�TV�jض��Z��UZ�m�m��{��p_ɍLϳ�AA�pv���f8;D&k��Pت���a&��� ���2y끯���1��n`�C��m��x{K�&��(:B
FH(:��; ���qކ�,�
�7*(17\�P�^A�pH�7^�jN��9H�}���PBA�P��Cb"����L���y�����<�:m�G��8�Ā�Qɰo� ,֬Y����n�dל�R�k!��$���1ѹ�EܑN$��� 