BZh91AY&SYlÅ�7_�`p���#ߠ����   bA�t�            ����Պ�lj�mmfZնզfD�-��"�A��V6�Y�����,�	e���2�Y��&�AY�R��5�-�u��j�۶���ٓt��\��YJa�ZLٖ�V̛ml��E��Yd�3��-���5m�fdj�ڱ�jj�EVʲJm��m�Uk�@<  � ���u�����jՓ�k�j�cS6���u�T�6�.a�l�j\q��QJ�sEckl����]��˃��"���ڲ�le���*U�m0��aR�����׻�]�چ���q֎k[�ڵ�҂ݗ����]�Zr뀪um���i�v�������-�뮺7\���h5v�����^:M�6��-�xEw7�G[� *:��P�U^׏�E%Q�s���P�9rݡ
C�x潲�R�E�t�5�ou[���S���ǀ:R�3����T��ؔЌ�T֕f"�a<1��QU�p��T�kW���� U�����W���B�w7�뱪�[���3�AU#ӝ�� ��wD�ƭm�F{����V�yy�)骠'���%(tm��w�<�p��jɩ�z�T��w\��)H�m������W��w��P�>�}Ӏj��b�}�ꔪz2���^��*��{�!U�TY5+Cm��3�uUJheZ��*�J�eRuKVh[�jimKMj�xx��R�J>�hj�UV>��P��]XJi����4:I]�\�QUJC4DT띪�P�T={���P�����	T�6W[mf�mM}���m���mi��JP�R��}O� RXJ�m���JU{�î����{���R��:�gJ���K�ܫ�CRu�^�� �'���0�U��X��j^����ejZn|Ҕ)T�u���z�8 ��n[���3Gm�۵y� :.�n 4	�n��m�M�@����� �n;+Z��kj�ںl��M�O�*�UJo>  l�p�@Wo������ ��  7F�4����
=� �-&hh�@ ]͵m`2(���A�(x�}�UUD���� wox /)���\  s��EzZ��Pn�s��o;E �=� w :��m��-U[el��ڵ��:�ꪅ/��� &������ t�� ���P�� h���Q��\�wI�:��  �   >   �� L%)J���@F2i�S�bRR� �L&&ba4h5=�RUT�U0     	�h5S� IQT�  ��  $�JDd��@ 4     D�eH�4�2d��)�@z��1���z������V�ן�����?����c[�^�O{۽B���̝*M�9ʻO��=��{���>��B�z�I	#�� $�����I$I?���/�ϡ?�~����������?���Z�mm��ˀ|�U[m���O��D$I��`��,��%�?����XO�,'�O�(��)'��D�d�D�R8TN�$�a8Y#��8RNH�R8Y$�Hp��(�*'"p�'�!8TN$�D�Q8Y#���N$R�,'
'	p��*I�Ȝ,'"p�G
���p��bG
&�	¢p�p�'
H�dzR)EH�Q8XN��N����D�d��#���I8Y�
'
�§�C�	¤p�'"p�'
���p��,'
)Rp�8T,'	¢p��*'
�K'
�p��,���,'
�p��bG
�T�N�D�a8Q8X��Ȝ,���p�G
I��p�Ңp�N$�,I�Ĝ,���p��Rp��,'
�p�����a8Y#�����d*I¢l�G	��p��,'
��c��8XNM��$�dN��M�#��p�'$p��D�d��D�d���d�N��<)'
�8T�p�I¦ʇ$p��,'
��RN*'"p�*'�D�dN!��8Y$�R8XN$�a8Y#��*#�����2
�EG$p�'p��"zY���dN�P�a8TN���p�'���d�$�d�p�I��N	p�����8P���Ȝ,'	��p�'"|TN�$�P�b8P�,I��p�G
'���RN4T�	�Ğ�$�Q(aDp�I¢p��,'
'
'�D�I8P�Å�8Y��N,��RI�d'
�p�'	¤�I�Ȝ*I�I�D�D�dNI���$�d��Dp����D�a8X6Xp�8XG
I�a8T������$��`4X�p�"p�!�dCE��bIK"p�8Q*I��p��),��ÅH��p�G$p��),G"p�'
$�I)bI¤�,�¢p�'
��Ȝ,I���I8Q8TN<),'���,�p�p�'
��Ȝ/���RN!��p�p��,I��&�)
�K �Pp�H��*'!��*H�bM�p�Gp�,��R8Y��p��a(p�,�¢p�I�I8Y$p�&$�(G&�)¸W
�^�p�8a���,�<,p��NN�'�X�§
��a8_K8W
|V�8Y��8V���p���*p�/8W
p�p��,�\,�g8Y�����8Y¸V��\+��,�g�p�p���)§8Y�N���+��+�p���+��,��¸Y¸X�g�p��Ne�N¸W������+��+���p�p��p�¸T�M��N��e�g8Y��8W8W
�\,p�p�
������¸T�\+���)��)������p���+��p���6c��+�8S8Y8]���¸W
��8S�h��/�'
���++��,�t^p�p��zY¸Y´^p���+���+��8W8W8W��,�XW8Y¸Y¸Y�g8Y��+�p��8Y>(�G����p��z^p��\+�p�8Y�xXp��N�f��p�p���G'*xW
�N)a��c������7���*<%`L3�TC~쵿՗��fPN5��d/Cӗ,0���j�h��շ��4غ�l�v2��r�V�ċB�����%�N��H�¥ᗃq�9Q�8Te٪yx�;���Qƅ�G��1���"�"m�ǚ�^���p]k�!�
,�B���U����j�1�Q�a*�*�W�xbU��'KK{��hۣ���Q�?�̙`��aK6�]ݪ[2�5�<-�(V�he.�ӎ�7�ʏL��%�[Z˼ܔ�������e�T]*��Х^�*Q+�V����]e��X�����OqJR�M��j�lL�X{oJT���c���$ݣ���7(�Kw�^7כ��T�UF ����$�T��;��57*����-�l�`�X۹��-\���6[��2�e#z`̫��N����NѣOX���7��505�b�F���Nv�YeR�Bݺ³pJ��;�@F\����*��K�m=���*����kT��Wut�n\z��[mִnȔ��S4�[�1r5d��˥��j��8^#�6���X�#5h�U�=Tql�髕��Ȳ�l���M!�,�-ܱj�$б�ɮ���(Rȍ�KU�h�h9�X��2���6��W�2��V�x�t�"Z�oI	�O(Т�5k1�Um4�q]kA(jeMrR��]Su���N��Wf���#*�[ID%�.�P)����k6��3#n\	�JAt��30�V��G1�弭�"�a�ȯ6����g\���e�$S'yD;7��h:,�v�ԭ/c�8/0а�潇5װ̷[�d�cZ-�P�S2�e:5���wi�xfV�m�ӴDwOu@�	������$���d��������,�A�Ku���T�51���ܧR�LʳV�쑑$!�$���٘E�5�X�5wU�u�,u�Ʉ\5tq�G5���7)rJjQ�Ecb^h,t޿!��7U��찁Q��n�a�&&2
3��q�O(��J��o���<}]��$	"�t�����:�h�h�KЋjP,μ��V�e�&�q�2л���)췸��N��2�*Gh�j�R�p��J��jd�/R�hݪ	h8��v��j\K���r��gL����ڢw��/Pe���h�(V��4](�p�l�r�M"�I�j��)�&0�#Q̸�#�U�Z.�|�q�5{2��-Ё0',�6�(��*�V�ɔo?6�&��^�c%���bdy0�d�O#��lfBn(�ݧ/6��kw*2��i^Y�ȉY��/hoK�.;�h�L���ʹ�j�ս���v��@�m�rd����jR^�����B�w���Zcx��3��Tt�wK�!)��$��1���F�Q�Wj�[�b�,��f�-�N������x5�Jעeƥ�ܱF�kّ��������[8�H�č��;�qJ1�:�;H�Vإ��O.J�1k�V�X-;Q�E╸��nUJ�kE�A�)<�0��kNP����Z3V:���W����VV�\QК~Te�|�u�^b�Y,a�:�n�֩��D�p��C���]!��z�y�ł�6D�AmX�õN*�[M��n�E�1\�]�M̫T޹G�r�G�rk�MD`U��DGT2(��f�v)4��X�n�#&�,�H���.k�x�����)��# �t򔸮d�D2���"C�0νYQ��0!T7&㦪-�NU��x�ě�4Z�4��R�4.��-��D�4�R���ۼohi���Ә6��V��x�mc[E7��K7"v�B=�<�{���X�����6�(Jo�5f!a��&ق������˄u����:�)�-�IK�2�(��]�G�b�v�K������WU��I�KT�m�(��fe4#��S/�	UK�C:�+R�5�Zi]����$��!���6Ee�^3eВzMn�K�¼�n¤m�/Qy��J�ձ��؊�F)�2^��ѩ')F�R���v!���M�0�k ���)d�}%�9G��7IM�r+�̠�b�K��̖�N�b�U�	��h��e�����H�n�8�ڼ�J���f�+��)�f3�J���QV'�m(T��)H���A��)�jْ�o7-i���M:�kYK)����D��=���T�bYĥJ/ib��r�_�^X�T���V��V[IZ�i\�8z1�:��bv*�+��me�苭{���I�G[�V�є�Ǒm�)�wP˺����^*3v�lҤ�]P�n�*�/f��ME�R�OEi*T6�Pf��C��պH�7���6�%;�-�Oi#z�q�e^U�D��X��i$�y*[n�a�%E����X��y�L�CV���ʌn orK!��0�ѹC�r,^ܣ���AD\V.�K3�i�y���cT�WA)*H�o0ِݠȭ�;�S�{��V�\wU m�7���t�I����	�-k�yV"�a�e�-���s[�I�5����(�'�Q��-�y��[p0]ۧ�t�W��0JY��Jmam��SPĬ�uR�-��a�-ݨ���q$�2�%3e�e�����Ny�͚V��7m$b��6�n��ɏJ���*��Q����2�E�V����ڀ�J���L�%�&M��&Ҏ��ۗY�����ܘΨ ��O��M����B��r�F����c2V\�
�b����$�Rڼ��O7&��ƶ�#����JMky�n�nĪ-V�e����M_�ZǐE��qb��wn�1Y�.M���[��H�e� �M�,n�\��aP�.�'�˳1�X�ܫL)
�ӑ�	�D�Ve�(�kM��V,���4P�zJN!:\8*��k�%�ԛ����LZ�� �~9C�f�!+��ҳ��[�S]T�H#�WW�\�w焱CU�gR�jj[��哳̸���0R̴	R���လ��ʴ�Ȗ��e��w�$�.�aux����,ܔ8�9O/t�ٸ��dGЫ��GiީQc�I�����č���&�[�ӊ�*Z��6�q1�Rg��T�y�ؽ���ȃ�-avLx0^��p'�R�wYT�U�q�)y
�Y����Y�=�D�J��%���*-!�'A�~*����,J����h�с=N6n�n`�D֋q5�K�v�]Ik�f6�hoM���f�a�������&M��Ԭ��5���o4Z��j��ux�k���Uvkw[�4��:�J�X��(#��L�J^Q��N�9�;�	G5+�UY�j�#H�̘�f
f�DݗX��p+��&�x�k'I̓6Ee(A{��T��6ܹ�a`�����
�%T:��/J�M�Ϳ�a�G]5E�k6�V��]n�;5D]\z�B�|��w�'i�h��؆$��k;N�k(�E�v��6�u�ml���(�#W-��O\�)I��0-8%"m�v7�4]93kdXʂ�h[1�y�ݹa�.����Ѵ�0ݓ��S�.D�QQ�vE%�2��$(���v�Ei&XAKY���Q[�e�p�Ğ��M@eZ6�j=��9v�f+UQUbX�3�[�F0���T�&�sR�5YU���<�tI�v�J���-��V�Խ/iz�%�$���{Vl+
�̚�Q&���km)a���`�:2:���[N�J6�ӣme7i�y�{�1�6�L$-ˆ+{I#���r���ѥw�/#�ݡ�Ҩ�h54kd5x1k%�m��uf]a#$NY
���MB�����z�;ں6)��zą�Y��BcW%�q�W�i�mɊ�xF����*h��^8��m����Uo�xV4s^��ۇ�ȝ�u6M�e�� [d$6,vȵ�����p���b2�Wr�:v��wȩ�X�'F����T�F��j
�)�xXEd��o����ʽSq=t�b�q�b��p\���e�X���/�oK�n��m���,Z��M{��u���ʹ�=�jn�	uM�k0� ���3`�Q]e���.e�Z��K
���O\6n��{n�m�(,,�qכ+Xt�V��ח������ݧ�2���4N�)dE���Sss#i�f��R�kF�b8��e��.����.�-�;1J�r�Q��{V��L��^ �3�.�V]�.�7.&�i���6��Ή36�͵����h:6bT���֓�4ji��{��5�
	#�se*�G�A(Tb���͉�gr�q�06q=6�k%軤��Pԫf�4�K,���ńK{q��GT�r'�7+�i�KU��G��V;J�w^�I�׺uh�Ԩ5�m��hy�:��ݙf�el��[H-wA[��5�É0H-Q�Wtv�F�lb��uy����n4�EP��b�[n3Ipd�Xj�_�j�z��)���i��f�3fE�I�m�l�WR��eVk9,#�r�S�Յ֬h��vwwlJW���jߎ<@�W�
�@���/
vbG+){Q�71m�y17VTӲ3Qm��0��P����k�n~kjn�ۋ
�n�IՌ���0�g16lhf��]eI
��r�UT�91T������f֌bV�ӸM������2���%l�d;~Wp�7"�c&��'��"[��v�71`:��g��˼�r3�;U
5���|Bz�7b�^C��#(m�8qG��;�׮c1U�*Q�[%�ǂ��Vp����t�Ká& ���q�lb�&*�*ӡ�W�
�3Q��J�jM"�td*�hTl�I$�5J��^U�����׹�P����j��0�4�<n\gS�E[PG�\��UR�E���K7ٸ �BȨW&�]�ML2a��]�n�󩖍���t����n�"�;�K&�f�5��;:��ػt�X��[�����HwW,�a�1+V��,�����_�2�{p��(ĉ�m<8��m'�������R�)�iQ�x�T\[{�U	�lP�Fɢ�ie����K4�j����P�7U�VMI�$�L9�%���Z�XnȌ�5O˂�B�^L��M藩��㩋M�2��4��/cV%FB�
9W��w��	ZX)���⧘*ˈ�%q�G+�H$*�I���e��+%X"�ZoB��]YNR�+��F�RF�dcnhQ���u�>[D�q�/iᖑ9��c/5(	n*��XEؐ������n��v���uB��3s!u%Ԭ�r�+M]��smke.4����*\��u���t�ֶ^6�ӹM�r˗M��
�i����A��[��3��22E$�tÔ�`�J��2f�36Z�B�P��Ū��[���:��0�*�%	t��k��B�D�x�	r��H*Y��Um�j~gM(�s��-�0������o�WN���z��ɢg5�!�s���xfUZ�Ѫ3"��2^��!�8)b#�nY^M(8�%��@XFĨ;qZ4!� ʻ.��+3
eg�ˍ���eW��7C-�qe�-Z�.-xв��f5���Um��5h,8�N�[��XѴͥ�82lܺ5[p�R �uU��1�lZ�"���j��ô�m���P�
6�BV�Yc��3�O՚m�wZ���$-�yy�"��:��tF���5Wj��*hV��Eʕ$AU���γOj9u)n��i�%�ij��-�fk�Z�����Fff͉n��<�U(������2�?�R]9$��2f!�V(u�vD�DB��L+"�|����FQXb�M0��pm1XQ�6ȫ"R��cn��Y	���J�����bHPp#΄ �{H��\���օ ��D?`�����`�ª¯����~D^�)1U䘫�@բ�05Ո�yB&# ��Qৣ��~�B�P/C�	1�O�&"�I�(��Db�j�- ��������O���ſ�\)�V9X����҅c��""�
_� �x&Ah]`r��<���G&@։L`)�F�$*!�A_� �.�t)\DV'�H�8�R	p.~�*�E��R�Q�U�ߵа��>�#��
L[`�4z�|+ �e�`UH)�\D��N�b!�&Ax�Z�As�t)�N�3�\X����J�H�]��3�����煂)�"CR�)hS�
hT��X�\�[���Z��ÿ�0]z(h����4I4�G�!8U`Ղ��>��2��DoW����ë*�Ia���`���c/��<�|��¡��`��{�4U���bn�W^����7��-�VTao����-�)�E���׭�u��0g�=�,�8��07l<�e��h�`��<�hi�Q 6������Д ���ǬbA:He�J�جB����:{��}Z$���(4��A`��]AkD��1�D�/~�)hR�Qp?����b��=��>����!�A���3{���l��~����Ub��xcB���V&pg����5������k�����^�A�h xuЎ��ځ&�uXJĿ;B��P��/�|K�c/=~�=%��!�&p�Ķ�[�cEU�\/;^Vрj����8��ڄ�>���=�
�,�Y�^ș���v�N��"-��Du��<���n
�;H����P)�!":�>�aJ �#�#�F�{}����D���x����]�x2`۞8"�yA���
z'P͡]�]P��R �l'��+�ہ���%���eH��]p;�SK�´.hZ�=��fp�B�"j�7X۱J
,&���%�l�x8s�b,�O�.�`k9LP@剳� �f�pl"n�
�(c�T`^�tAlt���@G��aV����t2�B�0�?k8f������ZA�`9a�E���3�NC���l�3�����aa�9�?.�VTP������yow�������7�B��ߡo^ �����8�F��k�>w�7�<�	ƫ9L�u
�@�N���E�8ȱ/*f�$���5g!Y�nQ�Ի�Iz�u�r!�
��Eb�}��y	Z-@��Ԃ"�&����c:^�(n�yv�U�����7i�S��3����33�ٝSL)Ja�1��e�ʸڥk#f`�G5������5�Z�u����P�l2�
��fp�����Ė��8XWUʟ�0�F�&�GfT��B��	��ۖ�H��ˏ�����@�Q޲�����*���qg'n��oBu�D�����y������Λ�]=C6��� ��P��q��xWz���R�ګ�S���"�M9��7Sڙx�vY�E��we��g�}��h���o/�y��WEi��}�ޣVd��*Ш�4���<�_C��e�� ���vp��t廓2`ڗ�'LFYG%�q�=^ʪA�h�jsry�7��ٙ'!uH_p)��ت:��0r�)srɮ��O����r�r�{�we]�AF������ʋ[h>!q7M��JҪ������˸�,e<�gUL�4f<Gv�뻼�xuq�z�Av;��l�|�R�V������B��{���.�Jr|RQt�v��uy��O��o1��]�qvoYA޲��Zj�(3C��y�;�\M���%Z�;CiT���=��U��
c�!�`���yfJ�=����AoҠ��v��a�5gPvw+��#�ZB��t�Tp!\�WFX����ys��I�̣����n;��mo;ۘ�&��9��/*�zs���m���,Pf3�����n��ϲ�5�Vf��]!(��#2���U�hr�m�U�w�l�c��Z��NVM���/��_`�����ݵ��k�rsMW2fh�Ń�9�Q�T�Ya�]�ط��5�5.	�Ǖ�^�o7m��p�N����gV����brD�!m��(o���9p��P�Q���-g\��6ڸ&�0L��b��F����b�AN��-F���c2U\��&[�J˘��jV�r�#]�<'�+�npi��c�e'{L՘���6��J�
���yU4+3�"�I��ꯟ�UV�T��P~=�i`��8�B������6�d�} µ+e3���X�ԣ���|�7H:��H�h�Ὂ��})a�r";�y2��Դ�:�����nn�Ջ*r�W	u����뗆$WI��E��Q�Ae=�6�*��A��a�G4i��|uQ4$�r9�ޮν�s��/4N4;Ia8��w���]�Na��)蚇s����Qy_;ۄߚy�Da4p9�]X����<�l��Z�`WA�i���zK�� �2��G���U������+�R�Ÿ���0|����f��7���]�]���(7-5� �+Q�$�����}�Ij�F͕dU�rW�X'����I�āī��۔iT|s��Am�o��P$}j�����踟b�}�_�X�8�q��T�o��g���Ke�v�VFԉ��g���*V�~��<���{Q�F����V#n+p�{� ���ۚԨG�3V�\�����Ƃ�u�-�hNh!��ClX���t���������ٙT���̹�����iPީm�%��l�2�\6w^lW�o��J$_q����ȝ����Mvmx/O9R�;�D���"�pS*7�"*B�vX��=�P����G�u���G�o��'P�}�f��nW>.�Y�zV�UM�&J/��,x�է[�af�k�K(:���E� �ov��ܗb�dK�D�v��E�赹��ڭ�\���y�m��IbY[4gj۲�<E�r$Q}V���)RV��cD����H�ǅY��ʲb��U�E�R�U^�bpOy �lfL]��t�/.���uqud���N�grJ/y��|i��R*�B3����,��y�y��r�:	r{x�qV_qT�av�V.Kp:�d��T5v�ᴕZr����2����d�َ�)5)ev����ݍul��ɛ���wϝ nݡ�m<�����W�7asA-ҹ���Ew+��2�c$�t�-��Ռ�s34[}7���ګ|/�wb]tS#��<���E��H��IAb�몫y1��u׾��Not&k��YR�Z��szVU�ޠ�0�}�=�/��m�R�Ȋ�{)�w<�nu����:=�-��QϹ�o�Ց[�/KH���Z"Q�(j�v�q1De����帲����h�q�gX�\aY�*LF���s�[�%�������S9SQ�N�Zw�ÕҴH��s�7��h!wQK�B�#$ï*����<�7{������.�F�/��t�Â��CB�zD��4�����/QMJ��#��έ2g�Vb:�UIؕ�c���ݹ���]vC���ά�]�g;|���\�D��%�zV���[s(&y�텝�-]f6�32s�뫧>�:��f�]5�C�Y\�m��Ջr�/kK���3M��|�Ua-&\�Xf])A^r]�O�w���6�b�r�nW;�k�yM,�kVx�UM"��x���F1���z�t�Xu3��~���cZ�F
��h���"�S�{��k;��V���PY��'(/��i���Rm�v��3h�З(:�X�5ם48���,�.�:�9w��3�]�J:�y�u��%��J�Ȃ�\��:�=v��׏��u�̇pΌ���e�y�s5�G)$�W�'u_\�X廒os���m��w�.Xj��˘����n�-}�e[�U�T���]�T���9��2����������'+��ڛn���a�K�Ŏī���������Z��B��m'l�w\��˨����cȍ��mq���F���z�u��L��6�i숻��
�n�R���9��m������:���V�=����q2f�k���X]��q�WUS�1��`�����k�r\;앑s}8u�\�m�ψ���c*�9E>W��v����f���m���ڔZv(����
�4�z�T�*�y�����g;[���Pn#������_�(�;S��R��N�1u9�S���'��W�ܪ{O�o[M�٫�8t�t���|�_~]����GQXfI���:�VrT/�u3C�\���5L��T-���� GfWk��œ8R˄h}Q�V�����@��MY�z7%b����<���)�U�.�mVM���:9�w�Zh2�޷�#��x]�����Z�`��.IyWn����M+��V_�L]l훝���ԙ}un<z��G/�U__I��3-�]���W9*�L���Y1��4e=Q��e�M5{Y���%)r�����5�zVnǸW.-Y�}Bt�p<��C�ڮ�M!��˲��(IZyBw��/!v���q54UvgkU�Ŗ�黙`����ʡLt�b�ׄ�Ф��'d�<(e������r�ĺQy��\5r���l��^^�8G����\}{���WL��ε��<�T�2T��9�*n#�*Ձ̕5K=�	�˳�I뻨�P7w�<�G�;�f�(��[��Q�7%b�e�a�>*� ��*�c]��"�D��yT\��9�ˆ_Z_g���}��<�q��(��{�0��3ݛ�㪾R=7k��Y*����z�+%l䶎q������2�%i_^N�ya�n,K��3W���ZHK��u�S)(���S����ô��Ԇ�:S�vZ���9Je�d<�oB�4���[����*��e<<sVv�H�V��QD�_b��Vn�k������m_u����D��$wQ�p�KP]���gQ�)z��M��:|*��E�%>I^�|����zss���NY�������֐K�S%�U��,���]219�t�Y�R6/r�s͜��������A�S�,ddP41�ТV7��H��Ur�rt�\)r��RkvH�&LQ=�*�"�=׆<sm�o.�m]�T�^��ؔ���Mk%u��]�H��ν
�)���;3P�g%I���%�F�o/��˚v")���˷4[�͑��:7�R���c��6ut���Q��}�ӗ+h�-[�F���m�����q�&�27�z��K,��F��b�Tp�ؓ�l��iر_f���U�ts����u;4T��wH5\�5b�gɽ(�ĝʩ���/���%U�''g�^3��f�n���Î;��؜9a._k){[~�9�՗��ғ5�l��Or�]�	Xx�<���NJC\�$Grl��vN�*F�&✖�r]Rr�3U����m�9��5�[]���a�;ʹr�V�M:��1����؞�ekѷ����;�)vWR�0���N>1�i��mc���UEm��!U��J#��.�V��ڱ;�7��7و%�o:,�vұJ(�A�Yn��n��b+�78[km�9E4{޴��i��yQ�vB�Y��W�YŔ��+,�@��2���b���n˧U��z:�M�����n�?��6��!�j���{�WҢ��u�>�9�P��V�z��s�����\��y�N��m9*�ƺ�:���q�>^u�|ꓤ�ٶ�(s�"c��c{~޶�%��\���X2BK��2gNV���z�),�:�a���f��pي�A���8�i��ᜪ��L���f5������4�m}2�vD������n�Sv�4��/z�T^�����g1I,�f�M�$�0H��[��D�*oRT���V�7Z��s�ͽ����f��ʜ �Hڨ1��B�G'����m����w�u�WR��i뀨�\�d�D��:�o�u�F�|�#�@�֞�-7�װ��������T5���Q�5��&0�f)��TЊ�-�Ϊ��T��R�
w�����u[��v:�#uE�9u�*�@2�ٹ%��1�x�u~�m.�4������n5}�G+n���O�#��s<:%حv`v�r�t'6t��2�9��kɗH��.�wrͫiN�CO�)d�7�l�{)�M�.����k�9���_oD����Wu���"au'Mm��orhmtvˊ�]!�vJjNu��7\�Tk���YՅd�	�p�RH�\(�fr�;-�b/.�REf��èIw��[�#udfj:�u�V-���e�i#���*qU��N�2������n�o���+��6�]����+����+����	��4M���](kUApM��r'#�ŕ&�Y3��T&P�\�-�{6�x#�Й"I��K/�9�*	��[�:Iĵ�Z��^V�3���j;�w�Ӣ7R���%�I��\-I�x��$�1v�\���-΍>���������f.ٹM3|S�(�v�eb��IYk����V�!��&#��׹D�曾崤����G��u��y�-L��Dd�Σ�Nv^�	fO���yAe�oe�d��k&�HM�/�PcRU�i�]r�c�{���f�ld��2z[�=��+�A\�Sp��X��h㝊[����`('2RǵNN���s\�d�s-nn-CY�v�b�gPr���b�G:Q�͏��Y\BY8�؅�"��`�[�'��g�I���^%ԮNR�j�&5�">�t�qQ��wB+�m]��!�-;'X�7���9Lm��Vqg�ݕ�����"	��||�'	v�$�!��͒D=+��5wp9��>�j�T��n8�p��I�I6\�N��&�4Ea4N�$�I%�:X�4�N�$�NI�����I"t�N�����&tni��0߲���>�3#6jsSw��I$�I$�I$�I$�I$�I$�����t�I$�N����I$�I$�I$�I$�I$�I$�I$�I$�I$�I$�Hg2l�q��6�E0���=SשM��ښSF�cF+�^:�q�UV�h�M�iXWZu�޾|�c֛V4�4�m��M�����x�1����4�f%m�m+¾x��X��mZiX�m4���ڼ1��4���ύ�1�|mXҪ��L6��j��c�<~?i��M�Ѵi�����Li�h�U^?��=|��LcLm�Ɠm4���&�l��b���]=i��1X��UT�+M<m��x�_=b��i��Ҷ٣��0�4i��i_1�[|��M4яT�[OV�M4����+lmX�b֏���x�q�ξW�)�+M1�M*����M4�4�a�m�cm��Wνz�O]x��1�i�*�c�ͼc�δm��4�1_+m�㏞��X��4mUX�1�cOT��UZx��ͼS��>u�<>i�Ǎ1�6��<|��f*�<i���J�J�j��1�6��=c篘�m�PB�A80�c���[�2��B�ځI("3�#���oTn�J�M���( S��܂So["KV!>a�waF�����"��䩬���Ge!��Tچ:e�F�S�,ʷ2���ITK
�t��ca�b&�UPE7�y���Ae�C2P�f]7M�]��'� ���ǥ��"�)�ԁ��ى�Q�	�E�EF'��(��!8Z�%	�1l*N�I�I>A�&Rʟ�vX���-�#qH�a%G�~Q�r���45��x�	c���?n^%a�p��p��y��6��P�#�	NSIt�h��]�:��D�N���yAU�z����?B?�H��~�?�~�]�H�S���!	��bI'�O��d���������������=��J{J�J��w��W�]��7�u":ޤ�DnfMveQ5&]!�{R<��9��syTh�; �rEJ�}i�]&&�>�6r^8+�W�9	��P�ղJ�d����7`�\����-���K�b���r�5ۉv��!���w��W���?/_�&�RfLH �I�I\��/5�=��F��2۵��6'�֘mv�;A��9ݺ�Nj��)]�|qֳlL�G�A�,�8���К�p�He��v�DZ�m4%���wXF�W֝�f�|�z��ma��@�Q�}��{MCMiN���U1�'U�{�����kD�;���8��a!�[Ѵ����pn��D7Q,8ļ4�n��v�������15���LWy닏�w�F�1��90��H�]��T��=����XL�\r�Z�Iܳv�	(�K+*�$�#i�"c�1�M�"X���[(d�9�b�1u�c��aUg��d�U�����
FT�����K�\6S��9�ԭZ��R���B�0u\�Yٗ��O����\f��VƐf%p�Y���[N�f�Xr�ƘBƹ�V�bQ�E�vb�ؓ�+b���w.�j������YR_e4�˕����FNN��5����U��狖� �@h �� �:t��gN�:t��ӧM:t�ӧ�N��ӧΝ0�ӧJt�ӧM�:t�ӧ�:t�ӧO�:t�ӧL:t�ӧN�8S�ڻ��\�əʶ�mv�8o�_d]�xԘ�oi
�ʸ�*"� ��r}}�qi
�K�og���]���u^dLZ|j�\)ǉr��]u�Г�֩���R0k��	�f%�^!Q���z��.uƢ�,�W[SF�v�;�)rK[zm
�NSg�:�u���ukd��+�V�&�U�L�Dx�2����g^
'��R�hL�j�^�����������쾴(l�hjN]b��9�)pѫp���5U݌���"����J�yv���ꚸ3����9�p[s0[Uo�Iؗv���X�I$i�f����.X/�>�EԸj�4-����瑨@���\k^K�cřC��Y*ĺޱ�C����cCz��6�ĨV�cZ*�g,ֺ����Y��c&��T4��r�.�߅O���p��r��� ���v\�8t��Zy�Ԑ�'^�:ag[�̗��uQ]ש���A�zV90^vU͸_h���l�瞞pX�5v���Д��W5�=o*Iz��NmQ~2�}h���\�+��oTl��N�m:�ln�v��y��f&��9Wj�/�a�+�u�H��ް�'($����L�i~�utsZ�p�U��V+÷-r�n�� �J���sZ/�c��wk6�`@����ӧ�:t�ӧO�:t�ӧN�mt��ӧ�O�:aӧN�:t���ӧN�:t�ӧ�GN�:t��ӧN�:t�N�:t��8��b %����2�Ky�g,=j��uf����𻖮����C�@F*�X�2p�-�+s��N���@���]��=�4�R�Ny��[����i����s���Z}@��X����ݬ�0�Z��·�L."�I�o@V�+��
�;��lo���(�N�Tc9�>��\T�r��0��π��;h�w`ބb�Z|Cv�W������A��p�,*=C���
 ��0�1nY%Wv��$���U�4�q0O�?'�!v��`y�^�X3@�zꇋŖg`�K��]LS4@�x@C>�Fl=��.�ۤ��� ��H�^޽�x�IEc˔HB#F�x&���%��M{ސ�	^��2Z�7��a�U�����C�`{�r�	�.��hḥ�	W�}�H��-�=��\�����Z�j�0ryҷ��h���lc�	@�=���]�ϟP��@��@�R��-���I� ����`�r��V��3��P2*:���)�Ҋ*�}P\�z��hFu@y��z�r����u#������n,hډ#��%p�2P~T4��������S׼-�[��F* �0�LL�b�{�U�t��x���4�,��6�9��HpI6E�omX2�ٍ�F���/�� �@J��͇w3V+�7uM�3��}�g*cO��������	V����6�6+��f -R�y�6UW���/��Z0�>״+�p�2�#��`����
m{��\�c[<0\<�@�q��� ��p:tçN�:t��ӧM:tۧN��:zt�ӧN�:t�ӧON��:t鳧N�:xtt�ӧN�:|t�N�0�ӧN�:|tt��]�
���q#�L��tOAS#�g$�D&��Ȭꛯ�bЙvE�$����"��B�m�.�R���"F�ަ�}i�r��7��+�u�Η����э㹸�J�g�rv)8��D�����������Aݲ�\0@E�`����B[O����Z?s]�6d#Z�DͭU��fev�q��ժ�)�ur��+���eJA��s�N� U[qε�k����.�lP�9Ex�ݳ����h;�/�ޫUA`��(\�yͰ�����jS�؎#�Y�����
W�lk�-g;S��;���I��cpS!���Q��:���շ�1GW�]W�`;֮�&�s"R��Q[�Uݑ��Ed�E��a�����F�O{�-�do
�8��;CU�W�Y}k[gq9�/(u�A�eo\�6F���-u����?
��3m�꯻[-�̫碫M�����w6z�/h���Q��yoWR��!r�:zm3�J�-�V7�6�<����0m�s���֓=ǵ0l��.Z��V���Vh�1:�>��d!5uwD5SJ]U�*�h�-N�u(T�k%�X�T�;}~2�jMT,#J�!�oN|P�{u9�E]S��#��m)���8�G����@Z�s��z�Mq�;'{vM�o�<7�Pfl�;���(T�cr��I�g.�2.�wn���k�5M:xp��ÇJt�ӧN�:|t�N�:t��ӧN�:t�ӦΝ:t���ӧN�:xt�ӦΝ)ӧN�:t�ӥ:t��GN�:t����ߵ]V_9Y�f��xJZ+-0�["WSr`��F<��͗�v�W��Ӛ�wJ��(�u�~�:�(��Y�P�wM��YL�R_f��U�r��|s�B����E�f�����^��o�{yI.�F�����Jh�x�I��U�h���IwX�j��޸�/-���c�+�{М�g:�B<ԎpM_E��>R�ބg�Á[؃N��7
����;�PoU�w��%ܥj�}��m�&�z�6k�����ɮO
[��/u�F���8sR�)�;v9�JW���ts��[�}���Q;�*�CxEub]H��zt�[s8�|�a�(����8��i��Z3�t��7hQ���ܭ/Yz���74L�+�M䊤&G�j�����%Dt9��d�WNǡ�Y8�hdUj��Nb�Wh��^�D<p�i��H�RX��SH�h��53��[-�E[�&�؋Q�J��k��s��,�k{^�!�-̅���wv��k�|L�3�g4n��J�Mo>m�b%���R��篒��"�KJ2non��>*�Y�AΥ!"��,�z�p�E�fЮ��rqҺ<�HV�ҩ]��:Aa�P�/wG)b�uI��`X�@��çGN�:t�ӧN)ӧN�:t��Ӧ:t��gN�:t��ҝ:t��ӧN�6t���:t�ӧN�ӧN�:t�ӧ�G@k�.�p���lpv�����4qw��6uL�3�{gR]V�vg�����ZeWfP�\<��3uMC�[Τ�Io�ǽrp1vk����"��"ysV�]q�w�z���f�e����p�}���+��=WWk�1���l�C��Y��K�j�-QN�z���:h]����f�H�����b�uҊ�RU�O��۽O����t��.�	�@���$�e��Fҍ��ԇ}��Z���|����4��`�&�
��u�qT���[Au5�9|��x���΃e��1��0�ռk����DL�=0p�+(�E��ym8U��Yۋ8�-�&;7���JL��#�<D����1>'e�ǳ���*�y�Њ0�{��ȩQmQ���,�4�z��u���j�J��~��а���4�k�R�o��pL��!�`�St��\�_E���V3R�kZ�b�yT$_��\�h`Ʒ)�����mm���n�L'�W%S�{�G¤M+�*Κ뤬�k��G�J��-�Y��[��=V�:�e P[�Ku���2�A�52�� U�W��ֹ]�y�Y�)$���1	�C3E�O��u�t�zFWe�v�A���ӧN��ӧN�:t��ӧN�:t�ӇJt�ӧM�:t��çN�t�ӧ�N�8l�Ӧ:t�ӧO���:t��çN�6tp]#3�Mj(s[8��r�]D*)%\F�\�f���;���:/��V��s��*�J@�`wϷ�VU_s́fa��}�;�e��}�e�8�H��3�y6���i��G��MK��;t�E�����ٓ/s^��X�
��jk6��;��(�����������z�����o;R�]�]���x_n:|���vq���_K/���g��)�Wz�7;�[|6K���?i���eT�$�\'fL�2�wxCToo�˭u�<-Ru�qB��:��9�e�� ��zuX�!����;���3[�x�@��=*��i��Zx���֒�3b̲�򵲱���j�����V{r��8���T����#�eK+��gBQ�*����]���fˢA�\����a����P����W�0-U��8����U)?(��ïS���u�J�,Qɀ��[�F�_HAA4��Ƿ���]#q�F�֪�-˻���WwGb^Uʽ{E��˨u�~7.�U���_wN"ղ���B����&����
L*(�H:`��֌ѝw��=ᔑ�ƌ�G����z�����N34nU�����\��d�+��.t����˥3,��cx��$Yot�][��}���N=:p�ӧL:t�ӧN�:t�ӧN�:tt�ӧN�:t鳧N�4t�ӧ�N�:t��GN�:t���ӧN�:t��Ӧ��,���<{��Ǚ��*�V����m-�tN^+�ʬ�]�OVn���[6�6�>bW�}��'��TT��#N�����hc5v�R�+�۹��^��s�μ����IG��-��,�JS�rN^�J���B��o9&��l/b�d�5�5�ں���X���n��.���L��
��VR�'p��m�8#�B���R��U�#r��ܖ�����P�a�k���B�u��N&�-]Q]�<|�ܤ���ܣxQ���΁��y�|�&���8�q�{p�SE�Y+�s���@ꖺod
����^�P�jHS��̘��F�G�X��JdCi�6�^jr���ڱ���E���H(;��N��Z��T�q�kU�G]��cR�5΋k\���v*�G��
��r������r*�c0m�լK.���-h˥E���j���k�Z�庙&_=ѵe�D6��TS����QU�[n���.*}��y��u��(F���8�z��<���%4q}���0��{���]h�1�ND�N�풶j)�P�6*��&J���Jyh���bT�"�m���O�d�����z�*mӜ9ڥ���Y���]9��ԡ]��I�PkElO�Tz�残��0��@��8:t飧N�:t��ҝ:t�ӧN�::t�ӧN�>:tçN�4t�ӧN>0�ӧN�:t�ӧ�N��ӧN�:p���>�������7����2V5��J�-Ɯ=5����>P�}J�Ӫm^�,y��c:���/�DV)c��Glf��`��)��Zhl4�:[ۉ���Kp�xf fm�g[x4��B��v�GVm1�X1i�1g`��D�X9,����3E���!�-���ކ�_w`eO>%볃���+4Q$B��qH�D�՝n��ąNF4��b]�ؗ��=���}H����#���N�W		�
�o9K��l�S&�Fބ(�`��\�9�O8��Tu�ck��4]�-��۽:H�z\勵��;��0s��2Di�*�R�;�j�A��G�fS�GpV�Q-��V��!��
�WZ���6ͪ�����ܪѸ��'k��-]�d6{�fV�A �8��t$0°��.}�Wn�OB�ZUz�L���SE�6�.���n�q�p)c�;��)ml��gx)]�ъ,:=&���8a��a�P�\w8Z�Wx�"|���ÏR٘������(�j�\�!�N��ݫ�b�\k7o8�;�;�e��q>3P�١Y�.��2�.���c����r���оEu��Qu��1q�{��uQr5�I��W)�{�Q�5���7Wb
��ɋ�AC)~�Q�R9y�P6�V.{�R�,@��4��k��Gx8$��iҧ5�w�v; ��������CD��mQ�8[5���YW�����
L���S(Z���,������,�Q���g>x��n�ö1�Co3q��u����ottN�'y ��Y�a��1ee�۠����w��	|�Q�r�ӢT����ʊ�2�P�Ns�������җl��MKmm�#OCN��ю;մ�c����"�7N�z��}�w��Y��1���$�8�Eu;��qΫ�S��k�mO�7i���r�W�S9#��
�s-5
�^��U�!}z�pe�F���V��pVf��;�wy('�/��vuj.c���;�bM����m^;|�l�j��rX:���G���n��m���R��U+���[7;�(Ч!O"��p�'J������PUC����S7�����R���B�3�|�������ҙW���]q!���ܟ���|�.%K�qVU�ʎ�˽�7p��Q�S]kF�巹
��9j칱�l6���T�4�l�8л�l���-L�J��다�S������ic
v����~�����$�v/��������/���)?��I�k��W��=\��\ ��p��~AFc	�.�(�2�C�%T�@���O��t��cG7���Ń+"eK�ǘ�p�k���}v�ekC��
$��1��nac�"�1T�������U��us�ʦ�:��v���}Ӎ)V��0L3/x��r�R1y�o_>������r�_n:[)��˪��x�;T��=�i�z�Ӵr\1V�u ��9��y*�j�O24㩁�q�Ӗ��7v�(�-^�ΡAu$w�j�(R��*\ܾ�����4Uu��mZ�r�Y"�!��XY՝��tJ����N��v��yj鎅��6�:a�4V�C8ΎѮ�:]�R��֮B�Ň;r�vR틃gb�N������wT�M�Br�M�.rk��BD%�s�:�u�R�/^�|oqcEw8p^�˶p�a��ش�ʝK�$6��3���y�x�j���Ra�m*4�Z�Q��� �u�[��&����5��)���}Ww���+�K��z��C�S��|�`���E؂b׍���od��]��g�*VsԍQˬ�*�����5�I�]޹#S'e�R��upķ4��]�Z�n�>%ꥰM6]:q�'U�OfqW��4vΐ�4��鸻��M�F�I�I���c¼b�xƞ�M6�cM8�Ǎ�G�6´���4�i��hٍ1��aX��±�S���LM��j��J�<iⱍ1�M���m+��eL+�֛S�M��z�tֵ��]J*҄REF�e �m�q��R4�lp*(��;e�陔�T7m�)��I�A�h�K�F~?��j�戶�n�_��Ҕ����p�ӝ��%���L�{g,{^�<�(��ԍ�2Ɋ��{�*����1KVU���:t�*�ԋUKV�I}[n���V�D�"��������R���{u��ʵ%�DJZٖ�[�V�X���k�uQRQ�F����"�K)d���aP򤹅U�b����1*��^֋V���:t���ӧGQUB�ijʪ,Wl�U�YFd�Z���7EK��J���]�;�y%/�%��z�Բ���sX�g,ªҽ�*����O�9�õ�Uh�*�,��d�u�<^y]��v�颊RR�c�U5�#�<:t�ӝ*�\V���v�ɒI7M���r�UΚ��KWV:��F�V�Xr��`�����ӇNuE^��F[��ҿU�W���)%Mؘ�1eW�}e��*ʣ�����:~�Y�>�vmwS
)�^.�K]�������W�T���,�SE4zt��ӧ�uO�NX1d>���oq$�7G�(��T��S����V�
(� ��{��n�ٔhP�A��7>[>��QN�T��c���$�@���x�3ԉO��S!�����o�P! �C�i�Eca����2�ݹ�bMio�/���F`������4)��X���2���'��NC��ʳ����3�V�}4�X�[o�*|؝�� 3=S�lQ �i���	�Cwni< &�1��` ��V@*�S=MWV�_�vw�W�#�Un�7�+MIO�7��@[�u�JP%��ŦT�j�{����� ��G,�S�ن<HW�օ�{��E���Y�{uV/+b%]j/{hg�޷cwU�)VHb_��\��5�Tx6��)<�����[8��^�di�W{�5ig��� �
��li��J�=�^Mɾ�w"�k!G��ݰoq�7����袝�z�����g:�f���'�w�	�5Mf��>�S͘��*���D�_�+g���Y1�h��e�[$� 0kQ � �z#��ٞk�>�唾���,*�q��Z�f"vb�� �f�1+7$Dx��a�KVa�
_��m��]���r)����U�tDd�l�_w�����k�cW&��Ϋ]���R��\�$1mҹ���5o[���t��b���՘�;x���&��be	��1,&��F#`��e���@SL07�S�>L��f>���D�.�J�2�T��hD�� fdb!�+j�>�Hbĸ�mB-c*Sj;������d8���V�i������J�ce*G���1��П8�G�+�
�}��ki��S�^ЋQ�@��YQ��!P3eK5i��<�X��+K#T�����/.���^r�8���>>�K�|&��l��U�3I*�4�=@qw�)�0���#�'�R��u�bz�n��|Z��(��(�|�&�%s��`�Y������2�{Ҹ\J��"��%կJs�XӒ&���6UT�V�l���
�A[�����.XD��̓G6��:�Q)j�V���j��lj�l�A��y�9u�uc��j���#�O8N7n�;�:X�N��c�AW�k���wF��6����H�d>��
B���I|��(��X���в���%����4��҆2�e�}N\�`��腷e*;�sU5��a���54i�@�%�����Y#5�Y�䑚��sN��FH�Q���T^;(�d�S�m�^.�u��4b͖�U{�g����ǩ����Od��QT�m��!��BY�	.�М͑R�����.nv��V\���}^�1cG@�-{��ܘ��m��3xآH�	���=�x;xlc�$4�<C`K��%�$�T���c=��6x�i�0.�5��H�������b���4�ɽU�.���ސ����}�{%|�'��Dj���u���@k�������[����6�N����p�t� �P�"VV�3r���)7WjU==e:^}�o�m�0V�}U�U��`�Û�u/�}��J�5�>���ދ�؜\��/�?9UV1\O�akP�ҮD%-�M;�����745Lтɽ髷i-��ojZ}�]��G��S�fR�#��u���G�窥 zĨ3s�T)���P��Ջ����7�uiU��:ZYH���a�݈u�����?HK�h����߾U�w���˘ҰF:�ڜ��C���ϥ����u{��]f,�k=F�,l���~[�S���/K�ϓ���}��皇��UR��@�+�U9r��FްFD�9u4���D;C�db������Ml�q^j����U�/e��M��j�H��ie��MmE��'�m���Ej�|�����i��Ό����c!����u�Zt8_s��}��>��Fug�ؚB�M>K�͐)Z�T#i�}��A���V�i�>�l���ɍ�Zʘ�L�6�n���ҋ�"������9Xip��|mA���h5ZW�NH't�4��@�����O���.�)n���w��.��M�$�L��>�+�HM�t
04��_jj����E�5j�`4���}k���m�h!+!!�]f�<��oOu�+e<��&���=/�}���3����#|�F�}�|�issR���s�#�l��(���B	n]'V��OUΧ��f��[D�q;ݘ+���Rղ�,��gveb����rջ,�۝j�}��v1�� @Z|i�+l1�G�K��Z���[�l�#&�S�/ۣ�W@Xq� /��gʗ�X9�Vʜ}u��3@a���"��E���2�l�1W�
cg���Mv_��ŀi�V|���&$ױJsՑ�Z�j��V`�Ԩ`���K�aܗ��k�,\>�=,0��謣��H2�,l��챽g*t��I�9u�O�Ab�<��~H�y�l�EF���dr����{
�'��*�q�7}��ry�+��d�W9��E�w۝}צ�f��8�ݾ~)C^cۃ����(�B��>4�FA񣛗ݽ����z�X{�b�"-�X�g�����T�U�$hN<=Y�t������5�f��Z�Uݪ��Oy�K��~5�*�ľ�n�Y`OR#:\��lV����k���p���$�g�en�7��$���`S����.�.)=T=sO@h�\����.��������D�:C
e!� ����zo7��޻��z¹lc|�^
S���8��
�._��ƺø��,p6����CL��3�[ⷹp��N9\}5�Xy6>B~:�:g!�f�w��7�����V��%z��ge���k}y{|�wZ���<��.k d�֢�@�^/%S��	^ώ���vӉ����E5��f �@A��h5�l`��"�E0�ʃ��K�|��mj:q24�%PO��� :]�\F@{ٛJ��5��B(�)4���d��Z���7זX��t׽_���,���ǳY�^R��a1&��¶S���7}~�1��{[>�����,%�{s�]�{�q0!E���B0�b�7�$#���d��VI.��峱.D�P�F�ȱf.� �^�L3^�.�5����U��D�;S�tP�e�y^j����ο! ��}����}��g,�­0�umvh��QFz��G�2̦��xD�E����*sf�ً�	Ԥ��=r�W�Pｋ�h��j��a�uF�ƾ��id��5���U�+2��S��c=.;�^{��K����ۈ��q[���q��=�܉Dn�4�<�ՏE�F��V��0K��c_r���tI	���Γ�1:��T�e�K׃�R�@F�K�*���`A�{��.��B܌��s�Q+�"5"��ʠ1�����n�Ɩ[d�'|�W��Vb��*����Y�]��<^6l�l3TD�QOcm�ĵM��+uҵ�'&��R��7x:f����(�yW�0�76[s��� �)"Jg���Z8e����pR�Ͱ�4�ue���͐31�K<����gi'��cR�#[-n"�Y!��N�m0�h�ih�,�m`E�ڜ���¶|>����ҵw�H�����~���o�Jw45LK�&�/��v��B>�5 �7�Py$�8p,;mǝf�AF	2��� #��\VN�.�۟lV/�'�'K�r����{��uLNW���W1K�Zr�Un�Ӹ���`�n�w�=;Rʱ=�O������&��b��Ҧ�0;��O/���6�x򪪦�]�_'�QL�mD+lM�У�(
���^ca���R�e���i�����+y���ܵùv����u�8.t+n���e��!���J%-��s���롻3�h]���X�V��d��@b�F�K^2��%Q�eBJp�B�����}���'l�CC~d������}���(z��^x}2�h�O��*�%>^x8o6+?]�a݆�B2�VыQ�f�[���}� �5�W]?��^,ļ:J����&\�,�M��e���1gi��4��|�L<  ��5ዑX;��o���|W��¸y17�7��V[ے�I=�U82�,�op��zƑS��LL������#�[>J���K@̻�"�e>){��$��ȣ���qG��g�+ba�~^@p�PQz��h�wݡ}��ŝ�#h9.�o��� ����[�f0i�7r������G1�\�L=�JQ�/����տ�;94��Z�J����}C{�f?��6���:�s6��y��B���OS�p��Nv6�ۧ��͗��LJ��˸mc��M]%�b�l���_��ɾ�� +�?�@0Y%��I�����w����I��i����ǟN��\36�h��D���n������.����	�ۥo+/�>lڣ,^�L��@�!b�6�f0�e	���d��{�p�A� ��Y��[�`k$j���y|��5�ysy�H�f+�VU�b�&+uN��dl���m�����a�/�]*f�w�rwa��sf�Q1X��YIn�Z�4�����Iw}Y�ׇ��}����o)�k�G������Dǉ�.��w�d�o_w$�~�k�s�!���׭��S�Ek6&zS-za�$�R�Sg^�ٯR���/��1���
X���f��D��ͥL+vlKM�e�7
I.�@lf�/q��dH>����N���V�����N��U�s<����B�c;��5��1�j[����?{��B��5�f��%Y^�E�N��7�#��X�o�+o�uv������r�'���d����\���zM�9���WY��V�\�s��Rbub�ws�vݤ�%��\V�w.����s�ӕ�]��o�pJu۪xq�2,����4�M�QO-t��td��9r2D�ˠˮ�-�s�'�I���GH�e��gt�e)͠|j�a{�؞����P�5Lʁ8��?ի�38jke"3$��d"��v+3r�}mW,W����H@��>�6���<LVF���N�ES�^Q^+i,{�^@l=�@��M�J>���~~p��4eV��-��CI���T��*�}4�ה	̉ʘj�x*�UJNovf++}�yD�-��,$"˫E�V�͆�Uߵ^ρJm������j�0E��e
\�B4�]�����za-eeM}�m;�x�PWMԓ�ɋ�>�d �P�P�sk��%�mT%�k�ѤU%F.��_t��/�#}�����	�}�x}�����t�)��%Us�o*s��a~�̔Ж�"*�-�i`����s�x�25��
�~��]�|W��mAG.P�ĞH�~������,{��o��	�~T���#3��h��0sn���ORU�	\�q�V��a��-�5�ik�7�v��*�Nbۊ��%SO͵9Z\۹H;���;�̩4�Y}JX2i��=�ˋ]�&@�f
�I��yj��y�����E�}kr&e�g�&�ǶB���cmr��ڦ:��7a�^r���w�s�Q�������!oz�Ccr�T��2�ɸԒkX]d���\XB�;ofcjr���T	M��(�X8����K�y�9�W=Sqξx�{��5�Ѽ����1'y�2����3V�tr�%Jr�iew]aeP��G�EM`�F�o7���RÈ�[egh� �	��X*����gVd���=���c7�9ݺej|�6.�f\;��S��0��S��&�<�s��9�N��xz!�nun��9�����K�.��k�fO�;���:��B{V���\�rT����W�@�E�/sXt��s���բT��
��b��@���ں{w^fv�a\�c�]&��M�ә���j)�m"��j�����yY}m3�ټ/e}*�Yrkx���J]uUI��5��b>�)�=�\�QyU���z=^f�����[����G"�Ϋc�j>|ѻ��*6z}R�,�Z��f����/�klf�V���.�Le]4��[fm�7W�6����ygϰ�cK�UjҪ�Ǎcni��Wͷ�3��X�ܭjy���u����
8hv4������� �l"4!�������;뱠���}]wjz���n�<X'$�jĔz\�uj����4�#9��;�L������B-Cml�Nv���9R��2�o����S[�]��|p����%���MYt��5���Y��<J'c����3@��[]m��L�5b
�q�z�U��t�C�'P�˒����K4�aT3�uE<�E]q��!��["�c��u����ȴ�2��VL�wƆˣ\��'���{ӗ�%,!�֬���7�!5�˦	˗|u�׏�u8��c�#�v�%��cdw���u�X�1�5�
�}���PJ�M��2�R��*wqZ榬��J���eX�����&؋��Հ����[,�)�������ur�3'.ns�N�:�������,�T�:v�ة[9mu*�ΡͲ9\�fb,���щ>+y��]{��4��7םJ��qT�YD�Ќ̵��5�gvU�ɪ��x�Uܻ����J�����p�[�[���׆���MQƯ�(Z�f�����)��)�����ۙ��w�S���;Ksp)uUk�թ��f�Vt��9)Ʒy�*w.$�wH邏d������/��k�ҏ��~3��C���j�kzk�j4[zm��6�I�h��f�����t��6Re5�>Y+�9d�,��&0��OON:rNY�k�(���OVC����r��-7g��1Ӈ�N�82��{�&��؞Y��u���%��:t�K,��<�e/q��j�̲=�<�7I0釆�O��:|;\����֪[-yQ�=�I�+V�飧�:t�qyd�{�zk��m<vߓoƍx�{dʔ�͝=:t�Ӄ��e',j�S�j�_�I�����rϊt�����çKbN�Y}��Ix�m�mzW75bX�I�->���Q�ؚ�ґ����u�m��f�Y|J����ؕ�I��T�:����gjf�:�el�+ѽ��G���6��_m漸���e-*�KJ��䟟r�s�0�s~�71��#F�����yN�U
SHu
#RT���c���*�g�e<���[t����?�������4vl�������&�֏��1�N4:�}}��k���%���0�=�ٳ����w��;�U���?�>�g�` �=�Y��6WF 98�t0�-��2�YP��l&���)*�K,-���܉ߢbP��lQV��+��+Dz~�����Y�+��գ ��dջ��,X ���������\d@������W���呂��d~Ɔ'�ud����k&(Zf��2;�-�y4ɻ̶��U�9=��Ļ�]��,�C5�fZ���Q�����;ɇ7���x6���}}���)�G\�[z-.����ܩ��m��e2h�c/w�m�vc�}�/ � S�`���k���J�u^ׯ�kP=���G	ܠ�+3!ޮg, ����5������[µ���p	�r{�uo���@W�ג��M}�S ƋoHg�����,W�������~	�ʐ�6;\��x�:�Q��x��y9n��=o<7*��K���S�{����Z���;r��U�W����o��=�=��S�i|�	��5�)�c��S���\v�����G^��u�/��s�d�i��&��6�egpڎ����~��@��R�=�
V���������_{�Sۧ���\|h@� iH�h+c`�G�~b�$I{���R����(CL�X=���?~�xD�l��(
�p�d��Xg��'�`=/%�xY=V�QӲ��Ib�V��@�3��&�;p���S�2�q�S�Y�뢤��yhfmѱ��@�~ƶ{��w�{��� Q�����c�<�5H�@ݕ�*�ȶ��.#��!\����Q����k+[�ݼ�]ر�PŚ3xj�yN�.�D�}�5q����+�z�I��T)L��*bas�>�78������%E�Ng߁G����P���sc�cV|@�N����?��t!���xw\z����
#r!�?8W*�Y�CM���?�v{�yM�S��(_k���5��^Νq�o	?5�7�]��/g?�|��u��Z��`	�`[�����\�l�������|��8�a��t����KHC L�:��d2��rB�Ui�f)nL_��V�yz�)�WE��ض�2��Q�Ī�7�m���q���v�'�g=��78�W�(��Vk�P��,%9�N��R[.��S[ѕ��L̻V�N�ُU�H��̬l���\��_��t?��2G/P�+��q23�򐽺8�O�Y'��_K�;�k�.�2����s:���#α�qo5�Z�p��np�m���ٶ1�����������k2���������
�Y�)d���)P��cϳ�~����>���?x(h��o�&}��o����� ���q��h<�NĊjnco5�I��P��q�']�c蝾i�}$�F;����A�ϩٍo����\vx̲��ʳ�t�w@��Lw1.%Fs�Jũ�e���n��Ϯ�+,��~AX���5��f�wB��4`o\ٜ~�'��at7����8,��_�D�����aR����kA�������~=�Y>4�:�R�����pXp1ͥ�9�M׽%�wOc��Zrvn\�y�y��bw�[�8+�.�w��ܴ'p�BiAN(���t��z�A�;:hrԘh�p�fnmWBe����WkO\xF8w|��xT{b��[�S��\�����0�֩��s�g�:[�V~��I���d�_�(��2���s��/���X羷~B)w���-���{�V�����%�ޛ�rx��ZO|�|BMr֨���>A�Vk�ƌ�+3yn�yk����V�<���y�s�4u���A��4�O��
��'����������Z�Kn��Y�`���n�l�l�]r���qBw��Z�d������*lB�r�FAbz�m.�Y��vb�W5e���G��v�֊�r6&R���XoA�!Pj��u�ѥr�/�sZ���H�0��Y#�
Y�"�"�C�d[$w��i[ܸA��m� �Ռ��� ��!*�<�J��D;A����?OL�>�h\�D���n����b㽸�Ɇ�c�}bt��q��������� x�G�[6;щ�]�!7��/��V-���zF	N���>wp"���E����o.~��p�!+�ay{y1�d�9�O
�G{����V�*���28ȡ�}?<���`&X	��J�-z�	]<��r�����q��q�Y��ٟ��K4І�����������1~�q�D�5{������ӧ"�oV7��]
�}����ǔa7F���Z�Fk���$��c�,@S3-[�������+��c�uS{Ίm��XE����~�f5T��*dsc%gd o;tw� |ޅ�'"��ss
�y���m�a :;�;j�B̅Y�e�����E�Y���bM@M-��*;�b��y�������8v�M������tЊ��'����e��;�Axe5қޛ<�E�OJ#Yu���f��3��m-ʸ��r�`��]!�$���6򕦢V�<�,b���7s�୙�{��Y�IC���{�u�I���� r]wf��1�O5N\�r��R�Rœ)P���+]˶���-$j�I��=�{/�I?E~�-D¤���"aI))*H��R�V &K��x}r|͟�Dט���#����~H ��~9��>l�Ńo��4-�.��z��N �y˽�9�Cq��a� sP'sX�Z@{����U���t�ŤF��nX�xY�F=2-��xZ��6-��3L{T�HD\�Jv664�!�̣��K���Nr�7�\D��7����tf���E�1�o��T��fƸ#��p|��S��VW:h��c޸�`��~-�Us��*�����@��F��Iw��]�{zz��PCV�"�&�RꭟF���ϼ	�����5��vl��^��KV�@ �Qq������9%�)�==ݟJ�g�Q}�%�%�D��ɗ��`8��ד��]�`@�oB��ì~=G�d#�2Uξi~I݇��۶�lg8�%�ې��;"��[�hpy�_�/,6�)����ɷBٜ�]�K:�~�g��Ji��nq��n��u*��/]3~��b��ڃ:��I�[�(dj�Q�1ul��N3�[��6����2e~+k  dq��U���Ҁ���r����X���o�e{/����
��*�rC���=\f{ȟb�|�/.m!}��PI��
f�G�W��Uw"�����ENj���(FE�A���]j��5J���pRR�:͐o��S���l���-�/�W������y���RO�
�Ց��Ȱ0�$�eI�h��&��I������=�,�x��@�pl�+|���G����)���Sm��{�Ӎ7���o6v _�>i�(N�?|���|����_>㌆B�K���/h`νa,�[�j��?�7*ѹO���B��l�W��1}��� ����_�I���h��������Es�ٍ9�ɅΞ��Ƚ��ʹ�}���n�ܡ�'*w!\���J�M����]�}���6\�X��Q�y7{S�g���7���c�45&��+c`��&�� ��-Ly#S�l�f�1-(Ce��౽~욒(Rg�
'޾�61�<���{aѥ�������z`��8s)��ymk��H�PXz��:yi�b�-�!�~�l�ٯI�O����u�O�o�<����k�8��Ɣ�gÀj&:�e��41�ѐ�BUk$�ɟqi�k3!�������	��L�^�g��A���W4p\{�t��ص"}���L
�T�O��=7���zz��t��_H;�U���ٛ;B`��!�;�B�~@c'o��=a�Eܨ�<�3��VM�R���Wˋ��������J��9^A�dp��������H �)q\�Rf���su4��u���+	.������$�9s-������/w��V��K�dG�숎�h���>����Q;8>t�4���xƚa������u��b���,HR��)$�I
Y$)R!�3�եo X!�
�ユ��z.07�k�y��/�r�& �����t8A�_��XH1�y��c�
C\ «�V�G3v�����u��R�3n�&�y���@��Ll_<+�t��h�8�qM޻����_��<x�<�ǤP�xga�R�w�0��=�[�{2�b�� y�3��7�#דxDjV7ލP����=p���Ꮈu�_�]
�3l�4��DC�G �wK����t�
�9�Tr�/�s����{�?Z�`�Lq밿���<7���\٭8=�*Vcߎ���߆{)��G��lZ���Y���>^&+<o�=������ύ>���f�M7/����ˀO��؂���D=)�_��5dPX��}0�k��lpj.��5�g!�2;M5j��)�\�s�QM����� =k0mʛɊ�N�m͌�<�I�Gs��t�u[Vl�xmop�n�RuO0���_����;�ZAowO����/܆�� (6;N�M�v|;�]��&6'����W���r�zA��F���ܨ��;>�#�kC^}f�<�8�f�?��<���Kb��b��p����^���u���v��WE�nE%��̾W(��iU�����C��OCB�\C���,��-.�!�������Ii��6���=-0�v�2�.��d:v��[wv��3$�-��$1c�5�܁�,$R�n�L,DR��E,"RĉJ�H��ݚc�wx�|(x<kux���	��ή��|�]���W���\b�L0lJ�z��l�M3J��n���8�� ��gL��<C�|���笒@oGK �_�s5k2�]}�����vk���']�2�T7���{�{X&������|m�ɟ�Z��r�jw���n�q�Ǡ9�SB}
�%"����;k�t
�laz]����14�r�۬v��p=8��5����[�<Y�ܥ3(�w�Ȱ)�]]Ǚ�30����� s������<Y��\� �O���,8����h �V0iJm�����cx�1�-?O&7k�`���wA���Y�VG���aπx��1	���J�᧌ �Z�����5P�D�A֝g��8�{-}���|���G��,�T�Z��'�pZ�M7���@��C�>5!2�%�8�k�-ȫK�Y�F`���ȟaP̪��ۦX����S��>2��E�������,ʬ�Q��|[�]vG*�hw�a`&�HA04�{�^ػΐ5�����k�![Y�
mP
� s�'��Y�:Y�[��lӝ���=M�c�g��v̬�[>
n�찂���|��	��9%Ẩa���� ��\��z#���5RM��W�d������2S��m�/�	K�Sf�P�ެp��Kf����oY��{���H��!)RB�"JX$�)P�Y$0�DШ�)�H���]�~�;o���Oϼ� ��sv��M���+�d�	Ώ�Sa�el�d_�ÕR/�C��7Y7������X��ܑ#�qz�?0��u̖��SetSc��6K�q6����0`�,3�D�[���]"�&�V쇟�/�5�TJv��X���`;�[���㷄Mub����:�VP���64�Cc�O�+��� 1w\ �k'S�PQ��S �*�Βx�����">kmY���#Ʌ��;@�GO'� e�9�ة�����Wl��{�(���qܓ x�)��æv4���׳�$4/�@|{ʄS�ƄP鵐g8�]ΛɹŽ;ܲ5������%�B����hrd<�����X��;_U����gߙE���b��p�]����$�]}�}ل�q@p��uD����e.�c����a�p���H����_YNt�����>����Bo�C;�Csb�b��v��U;��xf���A��qi��o��ڧr� �f�8�{ŏ��g�&�<y=�%��9�y�J��+_h�	UK���M��7�_;�;\���RX1:�H��5�P�ϐ�v��AF>�M��p��8�
�[v����aq��s�gDIFh��Ҿ�; H��'C���n�ez˷ϝ�z�]���ݼ��',D���I���,H�P��R�$ʑ0�H)d�)d�������Jp��=)�^�h�v������� @x�3z|k��c'�#�Ƌ��6���x�/)H���D�{ZCU�����0/uE򱃙/�&#��lQV��h�~��Gw��Bv1����-*Uz
W��w�-��s��������oD�_��D����*��+j�)�g�Z�!�%�K�4��Y�Y��P<��P _E4۠ɤ�ndVL�ovP�Λ��,�c��:�M�+,ع᜸�i�P���JU��>.� �+֦/��W����}�l	m�wM���Ս3���>���<l֏?������_� ����}��\�dH��q;*Q{���K�@�gr*���B&$�(ގ ^<0L�Q���~;�ed1����9)�,��6���.Q��+E�e��"�
�D�-�����3U���(
�����m�ho0�;!��v!�������f�Tm�[�3{���z�
�u������Q������XlA��5Da6���?�3��}�Ϸ�Q{6Z�g3�kX�ށ�i]+������?{�7���V�����T� �`��{`�=�x8D־�޶聱wٯ��j��5^�9F�,!%������\��T��2op]ْ+�Z����|�,��9���]aX
�r�.�V���=qn��\��N5;zQ�^^������V��_#ǈt�/��]��V&:-����5y�Lh�<lB��gt�s��A�g\k�{�Y�um�n�7]&<�cRrA�v�<p�G!�D\O*�ח$�rfu�ޮ0.�C4�H�ӫ������uS:*�	��L�-���U�Q�w��G��oC���5�^�+�5>�g)�3�o#}|��[eaΡy[ɵ��r�)5ce6�u+08x�v���*�6�#�2Q���=:swi�>\��w3��gw��I8�KqV^�Tz��wV��5V�������s�ڲf!�S�ُsnJ�j/6j�%SV���.��A�0D�TUJ�j�o&▍�fL&^��Q	����z��E+A�bE���gt8rm��b:����}:�I��~rT������9JՊR���4��)V�,��b��>�'Z��0r�鎺<���V�խ5���0�e2�Ռ:l���s�I��)�A�g\nW��YV9{�S��f�t�Uv�Z��]��F�s�J�P�r�ue�&nuI���j�_8	����2.����;kFwB5ÕeU��q�I"�Yߧ	����ո,�P�A����X(X&m��#�Ċ�d`O`�P"�@E��`b��b��!V1�V!^M
"�:�`X�C�e�6Ņ����^�Yu�jX�`vX�����cA qo��X�[�2�0��@��_�+x6�c��>���*N��׮��v�� ��;EUV7n�a���ғa�����\��T�̳�7z�쥜v�P$�#����d�N�Y�1ӭv^<��l��r��U��-]�s#���v�GA��ۜb1�]R9-�x+EB܅r�WJ��J.��E=�.�*�qu骛�	!W���M4���l�4����o��R����D�����kx����ބ⮺�|/�UA�����Y�7)s;ܛ�7�y�5n�N���M�V�/{G	�k�ٳQPɹ���QW����x��`R_7�l�ƪJ����N���ڵ&ʪ�1��޼����;׷�z�4����y����íq��Nd���د@�ׂ����*n���
��k��:�%��fI��ܫ���E�os4^_m��u��zv0e���NK��Ŧ빤\�o�r��-'Ԫ�R�P�wV�Z�JOP�j�xb�uLA�N��5v
W��ʾ�jBo���WK.��9��J�F�P�y�J�s��띮ٷ�k�y����ׇiͿc�tR��*	f�ӲΡs���v�iUt�#?;[z��F�ӯ�k����n;K_u�t�gU9\n,lL�#���gg_���r���Q��/�{����jww7}$�$�00P�(X�A
4c���ϕ��T�Li�1�b���+���6�J�ƛi��i�W�ѵxi�*�O�����Sƪ��׭�z�X��A)<����b��k���"�IK##k����]]$�W;,�D� E�,��qB�V~��?�?���
��|m����F�o}�~ur5�8zzx~���ڞ�v����nk�&����^.mzU�m�%������^٢�=6z|}����~���V�M�ߋsFM_��R�<��MYJt��çN�<���V��؜�Ư9S�W��ƮB�O>�����cS�Ț��fb�Xq�D߸���&��S�����:g8��-Km�^���U���v+��+Ʋc�d��g�>���3#*C�k��m�����x�ܯ��W4}O����Sg��p��8}V��7�~���t��ϊܬm��1c�u+��^��}���_/���ڍI�+�W�k���77���۞��F��4n�R��/��m{oB������O�	����bTJ���m�+2����;U�u�jwo�w���U�W�ٜ��t�h;�[��l�V��glL��=H�:)q�Ϲb��X��
{�J�i[h�M4�J�Mf�s[�o[f���ֳ3'��O�b$�H��!KI�(IK$IK��0�eH��$g���q���B �~�H�E<�� ��
��%�U�1�Y��+�5�!��#C�ov��Z.
U5ۯ�xc75�h��K��Q�<��N淥s��d[R0�Z�A(�Y;��jI�o�)�-����᱾}�gN�;��q#&>�6���`mfu�7C�U�j�ޔY����l�_��,=|�0~$,:��hT��'>(Z�a�,�	��\3[����ۻ����X�|��'[���xy�v������D�I�Wȁ���o����S�@��'�qm#:;���K�b�Q�Q��x@ow���)�y2fk�h,���A��wXc̀-!�^E��ZBP�ՈR�F�xS�R*�5v�?+��֞(�]�?V�Lx�ڲ2����q>S��0����W]�n]������ �&T��c]�)Q�:6�N��{�0^��k#NO�__�Y���~$a�[��`A,8��Dw�Iq홞i�C�6n���B��T>~�~F6 91E�e�z�^����0�]�U�d��',9��C1��h�ОQ�������E�#y�2fɌli�FȌnQ�
��-jGuq�Lu�c���ncޏM��ڝ/#Y�;"�E�3>m\�O0������,!�V@{߈ �3���<�f�wY�8�\�J�@�{�COTgV���uw;A:,�/v�Ejp���Ԏk��r���q�������T&T��BJY)bI)a�)d��D�~i����[Å[�:���+αz�=ٙB�\� ʎ�$?Q��y�L4��`�����^0�=�Κ]	_<8f�^A�6+es��-���t>�c�|d�v=��M�Aar��{h�������2c',�Ӧ<�3�)��7� �RM�0���K˚����#Й`��q1ѭ1�"�᝱�G��l2�Ҋ�����O f������<��P)?�N@f�u�F ���w:��w���{�.r�%�[�qx��)� gL�b9���t�-�G�^*^ޙ ��.�;������`:��1���X��xǠ)�d��;7@Q 1�	k�=�r<�P���������6�G,�W��kN՝�W�K{��p=�{hn��y٣^D↚� -"�x\��4˝�ap�
b�u��[ə7>�k��cz>���* *�����ސ�=��c�o.�w8���b���/ ?�����R�S�=����G�)��a�!F�(o��<L���}!J~��2�}M���D��mS�����1J�j1�,�ba�]冿c~?�P�<��n���X��#�]�?tS�N�~1�Dfu[�-7Ҹ���;V�phP�������Z�ݶhޢ�:����Wڲ�@	 ��D!)�-u�]4+'[��%K�O�sv���In%. �.#t�z��±%�)�r�=�q�5�uA������y�s��ǫ���#�YJT#�
��đ�H����$���&,"MT���<���������r�~	3�x`$5��*����>��C -pᫀx��i�6��C*(LMۦ�z�ʀ��ED]����0��W
�����@exю�|�!ƫ��Z#��gW�0�ᗧ�����|���V�xy�0���[P��]Xt�L��b�KT� ��[Ipi��3[ݽ��j~�@��D<S;w`J�{h.̱w����C�l%v�K�f5�W���d �<�x��~�E��W����~����W	�;�U^�T˞�)vV|���1ab>�5!���^�՝��.���pK���A��H�Q(�^S���O�u�ȶ�)�2��uТ�b.��S�5���[��� J�  
cK� -}������0����}ktx"�$3��@F�J�u����NZ�k���ǻ�;64k�<s�����3a��u�L�������-*���\D�q�(�'ǒǬl �,C��8��z6w�o���f!�n�h�Ѽ��:`�c�&?��}a�@;m�u�a	|���%>4��XKQ�%�pq�Y-�P����,oW�3>}&T�ji�2t�tg��л7��X���cnϳ$$�B��8,!�+_u�Fܙ@�N�����Y�jpM�8�5�V�nS��D���e�����k���`������?�ޟ��%(IK!%)!�F"JT��I&X�����~���4�p=�ɷ��&���F[�C�W�(����pN!$?~ 9�Zށd3�3�H>��rq�I� ����6k�Ǯ��zXg=N��/�`�����_L�t�q*�&����٘>l��}���4hE|$��������b���*Ň�l��(�Ļ�g� >~~+ν�q�1oƳy*����r�v� Јf�c��P��>�΅i��g~��$o��-�^3baE*��� ��P�3fj���W(��Q�*�3'��v{�'Ţ���j[���ڭ�N^h�U�.<=����ǟ�1�.Ɛ�䮟��vm����yp)�E� z"j=FT.�'��I�KI��m���� �pǃ3Ǒ�f�%��{�����;M�Ua��C�61�6����׽	Gxz!�4à5�.���׏����x@��S�ˍз1�#@�:�Ap��&�z#�hX��'37����͞$9��	�'�ۍ� �x�;#�[Yk���c:D
}�Ǡ[���1���mzK�CZwbx4y��5�xP:\5��F0��6,s�!3�M�����t�S���F)�5e���#=����9U���MnU�ӗ4��ܛ�8���{'���@��G� ��Mz��7Eݳ�#�ߋļ��PTD(�³(lhsЙ�z�mΘ�sww�U8�g�j.]��aW]#�6��'E�<�&WA�OJ��..�+i{G(P�DX�A	�k1��z��^˗5��$O�PJY$�RH���Y��H�S
�R�����=�s^���{�?]�X�D	�ƙ�~З���#�@}�{_�Nȃ=� ���-��,f�����c2ӏb���q -���\�{�e!ڹe�r!��@F���-"-�������mS7Ym�6A��3\S�!�u�f8�,�K�1��������I���&���?�^��8�ؾ~{[|��`/��ŷ��ڍ/^��nnF.�:�E���el8������ͭ��c���60�~O���k�NZ/T���,$e�1�Z�����{k�j�غ�Sכ�Ʃ`fkǖnm��ȄżH��PU�[�@���ʁ��(�*�h(�Qm	�3]�����'��z��;6p��p��8�?��͓�:����!�(��%�VH����s���ڒ��f/���>���?A��9���^�0�5�� <P_6 Hy|�/>�H�T��ԧ
S����޻ �!��qi�u {�.���(oH���̨D�򚐍��X�gP�>�G}׹�X��gY-�7{%�:��y��]�ͫ �>��c��5m�c2\��Y�;�]���%��T�߶�u��R��]-�8�^%�;ya�ܨc��QZY�喝�ޮWg�p���vU�h�uؿ[��
~�}~}�������� 3AJ��B�zpJvk�~�������9�%�n<�ԣ�[yY��!W��UD�}��g������~�#�T��$����D~��$�&}RFDR�� y� 
�/H�����X
aM�l�W���/|���A1���w�J�LL�5��e��xr�`0!x�j�t����z`y�S������ �iYB�:�&���#��Pa兵mDC�n]����&������yj�й큱�Zi�}�ޅ�T)�R��WzӬW�\`�wұ��)��G~@SV=��vJ��L��ői��Ԟ��_+ȍ$�L����~`L�r��X���2��S��Zą� ��aѨ��}� �z�Pc.��h/���0�ݽ�˭}����(��O�b�/֮�ؕ7���٭�_���ZՎzŀ�#������y�]�����p�C S�h��9���4@�݆��hwOoE�y�OBhlX�s�E�t�S�lh������7# yӈ>q�m/%�<�)�� ��������d�s(,�y��9�9ٰp_���X��<�ԇ6�?���¬�~�z����
G��H�߷��/!s�:�s<��^��l�m��8�x.�5v�,h
�9Ȟc�B�WK�U#ߕ��O�w�ߗo��)T}����k���Ig������hp߃Z\���&�K�6�ޓ!�w����tk�5�'!�g��6m������wf[��8��\.�S�ե��B���]�r����E���%����<1��w$��Ov�s�߿�9G�"�$Rɕ	����I0�
RE*#*Aݦ3��2�� �T��Ƭ�
i�2.?w�\�T|kȃ�X]�k�:�!��d��fW�9�������~��P~��i���K �]K�	P�K�b�vmr�H��sӽ����V����'�-#�g�v~�3�L
��*7�j�$>��<O�)P�ʵ�^�ݺ�������m=����$D�N'�z ���1(�E�S��i^��܆��h����'����R�0�_Ϸբ�e���ŅZ߄oTI�����(�|�Jy�; ;�v�,5�\���7�/�^�K��\� A���#Ӵ X�(��p�+����������7�"5Na��xݚ��� ^����`��??W4��8=��˺�u*�s�M�C���ga5�Vߢ�׺W+H��]�S}�#��D�J��
I;L������0
�߷Xo������U#m�W����-�N�xN�C(}���dt��a��d�c��.{��Se��+�;��^_'Nn}a3Š�V
��<�	큼"����\l�΋�����uOx19��m��Xc�.7Lr9�H�#�Wb�H�M�3%�H;Z���o%0(�P����31gtǭ
�A�ڏ�ǜ�L�vjwq��	�Mr��U����v�ϗ�	/x�.ߣ+�5oq�̾ª�Ev��]n�z�.�69J�
�ک�;����� @��,�K�-�KR�Q��� .�;���|����*�0f��:�my��	]>�;x�NI���4��b�Hl�uPyeN.+1���x����q��{����`Q�3�vƘ`a�����b��z��"y5L�a�L<q�cg6�5
�^7�9}Q�S(��6��>���C�i&5��;⸋����f�)rD�l?�>���������Dw��ŀ�|�L�cL����=�hw~��e�2��Msྩ��'3dڇ���]�f� ?���g�@A���Fu��r$�6F@fG�b��<�X~� ��9W�?���y`z�����Ǡ
y��k�k�L�1ms|���+�ڒ*��{5��3K���e�Õ�(HQ�񱖌���>m�a�^�oAO��.x9��b��}����ZN&
#�¾��6U���"{�X� ��L����W�[����TA��%)����D�_l�(��E����ZIV�>��xk���h��~y}Y2T��$Jz}Ď�L��'dN����;i:��=�N|��SE���:j/�_Oy�➲����ko1�n�x�s껜B�x�?w��RJ�X�^�nD,k����ܥNV��a�J�!���	f��L��=2�*�NS�Y���]�.��z�|[u��]���\����3A��1���]oYt��ɽ����JY%*J^Y&%(R��1$���a
U!�x0p��#��8�Lz���@%ǧ͆�2��(r\D�Ƭ�a���� rW+K<��:ޠ����$�郡�WxxwL�2)����
zˀS�P��ŤY���&R�|%�{��PΛ��������v�_ �5��o�ԾPC�
���	��d�`-�c�Z��)��gH��S^���A�]��24�_]�h���Y6pω��ܳ>f�C�����s�u��D���Z��6T�~���D`ķ�3T[��c^pR+f�[j ����� 0���17꟢@x�������A��Ϋ��>,�5��3L&��s�7�O@֎5"Ԝ���1���OF�B�|cV�]�q?��� UE'�Vny�7yl;Ef��s��b_��>J�o�{Fн �R�-#Z� gK��Gk�:C�4� _-���W�D�Ⱦ�]�Ɨ�.���#�s��c<�^�;��vk6tU��a#���飣�����;��^����{��H�����Ǟ�l��%�j^!k񩨉[=w<�uý���`lc46�h�40�Qm�<���7es��4��f�x����3�>+ٰ׹�v��mo��ol.�T��.���v8�i�졤�FԮ�^��
7�W��R�:h%ɟ��CV�k35 ��Aݪ�"�O�#������sf�'h2,�������s��syF,��*yQ�
TR��E*|�p�{���|�Q�����k[K�`y/"��8��H�,�	�����<�t���GT�YYj����7�;Wԧ|�?O���r'����<:4FE����ev��d�����_;i��fdǽ�>�03�y�A��`�j��|��K4��k:2��E�{�����2s;�/-�7MG2OcC��T;:^�'ˉ,~�/�����w:K�9�;��>���ru�z|�ߪ��c�缙���Sz �we��n��B� ZD�R3��t����c*�s�]�n��8T������g�%~�R���G@0}�:��n,L���q�#�!�w[L��Dx�8��W��%��ܘ�R�t5ew�h��>�����^1��B0�Hm�ꆸ�.ǭh��_�ٲ��dwU�q��+ۍ{��8ސn1�C�q:�
�QV�<���"���������*c����/^�3(W�^<�]P��X���2�Q�;N��O�n�xgiF��M�v@c?��Z�xSqsk���5��m��[��=�xH��=�J��u�s����vs	�F���l=]�5�x�:s�|���q��s��Ҹ�2Wi��u�gmǰ86�2G:D^�ɴ(��v����%o4�%Y��&仄�{��ϒ���k3�F?���ے�Hn�񺷣�|�w0�ҥ���*�hl�q�s�K7-���wTݝ&]쩯:,���ܒ�a�՜�%i����;{�L�<:�����l�5ڷuҮiE��x�]���x.����	��L���⯆<��zu:q��y��=�3��+��h��ڦ��Rc�q:Ev�5h�xl��#�	��n^�I���绶�!\O�2��Ycp
����ݼV
�Y��[�%,��v�_S�EG�d�f;�dN��]Wn7�Z�L�M޷M�D�����\�h�gPU)ժ�@����X��V#�Q���=�+;S�!<�>�k:0��xլf��rY��}�g��E�4�l�K�����}��ڻo�t�u�L��	�S޽U�[	0��fK�*�U)c/�q׉A��IS�Q��p�%�j�Y���fJ˕�M�;�s���a�̕�ݺC�4`Z�8r<���k]�Mb铏9
�����R�q���ڭ��Y�eڜ�c54�`C��yg7gM��X��;�����g��L�p�ܸ�� ڎ�3Z5�k�c��+�~?U�W^��n���|���˧ϴ�5�[�+��"�w�`�^�X���
PZP�Z8Uȗ-��X�m��[�3r9�G�C>�N�4�j�Ou-W���ނ�}���UZP[�٫ND�nuZ�gi\/Z'BEp��r���w]aՐn��NRa�T��Fȝ�8�1���R�S�2�'��< Й�c�>ۄ��\�5b��*����B/w�(���Qe��n�Ӑ�r�:�c���}�c\�VL��÷UzzyOG&�>v���UC���Iʓ�5%�r5�D��K������y�Jﻎ��+����Eu�Ȝ'
�CfRt^�R�ʷ����Nڱ.��FŨ���{��L�}څi�7�4vV,V.�hNU���.���C7�P,�֬&�HH�1pX�1�]\nf;|Q�RK�
���:x���h�w��U�d��U3�iثgv�����c{W'��1����!�rŎՒ����$��s(�6��}d�̰;�U(b�8h��mnb�R��QJ���v�)ۇVvi��ŗS�:���x���:��O��I�N4Qξgl�[eJ�Tk��"Oo*U�^�T��wfVTu��#�1��S-�d|]^�d�e�9�*`�#�K:�Z{͙���]���r��,I��ޒI$�
, 8p�p�F2����d����?�h�߫�}�E�b"��߫x��W��)]_'����ӕ.>����e-r�ݩ�_{kơU�j�X�<:l������o�[��g��,-�(77����^,h�soǚW��O���>M�˪9_�'�Y������J�"*�{��CG�����:}8����j�T�ٵsnE��j1c-�ް�Jxt��ӧO���Rث%��-}��k'+�m���Zů�o[9�ĕ�)M<==:p���[�kx���Tj5�����e_roL�U)����N>8��$�`�DW���~Y5\�d�/�&T��SO�������~LF5������>��\6�E`ޛ��e�h#}�ƼvW�q���f�
7�{oO��o�r�#�b���3�WF"��ӆne�.������Sp�7��Ld�Ŝ��V+{���Z���9'A]�o�G������$��cXX����}~��>������Y����x_�-8
DFڮaP鴽5<�|zK](@q��ѷ��b��iQ~-�  ���H�����,���
�3����k�5�����Dsض���ػ�}d|c�,�h~�i, �9��u
m�suȾT*��%8���zC�]�����~* �e���}��:�[��p �~[�bG�'����[�����ce�꫞F\P�w�woIoM7�il��+ӌN
��)E2j�w�h*��H��2�8�z�}o��W�֫�E~��k�<.i�9k���]5О��y�/w`���HfE�C�z���K-��������F<�����,+>�����
��&wO�)Xi*Ej�_O[��k�<O�� FC���r��?P�1\�Ǽ �T]J�ߓ���ɴk ���U�v���պ��-}.�,����j��L��Xk����m����u�}�>VâV�*�X�c��^Gn$�;2��_{i���c��D~֑�bp�|h�����*���,ݍ� OKJn�؜�;{�j�������|����l�����yO�[��;q����0q��ݻӍ��OE���BR\�P�hg�<`��ٓ�'�.nr�w��]K��Ƶ��e>����'�VN.���c������]K)e6R�2�ɖ�2�{��ߞ� m�݆�N;aP#��,~:�6��J�	Y�},�Z�O{���T�KT�^6�p�9O�c�4�C�ؖ�_��oj���Q6�����}�b��l/�xL���@E��?���9ʾ�>,V1���9�X�T˟9�uͰ����>b���]�w�+Qw�D��G;��E��ll���+�D�ބ^��~aAuO1=�M�N5��yOS6UJ;��_ם�,�Ò�:�����}��|��L|X��=<] �ܧ��k��T �|����q^��yj�eb9�=nZ�=�4$' \O�$p�G� ׸_ӏ�粒,궗:��=Zw�=��p���]aD����ml��6ޱ��w�q���>Gk��cj�$Vs�s�i�����K���2c��ߤ��mϿM��Gl�:e����r?���!�>w��:�X���%�,�m�J?��P@����SW|ǲ�#Q)֐ ���rfy��I�̆�O��٤�~�tbz�?�{���4>A��8�����eW��B�4�ڶ��d�3�%C��,���0紭�*(�����&�ee(ȦM����ұ8J�M��k���ڕ���4d]gu�ׯ���6��Vȱgƾ��6��s �]�/��ג��c��_������,��.n�M���uu�+i����t����v����T�oF�0!`1�m��d��j��J�˙��{������.���<gW4�e7�1�޺W�A�`��l�?�u�Xο��c�?8>y�CA�A�P�c��t)��tg!�u�R�9���H�c{�?.pF����&M��`!�8�øƏeC�*�H�#�ġ�Ñ�e�VK�$f��
���<��\���ÔKLI��3by�c�ly�khWl����ָ��6��e�Mo�ؾzK��
���ӧ�f��#]�ǥ��V�J��Z�QiL?)~��T��m�U���4OL��bm�\;�-Q�l���n��:^�C$��Q���џ�*��"�1ڠ�a�=��@���d���Sm��(S�<Q��jyLت�{Ϫo��?Zq���Z<��b^���6kbX�cXd���?Lg7TY�����J��pƾ���=��G�����g��E������)� ���q9��xj�#�۹U1���!��l������T/xd�kI땀TZ��M�8�s>�0B�m�ql��y�G
y��4*�''���f����9(�.�99�4Mr�
 ��#&�c��� "誚�A�2!��*�n�!�{�&�sb��ڋ�h��	���K�l}�(mf�L�˲/;Sj�5�p��+�`3��[](g���4��^ۮ�.K���j�U��i�Gy����h����QI��e�����	P��� ��<{���a.�\ҽK;���ֶv���K��JD���se�ܺ?�����1܀��5��z�^3�_����nmB%����*�D��_@��1��]G75$d��(pG�%�a�#N��a� [tu��kw!��0���yh���E1l�� P;E��[�\�7����x@9�Rd��5����\�2�����v(P�Ɖ 0���[�Ƣ�-x�!C2
q�Vz���4w,⡜�cn����>�G�y�I�w�F���خ�˺]�H؝�5���J�5�>�С����9i��x��	�(5���(G�ǎ�%>��q/��֞]��n�!`�wmo2�=���W��OM{ ANK������K?=k˾u<~���ػRu��ƾ�S�&��0`_�h�"�!��B�eD������];������T2k{���̌w�伀��'�2=K��ey��A��|/ʾ4g���Ӱa��޸h����/ێ����}_�i	Ѭ_P��ނ���<_�@R����і�4����!�4�v�"���\F��Һ�l�Cpȫ�u���%�l��év� �C��H��Y/\�y������.��{hݡ��g"��-6+�j/N�Բ�>�;��J�v[��l�ٔ�l�m��.N��_l~�
��,R�2�L�dU���Υϙ����쥶/TSm�b@ڇ.�m�a�?�<^��\���K�&����zU�8���7n�}c�^����W#;���/geC`1����om`���!Ja�}A����_���xO���=:q�����3���	��b��vfP��0,�Vq �l_Wʊ>=ݙ��p�aA��V�����E�;�k�9�)�_yt�g���mʜ��p�o���l����w>�,?�!G���'��=��^��E�!�T�	��s*|�N�^��5(S2ힸO�rv����]T��1����C�Ldl|sW|(��H�PS�(����e`9؉7��Ɠ�v���� ϟ�gOKC	�����	"9��l`�r�sՁ��~��yw�x������o��K��N��G0[
�W����ǈ'+��>�ׂW?R��Ν��;جn���6(����;�e��q^��J�� %ɓ0m[��`$e�������=T�U^k�����ķ�6E��v�c���u�T�gZҨ� г!����˻%S-z�/=aes�b�RX��jR[�]b�]P<�K��M܉�n� gnu�]�'��L�����}��I��7��w#�҅Y���{[k�!|�6+��o�s��Վ�c�g�떇2�ic�%������مR���۩���5���e��}��">XD
����=w���	k4���@�)����.��ǢK��������>��8�=!�;�׾VM��*�F��?%�1�|�����ٚ�7�~>�U�AG��`ߥ��]��X�z��)����tPoQk#�܇l~\v_��ڌ1&Z��w���lgn���D�ފwi];	��G=Q��"�� �ɹ��L�0?{"ȝ�]��)YZ�~���l�`�D�O�~?!��[N}�]�x0��U�Y��94[6o,}��|�׏ɑ���Ncz}͞�f�>Q���N7�B����b)�t�3�~a~��v�~w�}߻.��?yޙ3�OV:h��dk�a9�e��xS.{;����a�lqV�ʬ�v�>�{���bw�z��,	ŋ��kC@��`Pv��W ��`z�y��Ak3����g{$�y��ݳmԔ�>x1B�°�Oǂ�������km�u�YQ�X�eRvלr�z�}��Ϙ���	���߼�d�QCߏ�,���(q>�G	�0��!���1�rp�(x�o���yJJ���s�ox�'4�k��>3�\,��U-�X⳻��uK���>o^~/Ѓ�����VM����k�R�u����4^�\�;5�Q��Y��Ba�}�t�vb�p]�Ҳ׬0��" @��"	f�W�}�����KK�߽�sw��"��� @#��3�ioW����=�"�)��������׿8��l��jw���C��r�o3��U�����z�5t5l�5�-4�Mo[�]thߵ羥�1�4�w5�>�o�X������s;}��
�y >��Ŗt���G6U�1����JP'Z�M�%ͯqq�G9�����_lkv��Xe2��.[�Ǯy�1��9=����@1k��*�,Z<oO���̳P����ܜg_�}�`��U�@3�?lX��]�,�I ă�׼Y���oޯnH��M�y�Q�7≼�a���ߌ#���x3\���z�2j�κ�ŵ�ݫdXa��������>��\�SYUĚ0��B�o���|�r���!0�K������2�	���o4E�;�`RMӧ,ͫC��x�q�D�dT�$�[���!~(�Y|~�T���:#�zX0�3��fNA(M6�v@ND����cB���&�Ի�^�z�:��Z��y��s{����b�2�Y2+&[����Ku�f8�T'�Y�ȅ]`y)�v�)\��jZ���R�G�&�Я8n����d{�!����|��ͽ���cF�3��_n�'�vܛ�t����Y��N�w#�XG��{����w9��}���<<�@`�m��b�E�����^��9p@�W���m�·�/�閽�ϑ�,�ŇK�T��}���^����|l�a������f���%��J��=W���([��3���ڞE����a(�K:P���
�sr����D��
C��~��Յ�>Q�ex�ve���;�_Hi���u��%:��ѻ>�Z�\��R40�L!�t�x���!�4�!�������i�0ɪ/����y����u#�[z�~��,���=��)l������L��s<	�ާbd��Խ����]�zZ�}.���榠	2Yv/J �k�9k~�0���O����4h���9�@/��߇���`J�cF��9�����������Y��'5���w�R���-8K�O��8�/���Kqg�c��/�_~�|놻�7#�����5S��U(���۲,�+�`/�OWr��?yt��8@'SЇwΑ0���^U{WOU�>���,�"���ob�E�^J�����<�D�z��� � �_���g��X�޾���AF�`��O~�{S���k�*Q[C:���� N���-W=�"��嚍�ʓ����O����DK�m}���]�Շ�FwnL��`#%���WH��J��hΥe��)B��u��oJ�ͫQ_| `�`��7W������ #���a�[g2}[`b�	��H���?//奥�3�h���5���x_[GQv�n��DGF0�ܞ��~������ˉ,n�����X7��Ht*���~��ҩ�����S�@b���:>a�ߓ7hQ�@Y/���;��>����y��;��	y�G�Q��[;T�o~v��kW�����g�6@g%<1��za�fM�V@��h2s{N�����?� �/شJg�%�+/~�#�Z߱��?��Vn~V�\���xs���.���Һ��<�x�	i���{��s����T��s9�im�QO �+��W���i�Tz�������u9f�1l��c������=^�]{@�����z`s���s�D�
d�B�p�2Z�Rކm���E�t-z�oT�{�Jm���t`=�\��׋Ý^U�}��^_���y���^8`m������o�S�>"�A`X0f��2�f>,aN�P��6s��";�}};���B��P	b&?bA6k�<���# �8W�Y$'���j-�N�{���U4EZNQ�USWa1�p�x��*��ސ���[[WI�3�"��dh?)����E�����u��a�r�7�y��:(s�S�X�&��M���j��>������[���;��p�).Qϝ��ǩ�ˌ���RXNt[kT��L���`��GD'���T{z�u�0.�Xʵ�]��<rt���\�;��k�0���:�|���L�vp���K Q֥V��4�77��ZK+	��-����ym�S��ܨe�Ցi�N�kHJ)�Rv�^��*�ƅ�ͽ/���_����?��-7��x����qw�`��PoMgOJ�`�%b�E^���"r귷��Ep�Mj�h���,_������2 ?[�Νm���3�/#6f��<������iE#��<w�1�ٖw�M��Z(%���o��7���,'�.�.�o��m[��S=	�ȭ�Zw�)�׍`'��,�=���sKQ(إ�o���Wj�<�g���"�h��K�'���Wn�}gk���5	#T۸y�WH�64s�� +�F;|@�׻|�}c�UA��ͽ�M��S���:)�#����Z��ӂ�����%f%g𲾗�t��;$v�eы���`�2)�����>M����P��&�%���hR�������=���͑+�>��EŻ
e;�
�:26�Y}+�K+%me*86��x]Є��V�̪A�s�_��Giƪ+M�A�#9�yF�s��?V��z�;���7�M#2�h{T��/:Kj)RkY��n�7�3����Z2@��'ct�"o�i�r�P�kkn��&���T���7�pD���IFd��4���cl:8�$`�cHܺ�x��mA����G a�vP�󐻾ݤQd�ZM��;6�u��5ޞrr��ɕ��G �~�]���T'2����q��,X�ǐ���F�\�b�k���]b+V��ƳL��kNc��̻F�{q�$o���➢�7-cx�m\vu�k4�_-Xs��FuX^�Z�1.�ʉ'ӦG�ι[�.��k��`�*����C�':��f^Mc1SY�n�l�t��P�q�x�r^�z�z�Q�dN̈́kWL�Zq���F��TC���n�]kK.��T��Y/&���VK�n�ˇ��{H�6�ea��y��r���]l�M"�K<P��b�c���/jC�x���36v�jz�U�7fj��ڌ�g��f���:q���he����uê�^�p��\�MUxk�:�6��A��ಮ%Y�[y��:62��#
|%ΊSs�H�0r��-Y�z�+&�i*$�f��_�B�5�R��5y���}ԛ��Z����C���7�����~k�F�
��[���j�2l��`�A"R�g�N(XI��!`�U��P]�j�ͷ �:=�HE:l�ڰ���'��	z���00��K�,��A����N֟`��+�������X"�s*o����V�T���$S�U̔�T��}O&�j�9l�7K{�>��lY��^��3���ԻH�d���M����rE����qn<���C�=.5m�+W�]t��\�Q9Ӓu�t���bU�Un�v��b̝�.���˾Sm�]+1���a_�)�ypp���(��)��!0�qg9J��sm���ov�����݊��j���g�@���o��d%�����˪��`ͮ�펛W���QԤ�&�{���z�Wm�YH��݌GeK�L��YA�T�����g'F�ŵ\��|�'0�c��K^oT8o�n:�L[��<C�,�2u�bu5���o^n���yA�*�A�֮�ŷ�n�U\u$Q���%e�\�ʨ8��4�{O.2[�)j<�.��pp���=۝�e�v(D�1u���+���X�,��lɔ����lH]0y��XK]�4�`Y���u��T袄�&b�Y��z����%���F�7)�T�JӇ$U�.c�������a�ڻ)���,�پ%��J�����6ﻻ����ӻ�t�I$�4��
l�m4�m��4�T���i������6x�[ccea�+Ll�c�lۏx�cN=V4��JǍƕ��Q`�
�T�@�E�d%�.*�7`��LRR&�h�$b�D�2��R����ғje3�h������b>�x׌lF��X��{x�P%��Y��SO������}��&K-�wZ=9��~�q#�����1Q^�קB�P�u~W���M}�'�����ҝ�,�o�>�1�~y�8�.{��ɖ�-���)��Ӈ�N�+�>-Ȉ��%�~<���_���H��.y݋ W��-���0�G��Ӈ�r�f��׈����_�^/��5�/LB[��B%�{���L)�g������N[e��v�W�$LYJI�,(����}��i|��l���N��UH(�|We�6��Qs�"��ƕ�2�2�:t��ӧ9{�_��m�֬�S�@Q���࿻�'�ܣE)^��W�W�W�Ĥj`_�.^����q�߽я��h���܈���k�X���#��Ro;��Rh��1��]}��y�����^�\�Ih�����1��;ȃ���5�j䊻k�N�����^�h�ש�:�uk
yR��8q\���}�SLl�+Ji�J�٦�[g�(�0�YH������ �@
 HW�ߓPe|�� �����D�G�����@>9W�� \�\C�>d~3,��tSdѩO��ᵵ��A/�ȏ~������W�Bv�J�~,��+�uоt\���������
�z<�-kqX՗�ל�[m���T���w`���к<�8��@M�d=�l�f#���5��Q���p/��?Es�崅����z�=�WP/��l�Y�[���q�9��gjʮv]�Kz}vOX�s�r� �n��6׾T`��e*_.,����J���K��[c_OM��"M��l
~���+��[]wAc� OJ�ش��l����%]�g�*�<42|�υ�?1��y嵟K^tse[�<�|�6�m�)`w�ȗU];[��4p�`�n�y��(��=�lOm<���0�]�_��.�^��Gըϴ��-KQҞP���:���s���6��
6�H����3����?;�gPΑ�d.R��!�:16v�����Sݲ����E�`�ѿM�J�g\�.���b`vV�fj���}��,Ȗ�jK�U�L�ݗd�P,<r��/]'[����~�:}� >�� G����P t"M��οngkT�UD���,�8�:P(2�DW�#/$f�]$���Y����W}�� �0��y�{�+��M˲��3#�ݠ�cg��8����9E'����;�3;=�����Dz�G���9O���Z��~�.��A�l�<���2�f`D�t@wg3D�a�k�O�]/�5��©|��0=y����R� ~�����*;�h�',�Y��S0��=qՑ@2}k
���M�)RW��VZ�AT�
6��*�P;��ox�2i�[�)�p\�~�g�:�W���7X21���n��X�]�+ l�·���;r&+�T��%)���zO��E��M��պ����v�wn!��Z����r�5�횆g�t�s$H!�f�p�nv@7uD�0c��.�d��VWM��>�r^���K=��]6,/#3x�̈�W��0�3l�f��1��5���	�W>�I�`Mx�A�r-��9��,���7��q��3��8~5}s�F_}k���]
kew-�<��aNoY��_2�~������!����k� �G24��P�/�KH�^�u	�9�#'��vS�&�<�)�y���VS�5´�)�bv�E�R5���#꼧_�	�2ʖ-hRfcI�ƭ�0j`����M»9Pႏ����L�Q����r��a�#-�sM���L�s%V�I�oWq�沫N�
�vw��]�k/jkb�k&r�{��� � 	 3 �[�����*;�L������6f����/b^y��0zeX��Ǩ^��a��9<30�7p�wkfA�cO �>�=)����ͻ���A�G��:j4ހz#yՍё�ǈ�bzk���x@����&E�����!O���%�k���A��H����1g�d������٫q�zBy}@\{�p�֟>�P�@3Jo=#�����k��D�`�͡Zc�]Z�"8�
u�^��c�a�|!�2=H~p�õ�Ώbzk`��ԇ�|�`^p��%�ʺ�ݙT.��%��0��`r}0���g��e����<����7���U5����ئ!�~;��4���iey��w�����@���̴(��F��a0�𬿎%=�Ƹ}��1�nPj������r�[� �Fט�Y�Ĳy�~���؍���:v�j뭮�����lsu��e����9���w�4��
�p?�<���%��cc��n/�X҄z8��rpbv$SSs+y���:����qO]23�Lv;���w��+��Vr2�y{q��-��r�{/#o��ƴ�%)�L]*��렮J�g�3���
Z8T$��ػWu1�i�����aoC��V�ѽ�����'Rx��xժ����n��r�gFr9)h��?�\ ����>8�3 ��x�D�\8����HO��&-��[�d���1|�k�ܕ�]�e��4�=re��!uxEp��)(g�B������l�����A��f\�v`��`E7'+���r��`�&��x���Aܪ�{�cq������N������@�_?�ּt��TV�OB�@�8ȋ�<N���k������c��3��;�9�x�<�5�t��u������c���L�"��z�u�.2Yu:I`w����]�k4x��A����9��ǁ
�������.��)�Kz�8���!��%�:a���f�%Ɗg,����6a��rֶ��ћ����4�Ŋzn}���p98�����<Ui�'��ڼ��if�Ħ.���u(��n��Hy�v�a>��h��D��%Tӊ��k?<���kWt��w�HO8O0���ͅ����9��N�h��(�� ���_�	"��7˽>绲��~��o��l�HR��V�M���@.��g��1��X�b�~�iW�7��,��~������Zخ���!��p�t2����J��N������vclqm��]�°lwX+�3��`-���%Y�-�]:N�εws;�Ɲ����&����Ǒ�R�#�H*���w�.)G�L[�i*  ��!�����?�@K?π�H@I � "�K��������$��j��./�x���d;���C�Z������ z��рe, {7�.H�]��{ e�2C����.Cv�/Ɔ`�$���"����W��E]��疧�c]i呴��/�\� >�t�&�@x�s*)e��û#=M��g; #���~�B�kMT���]�;=�υ[��f���?q6�PW�/"�%��X���t){��X����P���l��k�,�����	
,PMr��>9�C��W�g�{2��|�¤�����Uj�>�5�Ke�����1�/Z�Z��@w�~��ÆZ�X��9��D�>q��1_!]X�ü�Im���M�-M�%�/�8��g����aȁ��4�r�Le���Br�Fq�����)8��S�y��к������ ���4z�b�46�{�H��3��}ٞуB�B	�|b�@/�l���`	X����F��Q#u����mw"6�*���ȁ!�A~}�u�XB��;�6������+�K89tw=�~�a��H2O?�|Z����U�>WL%X��ɐ~���UxȺZCb����g=~���}F�.�b���}��U7�q[��v�1�n�I��Ə;��۔4pB�ud:!�%��[������{2�#R�U������� H���\��b�~��Ph��H�rz������ώik�k�Ǘ�O�Tbڗ��}���y���~�<Ʊ���
��ʢ�U��R�����+�f����l2UD�qF��SQ��OW��b�C�� `d??�����ļ�Ç�m���T#��	�N���Ǟ���T�=�6�) �������ɦ�"���z��^�F^�3�>�u�2�2��]�2C8Mz��r�.)�K��v*}�,곘Y�~��ۛΛ:��
�L�a����ŋ���A�/���3�"0���5���o`�0f=��c�t�_����x��A����&��.���QL6F)�a�g�2���&%����w<8����^s�1�����nW;I���=�B�	j�LO"�{�����!�G7H��h\4eNvi���&-�p&[8����m;n/ W|�P���m����
�4���^�����&�M�3���N�����1���n���np�=ј��g�F��Gg����>B��"�B����~5�[^�k�=|2��(wfe���Z/E\�R}V��׳{tj���y���WQ��s��ts�,6�.���;���\�h���\���B�VbΩ\�9j�C�]Z�jJ�)f���ީTX]���X��W��{߀��f ��y}�y_<��|a������ats%~Ρ{B����Ɍz�M�>��������%��d�'_�߽�P�r*9��j+�Z�5����y�4wP-5�(m��E���*Y�cU���G���eQ��S�'�v`?�<&~7u�4� �OB���rY�ˡt�:�i�3����yf�r-1ý)�!�f��xE�_������э/^Q�͵r;���[�&���չ������ �M�G���P ��|5�A%d~y�*O/���{�+�7q����3��AEr`�c��g�^*KJ��zN�hf����Y�p��!�?���y5�S[��I�u�Gd�:9@0�
mrB��Z��d���ZٸkK�N�n��x"�y�{goo/��� ��zE�����%P֟>��@k�t%�5ܩL%ԉ�~���ͪ�����>E[�.d`�KʘE|�����M��X�g����z���Lb�����G�:c
s�_��V����1�����(8����`_���i�`�}�h`ʭ۬o5w��`c1�m�yM�Ǫ�<(��uO��#b������P�O_eȞ�D1ە��X�+�2��{h�F��6)�T�e��x�������Ȗ�*U`Kx��]�=j]o8r�u7�S�U�ǲ�w���؁�����3 �0� �gq&�n'u��|7n���𴻗�z�������*��j����ێ�+�Y�ca���s7�ev3�w=� Ï��1�=�i:5�����������T%�>TֺȞ�����/1_�g݁��A��?�i����竡2�UЬ�������ҝM��+~_�k9�$��_}�y�j��n��jd��=z�E'V��nzs]�mC	��m�9��ήTv:��}������'xI���1�I��yqC:��о̡���yb%3U��qo�/�s󸦷`W�zq��e���f4wB``6�sזE7'w�P��{;���d�w��fn`����_]y�#)Yq|p������>=x�{�0:~a}o���'�o{��2MI�=+�c��ǧ�O~�+���3Uj��9D��`&�~hO�/v6p~3��i�y��S�5�`I�˸8M�,(
#z��Z$�K*ϧ��^>/�~�n{�]�VcAI(i�����ugu��0S��\���c��"}����d��`0XVo���U}�Jc��8�:RF7�c�-̒����tZ�9#� n���r�yc�`���xW�5���v��4��@�`d���)��S�ʓU7�j���ߋ�ྰ0��l�t;o/�p��4f�;�fQ�9.��w��TRꃴ��^�vtȷ��M#t71ӕS�p���O\m8�o�cM��˭7�1��O[b�� >@~Dd
M���-S�o� A$�Q�Y���5� j��N?� g.��jȡBԆ�P-(ÁN���~W��)qBf��]'�M�d<���`?�����)��orެkzi�nh��w�v�<���c��D�a�3hq�:��~%|��`7 ��,�"?+"������K�e���q��kቿ{(�wwpY��~^��9�/�Ħ�[��k��>�n�3Ӊ�MczW=�vצ��e̫���^]�ҵ���k�"���̵��}��,�s����j�\*��3�C�\	}pP����h�c�a�6�v8۸���ȺzD
:���ϒ�S��wlX%���~T3���OzFn�*�[�!&E��n��}� >�	�t+��i�3�U�^}񐯏i��ߚ�����0-i�������}0e~��y�n݋�bd:P�c{pNtw�3%�u�Z��݃��V���?	���mO֏�}��Q*6`k~W_�c�ƱҸ�Ȅ�%�qw�f�yrr�n��n:hk�T�;ʮ1VT�E |�x���jC�~탥���W����V����n#6���R�c�����3,�����}[7��w%,e"�-�۝"A#��Y:౔�,6����ޡ�+S�:��CY։N�D���+R_,ä���_Aܨ&/����s��kL���E��jpÀ��,0�Y�c�gLqO�}�\�qj�2Z:p}��Ƒ��E~B�B�����pc3�2t����lw+~M����(������>����J��%öy����l�C�L�+�G]qt�M�=����Ғ޳�`m=:��F��
$n�o=1m	˻��ҝ�پf��<�8bg��PO����fb��&6�1�:�n9tWt=��0+%��,iC4���j�C%"x�?=cAb���k ?�[U@J��<�t�>�0<�F�s��x{��쒶�QOͪz���&3Oy�xfδ�K\���X��?�z��� T|sʱW�=c�d:��Ңoc,��A"�N{c� �L�}C��#z�<k��L|�]N��g�B�<��v4g�M:�Z��~�I���!�-���n��HM�#j=<b�Q�7�L�g��Ruu�
���hD��9�x��H	�>�f�#2��#('o@M0���wM��RTs���Z���v�\`�a�v��t5�{׆�]"}�_�}%�Y�%H��A�wa\�]�k�w��x{����
j�d���<��Ju9�2�i��δFBS�Қ'�e�wN�j�ŘЮX�J%�0Y<��k��_�Z�^9tf��h]�8240��5)�/.+kU�t1g��Uk�.�Fek��#�]�yU�I��:�#�k�K����9wq]�ɐ�B���=R*���r.�aC bqf���RRpݔ����﫺�\FoI��k:I��h����kɗ�8���Ӓ��3�1��J�;�.K;O_p�\C��nB��
ޠ�R�U�E��Jêw.�>MZ(�]4�tI�:�rÎ�=�I���!4�t���{Ի�А�;K��:�Ev�5}C8�O!�J1�A�qh���Q݃p��A%�z�-ʘ	��ڴ��NhҌK�[L�<�5}\wl�\e��oF,bq�Ҍd��5�*uڤ��K��f���Zf�ִs�,,��kx���(��}�%�OJi]�֊����[��ܙ��fI���cީϏ1g-�U��L�+-İ̷�����}ܬ�m�H�a��UTM�Fŝ�s+�,���i��:����&�37�묑�T���+Y�F�-����F���������ݴ�cyN�8��E����p;˻����/%$��~��Ny��^.�f1��~dx_1�i��g�L%f0�3hA+� ��@Ġ`"���
:#_ ��]�+�64`�J�"��(88.���� Q'��)�7���u�E�^��b0+X�F��p�;V��dBy�|�;��uΛ���s�ژ:���sKmTq����^Ǿ��R�����n��yfe�3�����F����~܋�]�C1��;SbeM�s\F$���zA
�<�Vm:p�tˉȦ���������Q��&��G�Ț���U��Hl�Afu�ǹS�S~���.�ś�S����Ru'�YTi�5�fou�Z�ECpW5qZ����h�V��lYKQ�����7�SuN��ն(q~İU���E�N�&
�Y˔WD�V�R�;�3�8D��F�&���]M��ηC����R��e�i:;��v.ڹ8��鶛�(I�.��.�O⩾�����ܓݜ�Uƈ�	_^�V��W!����uX�A�8�m��5䨅j6�3s%D6𹆪�t����w�c��y0��/Wk��k4�4%	f�Gv>����܋��z���.��m�Z�8�ըH�<�ɽ�u�E����2�c��uZ�.��/m�Ij������b��i+���;"b���rE�;�|������ͦ����w.���h�1�A� E cD0s�~Td�~6C F��^9����F�$)@�y݉F�����©W+-)��������`�B}\��^��dfX����!�������,�U��Jzt��ӇO�ydu)#3������I���H�e��)1�iXxzt����-�j��]�f2�񿥼(��L�W��y�ٛ<��?�y^��W�W�~���$ �� �I{W#��J��$I(Kb�:t�ӧܫ�e���j}�d��}�����0���ܶ�e�ۑM���:t�|�$0�6�u�}y��wl5��<����:��+�FfE)����~�~wZ�Rh<k���wnR��O:�H�#Wu�i^W��t�ӧJ[.\���ȵ-[�f	}y�/�]���g���;s*��~.��;�z)�s&�]�<��D�=���oPt,b�+۾�]ń��r�v��۽Qލ��m�����k[�����-=�2��%.�_��_������g�G�|�gPM�Z�,b��C�"��PS������h	p}�d�<�V���_<�PA�Fx���'z-�$�;�=C�@^�
@P7���A\�ʋC�3��7�?<���ܸ����q�\��ܼ���{�U"]̸�qͼ�sj�$��U�}�����[� ~ ~��Y�_���}��@��cp���1��p�3��΍���n�;�V���ٗ���E ���c8\8~�4��y�8���E�?1�����cp{ke�_ν.tCtf���2��>�'f˨,�[!�$�V���HOP: ��u��ֲ����FnR�!��I�q?C0�ǫ9�@��CkO��sM.�*�Pv�rY��c��3���3�o������	�1�"|�2�vތa�'`ܞ���P�� _���j�;9��h�i�w�h���͌�Sp�xy|���������$X	6D|��e7���|�MC���44񞫋��G���O��2���uy�
������	;��9��l��}������[�Q���7}n��8��5��uf�_8f>���/�I"ޑ3R���Ib�%��yN��q����w�ӕ1�ޭ��W��۹W���6����鴤h�o+��[�ת�7A��O9k�\���:'Y����� H����a�p�09Y}0���ё����������8��Ɔ5Z2��[�;��2f���ui�칾��/�tT�*!�� �9�T2 ܨa��/�(k)&5�����k����_i	�.s��o�Xy�&
_��_��R�����'OmG�T!��s������9��Q{ܰ�}d�eR�ҿ|���}�O�v{��ޙl���s	l��J����vh��P���n�r�wE�ؠ�yאԉ2;�mĵ�w��7�=m��L��o�XR	���x�s������-!�w�N���ETE����C'qǶ��b%^�kԀ�mE���u/B�sm���'�"���.�9]��=�MI�����F��O���*p�Z��du���0S�z��N�P����uNð����6�]d�V_
P��۷�E��eA�oG3S�&�\l�NDw>X=>\��V:��O3/�Aj�bN��;ֲdeD[㸦�#$N�:��ۂ�y�Q���k�|��iX�i�G�����]�/�U	�~�{+Y%K]/��ae��=�7�Ӗe�X�.�l+jY�!T��_G_��
�P�\+�TY�8�u.79!�����u���ơ̫�D�b<��t�4k�n�/p�#}1%ݫ}�}�z�_1\V4�i�V�L(�J��w*����  @) H/��Ui'��/�}���@�@�0�iivcō9�w*񲮁"acx��	��v�[�؆�|O���5�ε�m�]�4���nM���-�^��t���K��p����Kxυ��p@T�����]����`f�b�	f���՛YΟ	�Z��p5Ӭ)#%��2�8�zm89~S���_��q?*��R�}c�-�㎈����z|t
�V,�.pE�w?s���B8���O��x�3�g7�;�~ϝ�����a�/?�P��ɖ~X��s��3�ǡ���˥@���w���q��I�h�jm/���x{K@-oP��>?������_+:���W�^5|���WW��]s�=?P#	
�`1ϔ��?�����9h����.�bUэ��+C���ҏdV6��j�]0�l�4����hzO��=����S��c�{��C_�ѝQORe������@�RjW��}�U;�\^�c�縷}ο���Z�L���o<�������u�����#	O���}V�<h����7��Ao�$��H�/j"�9�#��m��>�^�mVnk�5�3��k�P]+=F��>9`���[8([�r�i^(dN\ۻ��d�i=Z��Ѹ(]��
�3P�ķ�#z�Yr��I��j���̺���,cv��]s3�����%���7"s(@Y����>8�`� �q�%���{����p��2u�\&��E7*���4� 0�P`&Y�WB��j��5�Ԭ�&�"Y�7�F����ON��8CP��o�t�B�� �-�����@$����,�d������n檣#�U���7(���?s��;�R��T�,џ�o�X��F��L#����h��X����j\9U2糽6�}sl%tY�/!���6���"6��:m띩�P�W��ݬ��P��矘�]s%���m�3�;~xq��4���v_������C��9�w<����$?(���)�<��h]�����O@v�`m�v�׆dZ����.i(��X��38�;�����>}oz�t�R!�N��5�H�~�,��w��#��oc�h_�� ����|z��9/�!���-l9tw>�ڂ�,��K�D�p� �̣`hhvC�)�2^K�W�嵦0�5gG6U��z��˒��7�|�0#����o6H��������w=,�E�s�y��L�=�4;���vK�� �gl��3��;]C�j�30���PU;9#��40JǬ�����b�\��:V׷��b�ԍ}�SL��w9w+s�gb�Α�j�^ʭ6�QVsn�.�%�J�""]����}��Z���v�����?t��2�Pw�{3ǹ�ۆ��q��5�-��ɪ��3�'MpG	o������g��T�9�Mq����Ȯ� 7�^���}�FìY�Iw���yy��&
#F��儳�fp3�������΁�#�����a�\tK��[�``���	�h� � ܺ}�v<���h�\�o�$�D���d��v{ד�����dN� �L;[>a����%�j^��(������r�������S=��L���̔y0���{죒�s~��Ϩ���Z�ݑ��˜�+򦬵��Q_�����[�X�|E���
Ws��Ɔ-����}�G�>�(U�[L�P��IQ��b�]�����B�<�(�S�τ?�X�k�<~e�|���Κ����1�t\8�y�i��c�������_c[=l
d����1��T��9�ΑY��=�b�pw�6*�G��&u�<>N����>�|�L oyO���.��i�����[�\�����lwP,���hx<�LO
�h�t��3O!V��������
5ϭ|���'$����̼������@��<��:`ǹ���SY�R'Ӧk�0�B��s�z�jgb�8����M�k���/���wǹ#lEZy��~� o��U�H �	 ���C�~�����Co�=G<ь"TkL9#��4�<CV*�>َ�6���mrz�E�U����p� ~7��@=�"9$p�8���'�L�Jܑ%�_@����'�7��Ga�a�=8��̕����F1b�E�y[<��׉��%d?�{ʀ�y}�>ߋ�����~�d�<��rp���c��b���?_y������B'ma#T ����ڧj���o�(�1�S�TX�|��]s���=m[��Un �=2o
�p����}�U\����7o�໘�0@��[V�{��-�&.��f̰4 ϊ��P��F�t��������'�-�@��|�����`�{-�g��}�^`̧o��?&��vUtV��n�Dz�>÷���*�g:I�l�}c0g�DU�=���y	���]���墘ש����E��|fl,����=�%���55����� Yǭ�*uq��;�y����kmgnގ��5�3��!)�prb!տ�sH���֫��jR��Thy���sw�W/ҷqЭ�S�N���~�V��_�}���0���&�>�|R3:=B�g�#۲MT�7Z��n�˾i�1��竇1�Y��=�B��k?�;.ƬH&�k���{l�SR���h�݃#�<�G��o��^|����W�ڱ�<+LP B�ɨj��-��?� yQ��S3ן/_o��w��쬇Y�v�]Kȧ�/�oC�(y�Q�Ьߥ���S�SZ�m�������]q�9������jN��1�ZD�z�2�/b��W#5t�7��娕A��1Y֧h�B���vDlc{�A�!�D�L�1��9#�{����lփ�OON%Қy쒶�6c��^T���5U�u�C	t�����=�"����	��i��(UM_u�&{i�^[K�o.�l�+���̘��zoE��@��li�C-z�`͕�_�Bxl�3$#�e��?�,'f9�4��槛�)G����0�|��:�Iq1�뾡7���);�u�;V�4c�dH�8�,M"��}\}���?�󣇏$��lOe�r����j��۽^�>�m�>M�"5%"N���!s�?�.,���{Z�[s
{,�%�f��L��xI�+1�M��3Zi���~�����j�r��u��3��2Kzs����0�*�N%�F��ͼ���N���ފ��� ϧ��,ށ_c��=y(�`z�ŏ�Ag�J��_k���%�i���ɳG������#bVMoi�c���཭T^Z���w�Y��Em��kT��P��|F$e$�=�g(��M4�rOiz�_s���s-N���>�J���ʙ���\�ғ��]����	 �	 ��v���G	\�}r>�R��C�$=�u��Q�kT������b�n����}��38R(�Iv��ݗ#�ah�O���o@�7k����;�!�P&x4_M�i�"1��opl���2q��F�&�l�h�i�3�B�/u}����nUB�ԇ4V��M�^P� �k_y�
����@~�S�4�{�#��8��,�C��m�����q�b�R�nr�m\v�k�^[h�m�w�i����YVc�����<���n?�vΙy�>�a	jFV3���8�Όoh5tz^�<�W :۞�]]����-Mu�Y	-���q�4�q��)�5˯ ��\?�?]a�5>u�U��T�,ky`�[Ɣ_�ơ9!V�aqk�wW~�`++�	��^5���s��x���r�@���7���P7��n�og��&WvmGqO�i��W|5/�Ъ�b��-V..=rޒ�����є�ލ�R6�5y�	*��X����U�fU�[�6����+��|30s�N��[�:�Z�1��;�,�Ε�r��2�z
�kl�Jɼ	l�[�]E��et��ۉ>8E~�@$��h ��S�c�����o�K�?�'�
��y<c�����fmiI�j���Ԣ�H
z7� �e���\y]DN�}i��ݛ �齩����ڏw{�?�S�N��A����P[���4��~侫����������p2�+ͷ�8�j$��#*��G-�� �0�Ӏ8\��c���mRC�����\,y�;7����>���s�bv˘��@�|��vq�	�����,,K�vfEnƀ�H(�v�`Ϋ��s�R�A�=�]L`�s7���{��U@�f(���ML���ݸ2T�ScU��4v4<�U�<�ٝd5��KE�S��<�U�t�,��$m_8���}�橼SG$�u�7a�1Sbg�jU1g��7R�o{cܳf�m�V�:�e7���p)b�-�3�kR����
���������<Ĳ���:���j�v�)��٪圖o+D��ĕRR6a"�tZ|���=��NN��uW�t��Q
�bŌ@|#A�N�e�����|�T�����h�ǻR�;�N�yAÃ�u.�M��rgh�1w9@��!�3 ��`�=v�uq���`Q�3ʃp\�<��}q�M�����.��P������F75c�Z�5�����ZW]�ygN�wb�[E[g3�}����0�>�`�"�;�`���Mt�T�h�,���K+ˏ%y9������L���5�i�/��U�����/�+B��A`��w�v�Ļ�v�06��W�;}HR�pl3��2e���0���Z(���x;�sy��o^��'h�9����L?��s�g�v��k���lGo�`�۾(�,Z�O����Ӧ:���8O}!-���=ᝯ筋l�{����������hG-������9Gc������V4@zzT�Uw�u�������}W�J�����'uvH:AÒYH�����~�u;+vþ��%���=? R8r`h����@�V�,x{�8n��8�+�(c���%K�Bn\�w��)A�yC:#*R�MM�6�K��p�=�K�l���=��X��I4u��^Q�%��iɡ]*ٹF�]ic�)61����1xH�:�y�0<z���ۀ���n~��ߏ/��v�`�>�Pg]қ��
��WZ�-�F�E��{j�1��|0�n#S�v����P�޾�v�
���A���g[m[-�����u1�Yo]&�m�.��.�����v<�&�X��kͣ�]Թ�Vs
Osm�E�,�p��j��K:�Lp��z�U�M�d��t/��L�@�,�W�YcN3Q���+���&476Rx2�rs��	w���;��kgP}��:��n*B�xh�x�VѤ���b�.����V{��œ���B���)̼�/����@��[��P��,y2,w�j
�W^�xen�u7��f�ue�b�@ݗ���m�Xx٫r�>�ڻ]�E:��.�34�EYhQyr�8���B�_2Q7�Ս�	���t�r��r5q�F��ô������ʪ��`�{gdDL���ȟ:�s�4�������Uբ�妹�.mZAw;.�խ�t����\�w�E񂶩�TxfȂ��Vq�-k�d����N1m3�lp��Hp�a��[�`� d:hp{a0z�Y�mg�i��h�i��K�4��$ ��\V#t��R���Xo��(,N�(
(�g?!B�Tz�0-�ob	�:���N�xv�cJ/< �C�����Y$Bh�O<'�B*�v �x!�:>X�;O�u�0���:�M���6Yw9[Nv!�WW.X��6Jc^�O��8n4�
�qI���+g7Gi]�gHgqf��{���yy�5�3�y��v��i[��:��k�+�к�yW��r#;rx�)�\1�7o8"A)�R;�=SD�r�K1�[&���sh�7�a�1��c��6�e+*�s���W��.��P�<`�v:��|��B-ّ�O6 ���!۲_t�[��ʁ�طE��άt�6�$�Vv�=e�:%����F�P��:�LAa��u�i���bb5Е��fVi�E�y.��;�ƾT�
t���:�P��̳�^�Q^�o#"��N�R��%��n�����v�6�Ahi)y����^�X)涫���%�u�a#�s+;��:MG�#�bV3A��EN��Tf��̝��0�Z��dm�Ǯ���q�_q{RK擡w��ԸN�Z�}�΍N�1*��̂�	9n�&pj����$^�N��p<��l\���lI����O�./e��X��hHT6ʩ8�k=�ĭ�]��+���T�6;r���7�r�wt�ܒs��:I$��uXƊ�^��lxяҦ��4ƛcM+m�4�1�)�G[l�iⱌiLi�b�ciXUiU��ٲ�j��b�m�hHTlC@��aL3Q���i3h&�i3
P�#l�
aER�_�����/�"�$��u��w���6r��xwk��w;9��˙����u�m���v�)������e̹Y�se�����'�W7�����͂�_��t_���k�2)��gO��9��e���*��qy�/Y�u���z�C�]��)�WG:�y_��~���|s3���l[l��ْ����;�G��f�s$��w��LOήL���0i_���W��_k�|��%�dƈ�\�"H�9���2,��)���8p�,[k3)L�P�ۺ�w\y��h�A�ƕ�W��_+�p�,��x�ǋ\̙f+�ʋ\�؃��]=w�iuw�\�[lS���O�����j��^u&�λ����I뺅����,A��3G�rd�a�x~?Ëd�[V�V/s"�/�Z���\̵7�fH,��"��ڹG�e��r�H������H$R�H�lD�(�Te ��y�VR��a��yU���3�p��B��Sz�I��yy�����������w�w����:�[i�a[Sm6lA�D�	"C,�f~� � H h�
L��Wyz��4X���C)�	��@䡞#!���_@��F�xZ�5��ۣy����u������ - ��k����k/֨�=�F��T��m.Ŷ�Fl�67��-b�Ѧ�M�CƋT�@��\ngn�;�]P�����.��`�gLsopӛӜm�<�4x�ק�{�~|��i��������Н��W�Bz�hҨ��`/���v�u2����XE�'����8���԰�p�VC�V^�Wj�#w��b���?�j��~Or �c���0��yaz�~��U�5������SU���ʅsW�W���n亵�m}a�������!�VN+_=�U�i����ox��YVvz�`���ZW��+��f�^�+��SP{-�-ĭߞ���;"�����$��GE����"l	��.	~�@��<�\��
X���!\y�Xv�^tX�!��k1�WE��-��Ϫh]�:�T%�	��j�5H}+��}�O�Ա�J8{�a	�B��m���2':�l�9�4�^_s諈�;�L��J�^$�Y.f���o2$y�Ů��v��-�]ٻi?=� ���y��zH}��O���~�W*Z�9���$J��ƓӦ���҅o�&����ݾ��[ђN���x�k��{
�#�K�n���o)̬�di�J������i����#�蔋8`��zu[gnd�Tl��.�Q"恳펥K�`>�b�X�U ��-#��!���>2ĭ�y���=�ؤ� ZO��ؤ8��p�E��"�·F��/�p&GU�Ӭ�ۉv�5Ϙ��0g%�5�R�>���Dc��S0aJ�]Z�4K PUdim���q�t�������Zc���۷�q9b^�n����}�쾝���A�_� ћB�9�??4�X�����a�(ƾ1Ã\�hn�͗���jJ���7��A�4���򤇤�S�`a�˱�P�w�Ƌަx�j�^�H\^���**�s�kdK�^4$n�a��:�d��G�����X��R�<�i`}����؎�WA�#=�p*��j��N��� P�]f�����q�U,�A�P֫i!�)���Z�uhv�R�J�2q���B&�o��Yt�|� $� ��Y���j���o��n�@ǹ��j�j��
�t���.����1��n%���#�(����ˏ
®��^E�08��U��ɲm�U��U��-�����A��r���=��XM������k\��*Jh���pa���5��vv�<�u��:�����]�y�H2$��l���#�k�3�݄`!
� |�|oå�q@���6y9�Z�9MեJ�"����,��L�֨ _ͻf��oGx9�1��C�6k���N�{�X3	m�cJo�\�e���{�m���}��H���M��{֢"�cSպ��.�P�o,�{甖�)��+@��!�u���UD3�����6����������޹��D�1������jyuM� ��h`�g%>Gw��qM͸
Gc�ة����R�
aH��(���ST���;���P�u��hHra�fY��*��$Ǣ�x;�wt��yW�r��C��q����&Q�J�0�0�.&-�&(�0���)4��B��Μ���ֵ�%E��^m�o��#�S�,�8q��vsފ�kqn�~��@ �H���@@":��l��T:,���Ơp��}�/��{!���uP�X�v����@�|�����: f�5��'��M�����w�v�ڙ�
�*y���c�2z��ܫ�#!A4�J�ǀ�?\���g����~�\��c�}�ϱ����P��"̲�Tޣ���0���j���YO��Oʇ�p*�S�����i✈�[/R|)�c���`';�0�:�x�z�{�����GW�u�h���\?��}s���o�Mt��+��è�� �;�G3��OUkU����A���W>s�D8�����{,]���d�e�u��4�p�O˭^D��9�
m�m� V�ܷ���5��e����c5���	ӗ-�|�^	�B�G��Ԫ�l?���$���#�b$$ ���Z�/S%z|����XO�\�o�܏{�s���7^�oq[���DC޶��;�P$�k�_ܕewM�XU/�!O�ӯ�2Q���!��&9(�V3x�;�E�՛cft�Zo
���a������A�u9��p��yu�u��q���:�W�7S��-���.f��]���it�N�΢�9�˒�_�,�1�6�M*�0�Ƙoyo�[���ո�~]u�?�����q@5n�rUo�8�*�0C<3��]3�[�S�)n�ǻr��5�-���}x��w�ںN��* �Y�^z�8��oHuo�נ0�4�ｵq38d\�񙨗i�H@1�yh=�1ug�n+���[b�{��H��E>bUz����l�)p�g`4.km�󍬟QJFv�us�UV�Ӟ���ʂj���}�;��|����E��5�v�FYp����fE��.��g����u�^�a�,�z��a��i��G� (zj�k[Dp�fn���rw�ުg�s���n����A���:�T��c�i�����Z��u���$�T�D�����e�9�x8�	S@0ֹ�nm���jړ�`�I���}�.�� �߼Ġ`�4J�[ծ�kUf߆�aJ�����w�iMF��WO����Sx�'B9 T޿�*�Ym�Z⵶*3�I�5��a�1r�e]v���N(\Z7z��T�3�UJ<P�{/-�﯈��1K��3CU�y�%x�Rܻʏ{T�S[#�{{��Q�ٜz��v��2d��&s�{H=r�j�NQt�p�^�W�{߀�\����u�^[������`s�<��agn���}ׁN�7@�VQ�D���ֹ_��V�u\����p����6(�����h7�w �g��zw_��*��\����ЅwLmÇ�On1<v��������f�Ĵ�7�X$�aV�7��fki]��vic+��w�Z�`m{�dA~3"��0�)�%��� ٕ��O��gRD�dIν�ǧA��n��j�u���(sxj����f�v �S#x��V�BY�Ӷ�XGd�L_�R�������Ŋ�(� A5�ҦƸ��p�����莇�&�.�3�,geջ��5�z�4,Y�*ht@��y�6���oj;4Žx������+Y�0�{���.�>�إƻw6�j�����/,۸R���C��U�މyz��BBJ e�v`�z~ |��Q�|�,�]՗/�,t� �jUP�QR����a����.*�ޔ�Pm�55�~4�Y�-qX�j���]R�إ�u�{�_M\���Ev����VZA�r�Y�R1w[�hN��<�}m���| @ ���y]���蕏gr��v�U��f�����t�Z�^��>K��eT���Ӽ�uK��{��}>�zbm]z����T�B�Y��5�x���ZU���Y��?��8n�+鐩��
�����isjS�d��m�i���3���U�U|+����ǃOc���Mq5�h��͢��+�2�`u�Zj����z)\��Q��Q�.ͽ�w�C�M5%�=�߫Zr�Co�b�N�*����f ��ʨR����������o��T�g�a@G�l�TU���T�_�ڐ�V�H쌂�yNb��'ԫO��'�G�
UM��Q��Od�b���s�
�k��Zt3���Jm�mj�淺�zjD�]��Q��Z-\�@}�@�ә���0<�� �U�֊/6��ܜ��3s�tl�q�K��\6�y/�r=��{�v-Y�U���b	���W�-�aTn���$�0��lN�:�Q�O-Cv���Վ
�ה�5��ѨS<{�~Y�'e���\Ū�VaKj�ר�<<.uj�Ѩ�S�H˧Ð�U�C��c�^"|�ޕl`�aN�ӻ϶6�]T�5n�� Ёl�At�a��'���
� ��h���;��~*DF�:b��ɸØ�d���$�eGXCa�
��M�mĤ`"�T���ېå�������͑-I7�� ��h��dP%w}�@?5�S��`O�	�7gLcz�N���a��+ �Ls�ρ������, h�~�a���oYon=�\��v?�z����/m�Z��/xS#���l6��?���ј= .�(�j�N* �kL�%鯝���١�4�	�@��v�ς����y�@k��4 ��CV�u�C��>�-!m���3��;�K�|���y�4��;��7F�xk]Q���Zt��o@��K��R�����/Nt��U%�X78�[��3� +�i���qV;���TZ��M뙾�r�=OV}	N�EH����@�l��d0/7Ysz�;�E\���@�ݻQ=��<^
���m��v��g��a�gƬ$��hm���WZ6��I9�j�X��]3�U�yb�XSZ�6���UW4t��A �(���F��LCk�s�a6���K�r���pyeXS��l*���طf���]���`�r1
s��ľ�N���9��*�Sf�J��2�3Ww[�ֿc� �d$�����?��0D,P^���I	 6���~CÆ�����Xm��t����s�m��Ssq���׬�ur�Ż���d.p.�;��3�b���"�+�C=|jF����`u��o��� 5���<�f���Bz���C���y�W���(c�.c��myֻd`�po7����0N����U��	�i�"ڕOZf;�	�9+��[M����w9�=���ˆFي'I���]�LF��b��go^� zU��i0,&i@l.�{��T;.�r�[��y}��)W�[�=�g#���gu�)�GS�]�`� {��#Vf�3.��n��"���Ag9Î�>����y�[�Y�e��f�N���
ʮ�J2��tZm��rx���P�+�Yk8.	#�hZ��Z������4Ժ�j�J_�H���G_5R�噊���ԙv�}p�t�r�7)w+I6�{���-Yg�L�>���R���2<5���,iM��]�@���B\=�-A�û:mu��J��bnS��T}q��h5jl��$ܚ��][MRR�2e���� 
n}�C��t�B�n���<F�8�@c����j�����<�8��{S|��G��=��oU�c�}���Y��23T�6씵V�C1�o��ը���Mz��`5���r�/��W�<!I��#���&�(�I�M���Q�x��`,�k@d���9���(�<D�r�ki��0e�\pr���-V���"���=� �å��p�V_C��������Ep\i� ��݃U7�uhB�Ȭl�X0�O��u=H�/�p�7�P��{�9�A(_��BsB;��j�ݿ�\�wЭ�@�X\�k�v�bꙫ$TW9}��X�z7��ܟ.z�ч�ai���v�h䳟���c2�����K�3��3���i��回��0�E��"����ԉ]a�;��H�����Y�4�λ(��}>Z	 }� 2����t���y�xC�M����4}ϥU�	�xĲl$ɱ�<��xE�w|�@����98_]ͅ��lrJP���U|�H��jX4��2���]��Qyuy���%��G�JŔެ��H��N*����;�(H��k']J*�t��8>��m��ξ����n]˼Xk���1��7���V�fu��,��d�eŒ*�+�Nk���fC���w��`��i�BB�0fv�Y�+��]V�bī��v���t�eL�ס�_���%|���S�UC8(u��:޶k�_9�H��Y�%>�{���ߦ8�f��Y-d:�`���a	�C��p�n�P���P�k8w.��غi��
Z���ۡ�&Ԝ]Vb�q��+6�J��j��ŕ��Y^7I���1zv�ad=�\�#p�'tZ�P����{��ͨ]��F����i�9b�sG#&����[6��F�m�}��҅>�MT�W`-R`��B�+c�yy*U�);#��nEkW*ͫ�4��u��]K���<�:�U\q�nggT:����*~�y�<�i*�Z�!��f^����ԏXё�d)���tҰ����q�0��"����B��ʶ�"9Y�Gkky��˽������}b����{1�UF6��N3S� .*�X���qU>6�{}��1O�1U�k�~i��M�6�������s/�2վiZ{�=�roqAA`���
V��薅~���£�кգ���2I0t̖)�F,J*����X��e.ta�v$M��,�>*��ۋ�f�8H��o�9�*���B���U�:�I7/`oE�Y�$���N�R��f7)����â�K�`�`�o�0���&�09����o�a{�o�P5)z�P�K�l?E�F%`5~�s_>ܶ�S�����<��l����[qr�k�"E]��d��B�g.اǸ��w�S�gF��v�o�!V`�{�����GR�<����])����P����N�ң����xЕ�-_��^eu6W��L���c3h�U��	Z1k������"�M�i�B�1��u�>ٜ�<��'�����es�(�7]�e�KM��wt�g{g��_��c�qƞ���Y��M�'��K��V���żzF7{_�����v�nv�T�yZ4-��]�f�YNv7f��E-mEzvj�([���Y�-+�q�]Y��x7�kwo�qS�j�_�g!��F8S���8���Aw��ƷX֣�����ѣ��N�Dް�Wt�{����1$�ޛ�B�����UM����u��ݡ�/B�UG�e�������=ndz��u�=�ӫ+{��ȱ'ӳ��������CA{0�)/���Ŋz�_��:���彵�dɿ�mU[j�le)��Ç�ӇܠvۮI�Ŀ�(M�~�ɼso����e���Ċt��ӧN�r�l5�+3rŋwv����O;�h�*����)���8rNKl|vǝ�0���b���^>+�d����h�ܥ~W��N�8st��j��j��!�\�6�����Ç��>��m�m�V�L��(��Y(�.^Y��yc<<8p�Ü�r&w�p� ������ox[%�YQl�Sç�N����+%�����&F�G��ָ�\�F=w|L6zl��Ç#��-3�2ʒ�F��&L����^6��+�w[���Q|sj'�׽�ʫa�yVfkI��~ʤ&
Nc��l��Fv1����X;Isk2+�X*f\�t�_V�WV�8y���x{t��/5nv�>�ǖ����,Cv�$M
8H:��� ���kS+�t�qQ�	�]T��,�&�i�B���pOR���<��SCg)6 ��=�2gK�����[O͌�y��0ʏoCb�y߀���~R�sgK�v��Ms7�����[tgg+�������n��
9�A䡔�v�FoV�$̫#���?��3{�^?z8���X�6
��!��ҙc�@P��q����50�\5��H��Ω��16����������3�]}8����{���
�5e�2�M��2*�Ds�f�u��,���N�G(��}���$o[A�n��&�P|��h=�MO�J^�a���/�bP�Oq��_�*Xz����7@n<f@����ۺ���t/[���^=�Z�j�2�Kc��������S���m<D�n��۸ԛ��$߮KϦ*��l�|���i(�J����㥛��#��Fj��ϦTSW-����$?h ���B�b{E�њ_J�{��Rk��w* 6�5J��FCΑ��b��+�!����N�;O��%��
�N�� H �0�9�fID����ԅl��$u�i��M>��U�ՒuX|��)��ě�c�3�x����͘�s�: ��G��"a8]�4�R	��anC�[Arn/��q �@]�N���|�Z-�5�O����@l�|Mt��D���y����=�x�Y�L�Jwh.�X����}� �/�޷�������yu���0E�J�=�W!��m��g���ᨁ�{r�&f�4���8⒙��5{�l������w�Y��öܩܛ~V_��C��/6j5>s0�W�<*'q��A;��fJ��Y諦g�s/�,Vf'��L�H�N��Bp�[�o���~£N�ǩ��h���<�j��Mp��n�@�1�~���X�J�����&�� X����ң�� �:P0�j`� FJ�,�z�v�mk���~����T5,ʗ���%ٳnC��y�3d�$$�W�����(�ԥ��G;jr�;x8�h���"�^G�Jї}fq��3V��V�;9]QYk�CXJF��Ew[LR�v�2��7^�/ulN�.�N��e�����w�O^+lcOZV�1�1���Oшa$�$�FO ,!�?
�j*�^���h@Zl�h J�N��уc�|U�&�H#<d5(���,���7gvGd� ����0e��x�g�
D�W�h@%}�s6>��[(vM�hH]�oT���
�)󫀡+��tR��(;�/�����W��eD�mլ��:��Ly�L�����i���]�Vǔ<�~��V��'�\Ea��"on[�f�9�"���߱Ҷ}c���״UQȍ�oOTf��{s�
��B�@���3¯C���S�K�s5�0z���y�W%%On�v����6T��Z.c�B:�#�*��O6�O�$����spk��;{ܲC����k���Q��{ywp9��Q%��Mπ�V{�����F�t�-����Y��Ls%�dm㍭�[	PQ�����@w\cn�L��z���-ۯ|:���j�Q��h����Z��]��h�*d���k��7=����7X-�;Orbn����O�m����2;ߛ{�_����y�K].�K�u��IKko-���2��q{t��XS�Ã�t4��M�˦��bv���]LҤ�3�!�)��7�h_h	s{ �Q������Oˣ
٢�bN�Cs 6k�I�v��5�Cg0�6@_@:�"�!��c�h5�Y�݈����wj�����7(�d�iL�2�ֺ1���d�6�H�&�x���ؒ�T�f2tz�Vl5�<C� ���5;���XήEBF0� �;�;�Ӎ�m�MW�x]���B���ןD�xU_�����@L0����J�s�����+b��Pf��v�n���EL�����(S�(i�s���E��,�n7dH�Hӹ94�V�����t�ǐ$��S��7Bا���I���jJ�UL�V�a�C]��@��2�@�c.��2oYbKQ����E֗�.�gN�g?�(̋n�/��7Hq�UgT(o�5%��
6s��DS�۾�f��	��)֡q�w/�����Y�γUZ����uYLPY��ϲ�o��E����b]:�<7m�̭i��.g)���擝��h�t�+j�sSa�t�l��U�,_�<�������w�>��Ѹwۮ{
��J잛L����z.�'8F�1�;W�����Ld7'ڨ����:�Ϙ�u���w�Em�4z�U���''��sL܆u-�ݜ�r���g� 3�s��<bT��l��.&l�}۹r�l��\��y�q�'6�Fv���KS;���;�Z7/Yqa݃ӷ��I[ػ�lh�cd��h���J^�އ�&�N<fWl��*�jR�}�6�PB�n��M��kx�S.�ɼġ�T��Y��n<��2�}]&\����4�@�`͡m	'l��k�UGOhmX�|��`��k�fWX���spϏ*]Pc�vK�ġ� 1��EUU�V���q?XƐ���:�wdس�{K'���^6�A�����J��I��>�Op��0�����Q@��x��z�\���8��b5������t���c{`<&�K��iQCw�MU�~�e'����ue}yYu���O)���U�]��G�c��4��e~���?`:�Ǽ-�X�vo*�^>�hT���o,�X.��| �1\7�������I!�����{��@������J`{�,R��o�=�����<&�@骰XzEp=z�ʧ}��a���z��ÏwV�Wfg�x0�3�z7�xR��xο,�kWTWS��h톪ɧ���)أ��-% s�i2W��7Y�Y#���}7 r�����IfЩ��Ǎ���L��w�]h���;���;��龺�hf�Vf�s��^����^l>��U>@`����|�X���<wq�=�5��R�NU雍5u�s���t]��v�%���ȓ=�g�~�]��sl�_&/c0.�,��BEh1�k���u+Y�$5xk�y��v��lŞ��D��6v�U��#'�=p�W�H���cN+k�憃S��[.�q���"6�����W��[� �ׅv���c����Q�-7y��i���[�5Z(腽	e�T��8o�4������R���ݕru��c��cx�4ѝ�;�J�x��*\TI�!	X��������]���P]qZf�
]J�QvY���w��F���It3:�c�Oz�4�Q'8^��A��QL�5Qű��B(`���b�l��<S�𹻶�癹j�;;�~/�����j��K���> ��y����)���ɹXx����w[$�P7��q��f�}I8x�[�v1s���@Y�J=Yϛw]�Mc�_nG��h�!�k�/6�n�Z�d3���E�vb����H�lOS�s��-׸>�cH_�ꯏC�{�Xl��,F�D.����ߣN�6�ð��S��Z��U3���ݯq�:ʤ��L2�!�^7��'�ly��i�#�{ҕ��#���������?�8��T�5��yݚ�2O9xԧK$! �3>{���l����QJ|UM�T;.LZ=[+a� ������{���j����@�I�Ttz���������jOk`�F,���Ň�}_VU�N���ǐ5 H��x8`8��38���Ƽo���n뒽z��,��
�ME���RÇ�d��>ȽqZ�sKy��nU]�i���P?�ë�Eǰ��z1i-��12�8z���o0�Qԗ����^� ��\|U�FIݘ=S_F��r���v!W��(��`�#���9�P}�pخ�u8�qX��lo�q�w��p �j�����N_�>�!)��=@ml�5 id��t�NC�l��E���v�MnB:a��Y���[��4�\;s�@��~Md�1l��:�>���\�^��)�r�f���]t���P����̛�W��1�nR�k ���� t���p�o�S�{jҠ)-��=	�i�xƼ�֯T�\��8�C��D2ɘ;�ud�y���@]��S�]��P��i4x\�Op�F���&|}��@mN��G(�.�s�U����j���'78���Ɔ� �z�7t(��ʀR�)dh�n�l�1�1h;:��Q�8�1���p�:�����о���� ��ȧ�;M�uۍz���9�$��ܱuMZ��"7X��B<vYahx�����W����2�ς��������Rg�@x�`��X�l������Y�}�|�������5���s�^�4��������X*K�{Wzwot����q.�v�@�����]95oV�J�1�����_Lk���7�ؐ���wp������5�#30�4��[V`b�%�?(D�Mae�^]�n��Z�?d1��c���Q�y�|ޑ��3d���X*�kg��[�s���mWp����5꼎*=4��:�l7s���c9�܋[�d
��L�(^.��ŏ�z�#�̰o!�����}j���A���ysM�m��\�º/�����"����{ț�j�m�W�>]ó�0�)��� c�l"J�X�n�鱩���'��%�0�0S^0��팬:dq��� n$��h�������uy��wpkTG.si(���w�΍����v���Q�8Y�";1܃�򷾼ZNFi�2�< P���/��x�/\�ǝ�W�5���s����f�Db�� ���=�Ϛ;[ـ�C�7jw�C4^�V4�S���L��X#s�(ou����r�4�*W2Xb.��2����Ue�-�����պz6L]}2��w����~���wR�-���Ȭ⌁+�ɨ=�}da�*�~�!��ʛ����R�ڪ^�$��3��t<���OO!X�����U�-���-�| ��`���'���[��z��ʶ-�]?t�>��w#ϛ��9�^߸+�	A�c�mH���|�ك�@ZL���w3~�frb�l��-����!�ڜ2.�d>s@A�1	t�ś��VS"<��P�Cr�)�L�d�� /+�@�lhks棲#�@x��껀n<���k:�Ѵz���O�5ǏS4i���@K� ��HY�tW	���[;�����j-����{�Q�9F��w��Ԛ���.S7}/��T�'�|�Rw���p�ǩ;p��[+�$X��q���{R��45�4����6�� ���Vq��K9����)ri���|N�C̴bc�&n�%��!��#j���`V*�������ĕ���U�����n���b������^.�׀6H�Q���ڼ�x��C�4j
ȶٹ�����*��ۓN<�]���W�VZx�,�r�MU$q,룹'%�ЌB�̘Ի}�we.�D�2��T�C�mf��N8��!j��2�5�3G�ss���0�e3$ˆ�p�������Ӭ�le5b:����֘�7�\��v����Y2!b���YU�[^6�Q�*[D�iJ>��g�j*x�L�/xߨ�y�CF	.PyG9��W�Q�ǉX��V�,ºed���(j1���j�����z�,��HH�9�Ғ��b�JY\O6C�J�6#���˩
�Z[�\봗C6]d�֖$�}��S�h�L�n>��gL*��-Ok�՞�Aȳ:�>�e����׭����B�����5�-�/{1��f=��LE�7�ܲ�[u��P�y�ڭ�J���;^,K���J�2���r͒|�2m�֔=j���jU=���wYm�b�v�!O��Ҕ��i�ܫy8���[6�-��J�j8(8"��R�c�\iI���q�p���u>}iSʠ���@F��2����qZj<uls�V�広�}ݦ�,��bJp+���+����ơ�鲜����0���ֳ&���ꝠѺe��U6Zо�I�R�}L��8�vR�o8×�-��w�P9tb5[W�u3�nGK%����z�%hb�KbU���?����	!�y ��ah:Z����b$Xj�!L?0�$�ª\B�݇v#p ����A�A`D�H�n��P`��!����¬a*C��C�&���$`X1A>VR_wY9᫤r��k!�%M�~�bA@��ߋ���\o� �:�0G1G��\���������)���;՘Q�\�
�ӎ�H�ʆ���P�e�W3��Mp}�M��L��E�S��d�1�3��K{�}.cu��b�U��<�"cVV-�I+X����a���K�8��U�T2݋y�m�aݪ�u���.է�u9�ٜM�D�A�CXgj�8%#Re�{:
�nG\�v��U�o0�����c��O2v.ݾ�1�dތ��ll]����֠�t��pgd��	&�1:�*������峝&��d��֖w��K��#܎�+��I���.�����r���:�yWv0�r�1w�kU���H�-W>��$�M4.R0*]]qXXtu�t�c�s�HT�sl�bD�ma�wX���)�tt]��c�H�qU৬��զfm[��69ae�ֻ%o �/tq>]3^嚉$C{�o�����u�]��88WI��t�:i���]mۡ����5���=v�����Q5+I
�y���mWI�qi
G)om:X.�U�1���1Y;��fy�ɂ:;���)��*�j�<�Qo/�{QfK��`�>�u�:����o:r��q�wl�|��'.�$�݄_��X�DX���^0��:���i�V4Ǌi��b�h�i��i�[|��oO6����4�x�4�Zq���`�@���Q)eշm-̭jҠ�u�/^�I̴RM���dA#`��Ԫi������~/�}[�`���F���k%J��e����������6�޷61���V��e��)�F�8p�b�MfU|rG�rצ+�x����9r�6t��ӧND�Z�����Qnk����5��Rщc6p����Ol�IF/K���[���hѨ�J\��-�)��gN�:s�e�����F�$kx��h�Ç8N-��J�׊�6�~�7�m[AN<8|p�Ƕ��#tn��W,��N�C��ʌ�M:t��v�{e�j*�̱)���"�ؤ�}nW��+�ż�F��\������	�?s�9DBg�	6CF%)���ʱ��:��m]��p��K������$e�e_OJ�w�e�$�pnYΜﶩ`��Q8��'�p�W��6�ٌ1U����+0�#$�B��7#`��E�@`�<9�	XLX�\?��9���p��{P�ǘ Mm�{F�:U���G:2��&Z/�8�ڰ����d��#-80��x�j��_���_b�rs���q{"▁�.��T��ϒ�]c����Ɯ��}�N0'k�P顟��q���b������A������dg�*���¶�����on]���<BZ�U_�{(�l�� ����>(��f���~ �:���!�Y2�'8b��Q��a��1��:<��%}�E=��굢�jֻ����bY���;y�����j��1\U��M��x�B֔,�Ho�!��
��k���>?�Yx��Uv"X�EԋuX���7��t��SM��>ci=RL�bO��7�u6��|�r{Þ�p%����<q�0�p��{��9� ަ���ߎJ�_�s�[�p+�������/�(�������]mU�V1��2�(k{�{�r�]�)�/�,�(<J.��h�-M�U�M��������^\�kh��t���T�V:�wq���6�J�IL���PvKف[�����x�?���f��c3�w\ S����{����^�!�����g#�"!��%�␭�|��9��pdy�h]W��Q����챔ٳY�ƫ}e�.��Sn��s-�KlT��u��k�n�:5�Ľq�ΗIkDbm�@Q*U��U��q>2��z�/���J��ҕ}���X��4�����'@��[F���-��gz�;(�eZ�^��	O"zJe��m��2;6����r�߹bE��|v|�qP��6^A���0;<���Mh�
�8́y=��;�v�"W25���s\����9R���l�z��/����gW)�3�0*�X$�eY"�Ui�Sٺq�/F�	m��`�[��E3Y����[.dM��SՍ�q��.&lR7a[)���(|pBh�w�΁��>3�e��?��/4�][+\z��KC碳��yo�-+�ǅ�W9V�[W�0��o�BT��T ��YދOv��y��_!,����2���Ŝ����i5��u�!\�����z�Z�������w�+�����	 |���5�E�:+��\�S���)BP������w���y��9WfWV���%@���Gr����i�#��ڥ�5��Ԉ�z�ֻ��!�W5k�v\�,�X�j.�5��}��BT8N^e��^h�<�VWBS0�	�����	��DM�ո������Mʧ��(z�Q���� �+߷������z釣�b�&v;�
������;v�j�P�K���\�oa��n�e�#!����w#�����/2Գp?������l�yD��^xJ뺫X�>��U@ʶ�=� �j�ׯӼ2��18��Ǿ����zsz�V�[B+i����ZUP����	��s�d���-�=�On�*�n���x�a�����m��>݋�0��;����%�gwH@-4@a�;�<E�p;r|_r�|*�L�պ3�^]�ˣ!��o4.ԍiMS�(�40i�����{��Sf�w#t�Mn�tɤ+F�#���6.�NyWeksZR���k5�B
�XS�YӮ�&�����C��']�,�+����E��]3{z�*3�X��;�z�ޝ����fg؍�^��΃P��O��O���@�w�v�����XS2�w�{����OF�f�ֽ��}��Г�Lٰ�L#\��dE��<�,o��,=��(�
J�OZ��o���|�����ʊ6^*���U����ޗ�����p򦃚_�!ʣ��|ymIUԮ���N��Vs����J���nTn1�g ��Ƽ�}�A��ô�o����]R +Sr@Ƒ���R�sp�`�8C6%�/S�#[H5Hh��Qn��k<����O�x>u䁀�2�Kn�&��&���";|i��x?Cy�g�; t7��[����9w%����k���HZ�	0�L��L��K���*�
ֹ�j��Rj����QG�K�H��F�@�YX�"�O����k�:7�n>P�C/j�[f����m����Y-d��eX�aS-8p<UMaȧ�����횭����C�	h���Y�0Y����r�r�&IQ��q���5��b����V%̋J}�f��N��fa���ⵉ�]t���V�«m��4ccJjkZ���$�N| �?�b�ݯy��������h�y�f�f��S����Jb�1;	i��#��"���.��.���փ�=��C�w���]J󔮫���[70�,2��\Eh� Foc�h�Z���腸;����϶(���=[�Ȥ��u4���	���7q �:�6���X������Z#
�.���L�bc+:���h��7�k�>sl�@?ξ!U�4o���_[�w[s�)b�[���ZF� �-/�K$��1�U�eխT�ȁ�Hq�i	���q��@�a��V��\�? ��2m��Uk���-.�]��:���J���1^�M^�wP��@$�VQeYK}�?��~�h~.����7���Q���U��0�`ܩ�3%��\WdU��rTP��9���>����#��u����}������o�G�Se�Պ3h»�I���mm��A�i��An��x<�N<��g���n�t��PX�3�z;w�u���٪�2_V�@�qݚ��dc�ת��j�͛k�uv��ٲ�G{�+R�Ч���U_��;���������}L��k��~�!<2��E��p�`��Œ��������Cv�q��.��n[�f�ze��y���Pإ���_��C��k3�?c��/��ց�YU��~��Z���[3�P�%�N�������,��u��Ǟ]5v�>�͟D��Wl�c���9�#���DT�n�Iw�M�a�e��c�/]S�L�t����*D�
a����7��M��!���]�y��v�\�P�${X�X�;��+�8Av~y�4��@� �>��̟zvN�����РK[>�@u��[(�����w(�:|��r-Vt
ʥ���<j�d������l�Ԇ����+��+�^*�^��v,Y�x Q9v��=)On�f����]v��Kd1�O")�aH��q��7�w�$�1�Gpo�����%s ���Q�1�{�.�-'���&�r���I�Қ�K��a�@��'���5���j�jpa
���w��h]��&� b��0����Y�ɞ��L�԰6gk��\VXԍN�1�]ԝ��0�eX����[�-x�}�x� ��xS�U-*�R�̷�����^���ֿϳ����v���t�wg��������jO'"��$�G�S�!���di�n�ؠE��uC�^U���HFZY�A����զ�.�e�0pe�D^u�]���`��9Y�zr78�W'2�B�V� ��C˶�����ш�=59 c�a�{�+0;���x�Y�e�غ)�n�{����=Z�c��T��Z��W�mW4,��(R�Wʱ��p$oK�*^2�����Vb�:�춖ֲ�=W B� �P��c@�l�n�r�!��=�\u���m��V�0o�	�k[�DO�ł�tEW ��������0c[��oP���1��z6*D�fu��n���6L7��uC�t��L�$M�"��/oJ&�:��RMMױgNu�ǌ�G�i��X�0�Y�z#�X<�������v>�K�p��̈n6��ʎ�r[`�ŻfN=ӥ.t��~�	E����r�G��4M⇕�9��:�M(���N�����y�s{Y,f.r���s�U�����y�p� 
(@$�db�Ϟ��繻L�	���k�yZY�]�H��_�@��G��[��ʫ�
���|�Ne�v�7���.��cLp{ܯ��'��O]�fi-�*k�+^���]�z���c��x~ЀY�
�zQ���#d��=�a$�q�%1�P�E���N�M��D���`6�}�V otf�6�؎]tO�Υ1m�sm�<
7Κ�۴����d�qa���I]�_���|�
 �3������#^�
KW6����@k�h�`�h�˦v)2M����H����dZ])rKv��\㱣'h܌A��E3��W��]���J ۺ����둸y��5P�*��GL��A��8�<
�Қ�L3����#�p&3q̙ H��w��[T��w�y��5p|FD�vp_f4"=�;� �i�{���m�S�|掮[X�-��֭�p��{�ݘV���q���4���9+���gi
��%���z�Y�_�^��M�i��Q���*�����N=�MV<��o���h�,q(�yp8u�*�s]�o(F��p %Sl1�k�n�f�u��~�JHR@�P3/Ƒ�����>v0`@�P���-�2����
h���[r�3u�p�l�7lSќ��B�e��w&V��M���2H=j|M�N�~�oFKZ/��'�����EL�k�Z���*�g!ĵ_�`)����Hއ���YbE(�o��MkefV�i�Q��Dʎ��� �[O�]�4�"=t<��oL��BC�4���Vmp�[��Hw@���͠��n���ov��!�X�L��37���S��{�1,�UM��p�%b�m�Ff�F��b��F�<*��[L�p^nC�Eh~��x��̝�� e8{̦B���e
���JV:s��S����+���.��\	�~#8����ާ���N >��I�6��W��� Ml�� ��i����/y�k�.�=��Ρ��\�轋}h��Ȩ&�3��+��:]��+�D6���S���>8[wU}"������fp��v�]�UU���ۭqN�ė�C��ݿ�=�`;���Ly��ϞYw��qT�arv�,jWWolOs.��mS:�]-���۴�y;�^�ߵ�쿷촴��~fK��0	��ڳ�#��C�Ϛi�S���i잀�\������^q�c!>���$��sw�� Rcݱ�^�qX�
���0��Uґ�략���T�+a�[U���s8>�S�q�2��Fa��<e�F�>Mn�k����sQ8���ᅻr>����]�z�l��
����`8^��C��� �E�|f~GY�7]��e�]k�l��������� �=!��a�2����Nq�]��>����b�7���ށ��π�1ީ�M"3M�� �e���*�NN7k(f��c�	��@UlzS{�}��
A(zm�!��^�
<3ph�9��q����� �nU!���&����!٪�c�Ɏ��5�\f*tieVSW)�c�Uz���^��]�~��m�.���=�Lj���-�CJ�iO2����y���h� ��a":�Ғ�17�4.�J�N�rcS�`��l��Bf�|؍�-���v��o1�(��bt�9ŶӘ�ι��jxx.f�Lb�TP.�,v��۷�97��Z�Ap���0rP��U��s�q�N(���
M����U�G�t��|ْÆ�����ꜻ'Tdu�%�wi'�yz/��U�4]2�ơӵ�/��n�kΔ�J��1�}4���}N��ĺ�:�3�B�t,�N)�m7k�t��k��ٗ�`�oibtjRA��v͉^+$hࣧ�y��:W�kw�ͼ��ꮨq.�f:��]��&��5]�%�/VC����o�ӻAKF����rz������w�Vmp���:��j�������h��5�j�wd�������uHtS�*�)�kV5	�i�vz��V�q��P�c�v�4o낫�4���O��ѣ"�k��v�������J���o�`�l�.9T`=�a�=���j�N\G ȫ�7"Eo�Y�MI;zS�Nc�ػ��Z+v�C��<M�:t�C�e%R((1��깗�8�-�+��mWt��"9nv#0��`�֝CnX���"��Q�ud*�&Kp�	f��6�mz麨���$�4bʞa��X�/ ���G)��C�5��:0P�bƄ4`� b�Z�������A��0_�՛�W��� A����韖�Bz�e�����.�I�@��y�9���y*��C�e��Dw6xC�sZ�cʙ�ub�)(��/��*vG}������܊�L���ʊ���\���*ͽH�w0>�����t޹z�U�jY���zR@���vj�3)=���I,�3`KE�,��t����X5<��e�lD���э0�C���b���.���A�f���}������SB(�U526��wnL�9ցT���/1E]]���l�ّ�;�\��fz�'��6Xj��/��מ/7��V�Pt�[���;S358i.�Be���,f�}x;˔p{�&���<}k��j�8����K����x���/q2����L��D���%c{	=����ː�Nu�ShڕԤV/��tY͎��hVU\�˸�q�����ޒ��]�5�,�,����B�˂��f�e�-�s��X:N�GK#�.�*4V>_�>{�8�C���*���[S%c��	ϯ6c1�/jOE֒��opJ�R-U�Ee�:�m���d}ybWuG�cN��.�A}Kk�[��E���.Ӆ��L�Uf��$�I�AX"
 C�I6wo��g�dņP�$��Z��b-H��<4x~�N8�m��h��q(��6+x�?)1aN�<:t�Ӓ}\��b��k����vѣ4Q�-�[=�,��ӧO��9��վ6�v�QּZ�~/ajS�G��~��}ĵi*�f�oǌU��Z���m���S����N�8��[-�-�ũ�e����>̾d��bh��ӧ�N�T�U&T-�-Z��Y*����0��Ç>k|��co���\�kE�k9f��z��0�gO��8�������W��զ�l�vv���nj�j��4b����������z�i�Q�:ru��ޤ�V+��]A�6�*O{1Q�8��>�k[��U38>�T���2��N�e��_O~�"�KKJ�R�ww�w�˝�f����^ݣ��g��j�]o�M�q��4�Sn�n��q�q�Z��Co�M�~WG���pw/°A��A̙b�߹��q��9��1���T�p���y�ԫ�o�c�F�ҁ������1�0���68��!�޾�@��@I� ~O;տ�����*�;%!A�LO��U��a�D��E�
�_j��FW���z@�U��`��;]�xML���bd(e�9}����R��;{ ^3�Y��q��c ���u)k����	G�,�&\��֜#op;h�r���"/I���h�39�a#m�a|q3�mx�T���	I�(�hx�����i��'y�LҜn�m]�o|�z@�1��PSi?�`p��c�9���bS.zi t�_h�HF�k&�6�Fi	PZ�2��S7N�Xc@;�p.p�ɳ�ԥf���[�m1�o�w�Z೟��5����D`�2�]��L��]��6�/PT/cLU^��P�%��Wk�ыrvs����Q\��|�>�+Y߲��^lw���e=K]7X�����O�aT�Z[^��?]�~wS?C�텲�jx�H�<�M�x��V���(�h��3u�\�Ɛ�(E�O���0ϰհ0B\�j�����Q�@827���s52�Xa�l��1ƯGq�菺F��v3��w��\�]����EVa�̭�1 u������5۝Y���e���<|2iWcKZ#���E��	���^y�H��u�S���m�)ʖާepǱ�E�&
�{���x+�"��19C(UC{�^��u�]P�;9�;J�k�ޣ��Fo��p,���~ȢJSܷ|砤w���k{z��v67E�j������89M,�.x8�hY#�������0����6gPS;ˎ��7�2����9��zz�r�ݟ$Knc���>=� ��[��{+Z �ǡ�`0�6��'��;�g+O%LG*�n�މ�pG�oWQ���yap�H�s�[�!e�L�e�d8lg2��U͡D�I���i�g�h����E�A�����y�I^��^rZ0�8�}tN���n=�hdԭ��;p��"c�98Vd�v�y�t�m,�b����
AV1��oY�f�k.�o�[�M�y��]���00��|���U�^������_u�[���v4d���7�y�;��gu#6���:r9�����Z��u[ں�cIY~	uX)�`'�sVs��Z;[ ����C���|5�nᎺ����Qy�0,�1��ꁵ�~�m0��`u�`-�5��kU]M#q�t�Θ��M��E�/⡌���J|���|� Y�Gq�l��^�`�m��gW�J��	��܏�ր��4�߀z3�G9�Z��J���CaqT�]�+���7�]K\��iF���1@~�ı�����Qj��0r��dGL	����C>qJ���o@�IV�u\���֎�i8��0�`��ݻf@z���7��tM �v
�6�DN�����"Xjm���u�vpa�oI���Ʉ�^���Dl��o��@��l��uS��Ԍ���F�Wer�,K �U��䋁w�s]�ٗ2�66�Q��F������a;v'(��s	�X���:���P�&��M�s.�%�,�fnm;��Ld�4�sxN 3���^�oV\�6:{�k����iVW�W����l{������B��g��-baU�U}1D�;M�m�%��xwV�����ToBj����j�N�"�D	��ờ���ˁRG���R�a�tl����-��;a��*6�M'�x��ռ]��Q�bN����2Ǐ�k�����Ov_3�^fАx�Mr/W��Lv���KG�tOf��	n����]��E�Y��Tz]�U�>@#͹t�Gq�N�a��w]^�د��냇G�g��O��G�oRh,���۫�ʧyH����q�l�B�D��\Vh�@x��m�7p
�>קo6C)/�8�;<�	���Tl%�mj�/]�t�%Ht�pʴh�Hq�q͵��=��ʼ��Y�gO����m@�!��'^�:�j��^̲܇uE�����T�׵�k&ia���ٗ�6��W�|v��;���	���5�7ܒXD�3],߆ea����Z_���qK�a�\ﾩ��� H�
�)���2�]�z�$#�75�J쎺M��������S��}ǳ�3Wk�*w5\ﻷs#��f�ʫd�^]*n� K�������n?�<��?�D���g6�����2��"���5sZ�޹������x��z�s���2���Y�Vo���ne���@e՞{5"1LH�vvX-��@�1��� ��+l@Ꙟ�"F�0���{��ӎ��*�]w�"��&��@����T�d���@Z��w`]�Ǎ�n��"�.�*ؼk�W��K>��#�c�t.$ <��Y���A긐r��%�?C]�`#ב�.ee�g9��hy�{��c���7� �0�ǣ]_X�Q�����p�uV�����G�Z�oh��;��Ên�m��D�ߙ�6��wY�i ���)�dU �	�f;OY=]����wOg�ޫ;L�[o�.'�ã�9{���8j��c̸�[0ϣ+���
�aBz��V���5e�X���+�@Bf��WV^{�驐�5x�#���T�tl��55�^U����#���d{�oVE��{�{�͎�E�RY�Y����Qi/����&Ik;BѴ�&7m=��q��h�o���x�߈�37�v��h�.�4�/��[�n�ֹ�ls�A,���7%m�΋ၵ^�:ӺU�<uHr�WN٩Аl%&G��6���8���7����N"��PQ������ep �}�pa��u ��˥!����N���gZ�wM��@��!����T�Ř�|0f4"���%
��Tq��E�K	��8>D��f���ᷟ�u������N��4����&c��~S�[`�:����nSl|��cλ�&�U�u�w22�2;�rp��C,�.(ӲR�CZ>z�Y G����u�uk=�X�F��/�z�_�ya57@v�xHΧx[!���nl�ɬ��G�RFq��&7z+ 0*ˇ�M���>��R���uV��B�4�9�K��}�[�L�Z��	��>u���M������tO.���x|^3��˹�����4��9#7�	T�B��Er�aNNe�6�+t���l
�ڷ�+7�r�
��4յA��y�vC,=�"�t�p�3�0S�,೐��dO��Ty{�D��WK\�,A3Ӯ����Tqf7�{w���p`� �A�H7����)�<<>�9��R��9�wj����{zKL���Cgn
���<�N��g����.��-�O��+j˺��Ol��XA,ȑqP � ve�qw�[P�w`�$��ঌ�|���6���W���;���]����~k;:��w��zd�������OeSi�B�W�F�ⷸ�ݞ��CX̐׻$Rgj�w�>q�&ӹ�S�@�Ω�ut���as�ƌ�Z1�0���\��U�yO�~��F`�6�?[���l�7�[TVGC�sŽ+�D�WW_������7��yl�<������j#7<K�i�e��jj��:�*��X�������s�# ~N��D��Y�[�d��:w����`��l�K�W�0X-4�!~+���g��4�����k�)t�nf�5]Q�6�:�.���kֹ,�����f���d��JD���Ψ.�CT��j!�A��l_��4�Y�s�l�Se>��6eZ��T4W�{�����[ք�9����p�#Ȉ8ۖ��<CW_�B��c"�e�qW�˓0�Z��n����7�,=ȱ�3�鵋VK��WD:+���k��j���E��C��9�m2��:�[�'V��;�E~��!n� U3A4�F.�ꄶ�y�k.Ǚ! Kp�"ۛB2"gG4�h4g[�y�cK�Ε;:���GV�b}��e��WK� ѩ�*j�W�{�G�߼�d!��ɛ��Iy�i�vq5Nu���w��誦5@o]w8�01�7U��Y��E�r����6b�������g����F�:�ɱ�w����l�[��;�����״.�27�`�����Gr��?兾{_W�u��|�Fƈ���u�t�r[#sx�c����yN9��v�چ����B%cs��w�P�<�mY怈�Uug�+�Q���3���'�=�� �P֣��i�����٣�)n�<:�Z�_j2��zUB���n�}����!S�t'\V��Ç>U�u�)���+׭�yzX�%^G��*2�x����K'�'Ry�E�4J93�m�ym�:�)Мqm�$|v,�n�@��](vm��Gp�+�f��l.i��,Dq��TN�I�	���@�N�<S���-d4w���@f(�߾f~z���y���r�o�'�[s��-p�*��e<�o.�)�u�ʐ%���d�g��d����oWv��	�ͷ�f�~��6���4k��c��A+C��-������������7�,��Ɏ͛��-U�W�� �0˕��ٵi8�[j�Ҁ�k��>v��b^ �<V ��x�U����\�����[S��;�,���}z$\�r�<`����&�EV@嗉��հڹW��諧�:gvvdfm?bV��v�@=;. U𺩍U���;\fsh�WsP2�w�u֪�+��3}N���vPm�Saknb�c�H?f���f|+�O���y׳��]O�m�- �rI�1|�uګ��� �\wF:N��\�' mW�<��"*��ݨ5�u�".f��lo溛���w�x���,����42�i�a�O�Zˆ���s�2�f�C{��
�+�y^>�����m�]�0���覩άC79__�|���S��!��1}2�Sx�5uz����C ����-JZpb�iW=�;8�!�� ,H@�[����#��3�W�pݓVA9�ѵ�>��s�7 h�]�Ֆ���m�r�تm�V�y;[�ѧ���|쐒����^���fE]��`͡��@\v˽�J���D�U�s�/�7ߙ�y�C^�n����o'v��C_+E%�2-����,ˡ��roD����m�-C�X[8Z�p 4��q����6]~x1]�B�a\�!BZ��ػh���b�j��z�>kA���[^�w�6�S 67�g�P�\��m�-9ҩR$��D�����|�;��)��f�`m\6��.�R���ƅ䂲�6��㵦�d^#�LY�t)�#������vг8���;-e1��d����<�#d�+�{�_���w�����iIL�bH"�����H��D������27cǹ��JT�JQ^<�`�K$�$�E����"

$(,$B��"I$3^���$((�PX�vDCRB(*"EH��I$PY!"��E�$7����ZK��B����

B��bH()PPC5�5$Cʈ0��!BвPY$���(*B�
-"ҒA��Ȅ)-"�!I-,$I�ĐRZE

PY�ĊIiQ�T�AQAbE�%B�JJ	(*I(,I5��Aa%"�T�AbIKIhX���(�--D�����$�h��J���ZJ�Q*�)-"�(,D�ZU$Rд�!E�XE%��T
��Ȃ��"abO�������Oo��	��"�	 �j�������������{�D��������7�{����T������������������?�I$I7?�?�?�������D����d�$�H���\��*5c��3�2O�������$�$��~~��G��7�g�,)����'���8�4����#?�n?�+�����$�U�[M�F�K[3[[k�ՋTkfV�J�5�m�KkE[%l[c[%[Ime6�e��mi5������ڣ[%l���Y5�6�M��[3[%��k�-l�lkb�-�kd�YMlkd���kI��)[2�%�*ƶe�-�Ml�R��-l�[I��m�Ml�ض̭�l���ɭ��4��K[���&�5�j��d����5��ضƶm5�5d��V�Kl���l�٬�El�Y��U-e5e5�M�+f�5���[2�+f�J�R�2�2�kf�Kl��f�-e�+c[ٚٚ�U5���-����[-������l��Y����+e-�Zke5�6�M��Ml�T[c[���M��kk55QZ���5���m�ml�j�m�j��KBI-��BI-BD��Ȅ�@��Db�B�-IZ""�Ej�ɵZ�[ckY5�*�MZصd֩��-m3[ImF�3mV-�f�����Ċ�k�FK������ �KR	�"�$Z�A/�N#?�����o�-������$�G��s��>$�$�&�̏����O���w�f�'��#������Oȉ$�&��H��?����~������D�H�s�$�$��?�G��O�k�n���	�=���YI"I�,�?��)��]����f����'�I���n4��qIK�_���#�����"I"I����y�����?���ѮG��#�?����t1"I"I���,�O��$�$��y�y#"�?��bd�h�'���G���&��S���?��؉$�'����M.?�4����G���9��װ��O��B�A"O��<,j<�$$���{?����?�?������(+$�k.�� ��B �������3�ϩ ��Z����ժ��V�m���Il�1�ҭ-��[Y[[T�SI[X�f&��iV��m��������mRm����\Ym[,���5�L�ƑF�3m��	l�6��u.�IK\ЧG��=�i�,Մ�[`��[F�h�hڶ[f�UfbԱKZ��f�e1�dh�-�l�A�jf�V���/}��LKe.   9�{(��RcN���5�GiWu]v��(l6�鮝��9����ж�i��nRv���dٓe
��g����m�Ǿ�� ��m݀ ���m� ��w]ѡI�] #�l�VYd�Ţ��� O �� )ن�;vq��s�uh���[��`Wu������;�j�����6sx 8=���u����]���t4w`�.Q`�� �������)\��֬l֚�m�x ��ʹ�۷��l�hj�r�k��B�vqB�4�;���aE�[sV�6�H�cVd�  ���.�2j:�k�Ce�F���n�hU�qݖ��I�
�\ܪ��Ui�w+qU��eH�fd�J�n ⪽i*��©UT�iUT�����UBN��U*�.T�w\�ܶ��R���UU*\mT��Yñ��-����7o wQ��US��P�5S�E*���EP&wT*�u�UmPl������W;uUA!�n��4 �%�������� s��Ou�J��Ne�*��T�iU7l�
�SmUUZ7[�R��r�N��@TwwT�銰wYj�F(��^ =Ӫ�l<�Ԫ�T�a�S�΢����nj�U��rC��J��Wrݭ%J�k�R���  P ���)  * "`1)*� �     �{#R�!0i�`& �	�"��	J�� d� 	��&1j��@��(�M0����CAA4 f��h&��ɑ���6��I�D���������  ��6��˫�+n���ye���Iz^�ҙ�r�o�[�EL�
%���'#�@�U�j���UmZ�����*ֶ�,�����?B����~2����~��BD3kU�Ͷն����~�kmm�
ךm{`���k[[�m��AHDA]Ъ� b��)�k5^������ ���\��2)����[�Jq��tyOd��^�H힇�
Ebb�Z�*V��Ҩ��r~d����"S��R2�l�?T +�0�o��K	������dP��E��"%(Ð�D0E(����*8�$��o�4�m�R�-����i�-D\%�
iB�0)?H$��bE�D M�[�R?�f ��Qp% JB���M�c����Ut���V%Y\�8�,X��X�Q��B^뒋���\���Q��ҶiG�c��՚(Q�tte�˱�I�,#2F���$*4[ҁ���L4X4�.�҆L�6/�,Ҕ����G0�Y�\%
Jy��?�aJ�"�BUee�e];dZ�H���٭��Y<K�YZ�j
���b:Yl�u��,Zt�Dj��c���w?sɶ���azC�{�UܬX���T�*Pw�3m:%c��Ve�����%� 6�<���V[r��h��8�ma �C�.֍��Y.�!x�CP�X-щʳ��+��S#�1=8�ʭ�tD�4Ƶ�#pЀ��N�Eu�3KE,�qE+ h:�:�c/u�yd��꽥�J�k/V���[;NaK��M��a4v�ӆ�n�"�CV�˨�H˒V�b۬X�6�P^F�m E.�wY��P:,n�n�6ݴi���Vh��E<2�d�it��yV�["���E�4S'�:��i��#-8+#�؎��@���X���0�/d�aխ�Fokk m�ŷ��ik������V�6�"��`�ٱ�QʫաyX^�3���#�֣���9�ju4�i�[W�7-�P��a�Z��j�}[(�R�F���l�YIksCn��)�h�v)�m[7�*^)��0,x��\�vN��!�N6�+-"��7{�&6�a���)��X��;m��D �gp.S���)|4W�B]���M�]kZ��\S4�'�gA�HT��;�+ʵ@o�jF/���׺��%8-�;�͗�4il,�U���2��oN�{y6������uv�X�K�c��\WJ5�#��a`2�H��Yh�7?!���v�jE��c��\:�W�Fɏ#��d���c�P���(��(��C�i�mٕ��L�ͻ�~Z�-��Y�	�m��h����U��0�e&'�.���N�Ab6��ͤ�R��Q�Jf��X��3i h���Uba�{��mð�RFm��v���p�VU\�)4Щ���e�zn���3v+�Sf;�!4���1)}CN�p�iҒ���	��D�/FUUZ�&�u�@�0+�f1�-�6д��╩j`��̼e���7Z��a�5x�5x-��jk{�i�n5M��o��.9R�HuY��ƅE1A��(��j�	Cz����-"�V�n�"�h�8�я/�� �T5�����[I��J�h��ڙ�*PD2�n�t���)c�5�UM��0�z�%�a���`РiXv��LԱ��;�R#a��.�c	��c4�f�7g][[L��h2�ml����*��3%#6��e�⢪e��(��1K�=�cqDU�e�D�ˤ�����G��`��F���4���V�g̬ÊJ�V��C@���i�Y�&`Fm��`�����oR�fVFW�\��$\Ū�V��;"��Iɚ���H�q��e�KN��ކ�� s&��\ON8���U�9.S3V���t�x��n�oe={pYW����T�
�˹��ŕ� �L(Ez��92fk�q�iKu�5ݬ{����YV.�Z@
͸^$Vf�G&�!����n�#����7O7�������g6�Ym;q�E�"��)�.���b��aE�{��f��%aC*�u�M�Xa�nSg
��:�˔���Q��U�6&S���[� zɤ���=�3P��n�o�$�,���V�l�� ��^�^��!QE���#N#Z±6ڌ]��o�{&��q��SVm�-"�<��4�ݨ�p��k�nL���ּT��D��.ث�]��iC#D�m�O/cYD�*�;x̥�v�'6R���+cJt�@74Tf�c"��a��ܛB���U�f[v����ċ"�h��u�r�6�%��IH�W�3^�4U�@��n��J�*T�k25.�,��jrV�$ֺ��u��Q)�VLZ�Ce�8��]J-Y��,�Z(K0q���0��]���7���� �;n3R�Ԫ�ۆ��� YE��ni�KA��z'u(�;�1ME�Ɍ�T'��̐T^ͱ2��6��tK�0Uf!N��F���
x[���tt%W_�Ǣ֩0c[��jځ��*�͠�N���9EiӪ�f0�e0TB�sq�b�A�]F�[�����E�M�Ѵ�a���Ca7�<8�mUn�U���CbJ�!)ln*�/��%´^�X�e�Y���Zn�q��H�ɏ~��]Z[uj\`2�ݹ���k.�w7ef�;-��$Z��k#����%,�aZ�M�Pz�aǢ��cC�mV�T��.5��vFNmJ<_0���+y_J_LǛ([,ͥ%`cm�F��6�$ܠ�q�w���,��˔9%[0ǥ��TA��y{G ��\�����wn��aI�̕���2��w/���������׀�ө[z
�۳�bd�L�C�V�K8m�m�TS��޵G))��̹���]�\�i���9Y����E�w/P�$�`�X� �#�/~x�k"�p�%�,��co2:cY�Y�4�3%<ʄ�W	{k ���cYxH
�j
d���H"&�Mf��1f�*��ǵh��[Ʈ�X�*�i��cL���XĐ��+!�[�&��m�g��r30Ӌ�ڏZq'6c ����z��hU��wa�Y�-ꗘ�XûC�F��
����N�u�4`TV&�%e=��αi(�uA�.%�n��D8�����v�V;� ��/	/e��l�HaY�ָ2�Ј��u�=����t���^����+La°�n݈܅��{"��Q�3?J�๯M���PzNj��Lӓ(��9��E�w �K�=�ɘ�G6�1���z� �(K�kHdM�oi�	I�F�ր�-�+tM6��齊�K.�XŊ:y�B���ɹ�ch�I�#�b�W&���#�V�&P�d����2�j�%�˷���-4�Nb1.n�ʺ��#�39���3v�j4��N��Y�m����R�q�[��-�7	 6];Ɯ;xji������ҟA��#E囟^�k8���
G�.5��q�e�:. ���
��ń��-Zy/n����	&V�	�E��W�!X�^�d0�L��f��LoMkq�D�N�lb�T-+;.��ཊ1�!��(]3Z�Rj�i�Z۰F1�t	ّЛN�^�ܫJ�S����wS	cb.�W���[l���DX� 	���D����tF��v*���]\�7%����FT��,�Ҩmn�4b9Ykf���:7Q˚�)m�9�ȕ�I"VMHU�n�Ӎ=�o[�F!��ӂ;�/
y���鵐+5&�]`����)f����Ʉ�f����
a�՘���Ve�4D���`�=M�F��L�23��<J�4��$���p��G��C�&���d(.��� �%ym͈��],�Q��Wi屗z5cp\�)
+a͚bl�dK�oHٛp�u���f���(��4��츖�4���Ln�j^��ɂU��`]�u���ԩ��L������c�:�7wS)�����M�M��N:N��I���[��ϮS z��I�>9G[��a�ņ�w��FEf�Z�n��*+)қKp�n*B0)��<7����X�`�;2��� �+���q3;��tPyE��f�$ ��5[��bf��;v�+c��"�Ph�&���q0�M�9��
��]jf�֔ Sf*y������3.����)K4�{��X��w�`
��4>�--��v�fMŚ�Evi�uj��q��K%ǔ2�{v�m$\�X��
�1�-!�f����jR�H�&'��D�l�2����R�-�D��4��[�dr���8!�b�azɕj�`!k"�-���0�6��GiK#t6�(�3㼚�鷑C#�a��[�ur�w������1j�V�9�zT1��Sy����.��d4�P�6�"�%ᅙje���!j�b"`.����.k��T��0N3YU����C1#�����$�Pe�[u`���܃� ����+О �ٕ*jfc�6�enQ��W��1�Wt1���\��`���Qv�%[�PZz@�pMb�y��F;9B�X��m��*�Y{u�P���y{+v'1M�/vn�1�5j�l[tKs@5.E{��%Ɲ[1F�711W���&�ɥ�2�+Vv�Y*`8f��5T�r*3n�k;51sQ��F1�+X(����׊�3�g(q�4긍Kg.ձ�i�0fG��q����s,�{rhWv��-��?������w��i�v�͉�5�$�7�t[CqS  ���xn�M,��""V��q���47E�[>L,�B���F����w��A���c�pAY ���h���tu¬Z�eҭ��"�,�cU2 .#����X��/M鷒�D�FT�z��n�q��H/(᭘.7��<5�����e�b��(�r+�"�e�*����C��NR��@H՝�ǒ�V{Qciӧ��1Z���[j��aJ�l79h�*�Ң�C�<�,K���f,"��ɺ��o>��j �ͰR����'q][�	��:�$��˳X�yQ"J��!*�I؍S�*�h��L�=��#�5ա���&&t���b��]�:g$ 5�A����� ���3��e�A�đ0�E�,�N�'`��M��e�@�!2HAQ!L�Q�2�_�P��(I��H, �P�̅�a���2�DC H��d�q"�d0p6!�\%Jr9��`��0��
F��"e�D!���������g�I����� ��?�4e.�[��h��*�����ݷpwZ�$1�T�P�f��gv]Ϲ�t��/騳�[��m5L��С;	Ω���(��{_.:��[k�u(R��e��moU����:�P��6�5;�����u�ծ�g9u�ηٜ7���Kn��y�p�#]����Y�y�ćP�}���v� �Zy�\+1�lUf���v�ƺ�ƥӑ�y���Ya1�.��a��RϪue��&ч�&d�%�
9S���&jt����x�"��]�s�ocW[i��H^MFe)���n�}3R*�^G�	�R��y�ǁ�ۼ�]߽���|���*�]�FX���1��%�f2�ַ���J'J39��>�ܹ�ب��w���� ��zw%�U��4"8����w�I�&�U���xu{��v���x��0�w��EV��³�k�|�c���:���,�Ɖ�핸�#���/�y�pt{d2��P3��WY�u�j����a9և^EC�9&�\�i��3��x�J��@����eh�p������ �&bT+������Z3�sj%zB�T6HS:��0yE[u���B=�\��t�x9�1��}{!�l�K�]�%�bܝ��zBu�7�$�\ˤMƳ��Uoms�6�i%l��\@%�����lw��b:�������{gmu2�D,}&�.mS�i९�A�G���<7�.Mrj�����ηK�w�|H^�;L{�W���{�&�,�w�Ԣ=�T:�D��$�x+zgd�q�eб��`�6����fvaÍ\�)V]�l澧����1����-�8AҸe\�W"�sFu���7�1����j5��䁣˫?T�`苹�x�ܳj�՚s���q��I�]f�:_=*FM��f�Š����v�P��*�s��͚A��T���5�N�APpo^�D�|��g;0���=��pPWR�3���wR�����(�gvݩf�:��&�:ÝG�Ԙk�jM����	N��R��eX�Ki9���w^� �jWo�7^��?�S�Ÿ�z�����#�9�NkЪy�V���W����a���h��]�*�@.A���bBv�7��3rP��f!��ڑoZb�De�[��MJ&.ya5��*�����
^J��פq�+�=K�{}d�ͭ��\���5��;�������vbKgR6��v�(c�AV���v�Bh�l+L����)���H��ٴ�O}�$���K��9�n��X7���O&<+�Dme���-���\j��ΰu]f2r��E-�][jf���S��E^�rWk����R�]+�BI�X֎�d�߸Ĭ^e&���#^w7+lq��R��5��S-��ӠN�O�+o
�:�4J������,� 2`���5�*��4��R�R��\]�	VoNL�t+gh��s�՝#z 3S�+��i�ru�d��,l"��!����M��;ή+o�;����y�O#O��_j֥�0���M�X2�ųn�����W���S��HR5�r�י]���ݒ(b�%�k�=m*�4_S�	ŵwt��\�˴��;9�VSy����Agpx1��;o�V1�V$�F�n�#X��]��\�Ym3�v�͞9nA�;��0�^cS�7�8�)q����eNJ[��Yc{m9����^R=,R�����w���2Ռ�yz�ηW@�AsGA�=��6;��˨Un\9�ôhI"�͈���l��V��-�1PS��T���2�>�6�;Wbճ�'6o.:�חgA�nFq���^荊殣eW-���=L�>-"Oj�:�ڧlZ~u:�]8}ڒ���c��O 9��ҳ�,��l*�%�4r��Z����ߵ�VӖH_u�:��qv^l�JR�8nF�����Ev���z$&���(��Lb��8�e*Jnjl��>�y[ݺ�;��zC���v2Ts���c���[BT��#�":w�w��P�ܑ���+�f�ZΠ[r�֫kæ��7l]�t*�|��5��1�CjE#�z<iL%tw���R�ݺ�Js������wJt���m{��ofa��N[��(�,�x�\*G�^sݹ2�䡮^"�K�/{�#\M*$oA}g�5�\�ѻ��޵e}@��j|�鄈,-�smf��v���k��ۧ��w��Q;T�՝�ֆ�٧Wi9N��x��;I��� ��E�5����{�v��2�fv�R��t��v����y���o7Ϩ�ٳdp* 7�l��v�%I{�%q� j(5D�oދݘ{��u[��
�<ħc����0�WܕK;��l�jS-�ԉ���]
̓�1R݈��2���J���Zɂ8�h���H^�ʼҬō=i�yڂW�fA7f]��`v��s�,PװWVT��W��;:M�c�Qw|���t�d�N޹Kj����Y���v�V�ܖ�eE�T���}Aif̈G�#�G���.�&��{10��Rw�@�k�˜�Yb�H�^Z$s�7{y`�����ѱ��ON|�e-YA'}M��C]d�tX����i�4\����|��o��d�l���v��2��f�9S�����{�GKTO7Q�v�u.l��s	�� �MӬ��1Jz�]�6�lv7)����W$�Rk0m���%�0U����Ss�����e��)t25��չ��v�]��E��Z��.��:�DZvN=�,�-E�8
�3�C�عڙa&lg]������۝w�X"�L\G_s�"��R�:�㧗]�N��[W��GoQ`��ZDXڠ�;�^�}0��ءK��K�r�T1Z[D>�!{6Lp]
��Y�ܩ2#E�ta꾓�2�%'|(w3Zn��^��\�Q̰�����lg�SO�1��.�j���0�꙰^��]]ݴ��W�o�`�x������Z���Â��m^�q�EF��i��g�k4�o�ɄSn�!,7���feadj|�v��wf��T�Ҳ�<�*�v�:��6�.aP}�,jt��)�L�\����\��V9����[Yì�[Y�Ѥo6�~���:8����"%�9�T����xV��w»�e��f5��;��V�����������jVA[��1e��kێ$c�
��:������(2j�[ґP��?;uz�#mxZ���T����gaE�a9�<=;�-�/�b:�g�%m�7I�ۏ��5Õ(x�љxq�<.�0����K�u�o{2ciEN��[���&���ޅZ����X��5�fۣ����{�Zb��o��]�9��dJ�^��λ�j�ܛqj�-˯wb���Y�m��
�i�����n��;{���s��L䩨M���ݼ6�3,7�'�e˕�5�NK����`�k�{H[�� �|H��k�&���sn�S��Em�W`1׃�Z��t��cҸ�q�:����2Œ�˔�bJ�LV���o�hj=wy5]<�ֵ�IQ���qrU�@�e�q�by���8S������a��Fzvg��GZ%���������[!g�	h(�X�'K傢#�\�}�r��S/�M�{KTl��Mr�N�d*9����9����U�	ΐh��.�i��"}W2�%R��!�W���}�X*�٧6:��#���V�r�qx�j��uP��8_b�RmvbW�)���|Aب.#�b�hM���ʲ�i��*1�m�z&��֔VO�o6]�i�U�W=;�¶��a��-���Yt�3�7q�n�G���	a�����%f7����C������1�7��W��o��"���I���ȶEpˌ�~�F ���]hے�����Gk���{���R� ΂R�\cM��:�c�MǪ���(fvm*貭�hK�ݮ�_��8�X�P:�:��=�A!�+zZ���]Ӹ�ǋXW���]j��ٴ�v�0�n�| ��a�����q����L4��hb.:�Y�sR���;d������=���f�K�ՙC��Ueq��mHl�y�7��+Vf����Dͮ���N�cJ�f�v����7\.M�ヰ(t�ƕ[�c(���]<�+�3(�l�!��ܾ�B��0aT �u����:����Nh8�q�ͻ��˰�f���ʏ=�c�l/���&p2��\>79���_nqb�o ��KJ�����O�u�O�]&����^]zL1'�$�F�%���I$�I$�I$�I$�I$��vt��;z�/@��om�w)���{�E���S���+*�-ZKv�7���$�I$�I8@��d�@$��U�$�I$�I$�I$�ID�I%I$�I$�I$�I$�I$�I$�wL��Y��A��.�e�Y���I��o]`�2�.�-.v��-QSgI&���I$�I9��I;����y�KMM��h���7���'ӫ�n�N�گ�r��m��"�0^,�3��ۣ���'SDU5�1XY��	ج�I#@:@k���ye���-N2��rj̈�'	$f�Nu-\�7��Ӂ�K��ڵ�]oGo�TT#@��&�uΒi�ij�iX��"+9R��R�L����)�$�w��ko[��B�ݝ�WX��yb���h�*y�"����r���D��QM�ͭ-Ds�g%�$ݴ�=�S�]).��W�d�զ�P�f�x�Y�����Ce���!��v��6᫙dZL|>�S�t��D�jr��;��a�j�wy-H.��"J��w+�o�{��c�� *��1Z*`���u*"�v�9�y��b����el�݌S8���r�Y�S,eLJ]V���!�l�̊J�6Pd� 9�p��!ǅ0?Jv�q�˱��RC��S���r��U����=՘�p�{��>vy�%����Ct+�2���e+o+�݁�&������l-�U���-�X����%�ã2��Ci����,�[����gP��Ϩ�8wg
�A�v��eKK�g=,��\�n)m�[{iD�]���\8�:�$���7#�2�=lPԬ�`B��יO(�܉͸ �X�����>J����CX������Y���۬���QgZ�WP��0�f)}�(%�m����fS���SkE�n��2������mH5B���XWY��쮇/�Ã��v���*��H&��=�d��x�4]�ґ�J[!M�^O�V_3��gR��Cr����~�ӯ�ȯ�e��C���q���/,����\���a�ff`z�]�r۾���F`��K�I�O1�O�R��]<a���V{p-�˴��]��f�D�\���$:>.#tQ՘��.��;:��
]��:��#���L40�}���=�	
k6z�S=`IE��*��i&����n�+��P��zX@���mB&�R�R�:
b���lܡ:�*r�
ꓴ���M �+����PR���ܥ�\e�b\
���wb���]�-t�C��n7\�Z��^θm>�lnF�Vgv�Y]}	KM�LM}u�n�a9fe3�N$�ꖶTwE'��2[����A}�U2��k/�b�D�݊��[��n�ŝ[
6�"C��0��a8��v�μ���5:��W�{�;�b�+�R��c��[���秬�es���������,�S���R��}}&Ü�}ڒ�69VN�;%�+Qc켔�!��n�}�W��0qc�Vº-;�-H�m�d��g��5���Ne"gd����#GX�K��*@oqF�t�s� S����L}|��voV=<�-�m�OMp�\�fP�euf֌�|՝��ky���kj��B�I�����Mp�\ ��}�*t�d�(Ѝ3r�K�+<�/���]����W��u��;����y-���G�d�/�m�Ԫ+�h�8l��(
n�RǍ���r�A2~#�sJ;�L��{��h$�D�Ko���&K��fu\�k���t�4B���ռ�U�w��
}�`2�lk`�xWpc:Ն�]ώZ�<����\�$s�f�<����p__c&�|���C�L��f�=�1��g�.�Ѯf���c۸-����dcwX
X����W�����L�7>�i[K]��VmA,}�����q��1�/'RH�R�Ζ�}kVIu�'�m�0��Br���ț0�!� �LS���&�j�2�����;���'M��ֽX�ڝ��
�u�B5�z�.[J'oe]��L^Dw{Yʾ���������Z�Ŏ���H��p㣮��n�<�K�����@�.fΜ���;��Be�UEW���U�˯>Wg��c���lK���i���.��37Y�v\�����\��u��H��!H��i�Gxf'�G�L�S��w�5S�9f�b�)r�(ݦ�Cw�ղ���0�6k�̻�Do	+��Q}���:"�a�#�\�D�r�7X�w��sC�i5j���Ika3���Ի�5I�.5�7=l-;GSRf�h�A��� ����w��X�L�����6�H�x��Ƕ����#���ݺ讷���*����+:H3];"q�>q4��-7Y����X㒲K�c���/X��z[)��c�,�渊��GnMT�6�<�s�M�:�n
�E�a�{k�@��r�c�:�gPc�Pk���˓V1-��8�dTeV1�L�w��p���֍�J��m$ɷ�C��U�2�71u)�|s`˂����p>���v%�Z���{$������wftf1�y��R��N}�כ�pծ�=KF0C��kWeX�ī�mN��`yz�;��A��kzWKmu��J��N>��s0]���Iq���.��pu0�Tݬ�P�z���LS5��B��#T��W>��}j���4�3�$/������q��]��0,F��O;��H�ya��͚�"'K��V����V6>K���8V5Y����Э��k	��e�|�'�[}�c�Ԓ��`�P�
����N/�L��J��.���@���Kjo�X-9ہQ�sX�u��כ���(��s�M��~�;h�m�]��k�G�9��"�ʹx	6,����Y;��&��!AεX9,mm�Qq�9&���D�����4~euS�σi�)�7-d�-�w0DM�@�Dw��Q�.~��l����	��+
{�H�t��#�@�
�M*^�U;ǝ5�9��{�D�h�mgo(i�S�C��t.��{�h���L��I�T�gh�1
O^݋���l/݋5p��J����[O�]�n�}����f���\ȤuUK��W[�D�f�T�F�S�-�I�����AῪ�9_"U�L�Qʿ���p��CS�� i���s���wi#f���_k}��T |9�9�}D�<�۩P�|��m��Ԑ���wEv���9X�T���5_<ۭS��T-��`v�$]:��7�-{B��W;jEglx(���MU7�˲�/rJ�������S�aZ�N{���x�����o��:�n��D��Ox�2� �V����c�(; �X��
�~/SN?ߊW���r� �!��J����G<��+��l��U{��2�<��ZO:U�������닲u����\�+��)d�Wk��uf�x̾�ZɇR����f�t�.uV�&[w�T9K�����;)|�ٍQa�t���6[���-������u�}cso�j[��ܢ�_��8\�l�>�B��VW<��c��Q1�@��QaXr�q@J�vu�Wχ&R�RCK���wu���u�V�T��?`��t�G��~��U������}ǲSx�T|~�4��e򯞁�nTz<83>������Q[e4ph���"d~�T�#��c�h��[k(+�:+�B��;��)�/���z�x��v�vf����n?e��'��屭:ݬ��+����j��]�E�n&�Ϝ���螺�����M�o~��]Z��S��-�URSO�������"u��+�2��4��@���ӣZb&��Xک��Y�p�F�ƭ|H�Xܖj�}�y�6}v*��BA@���-*����-)PB��x��P�AA�+�:�cU* �Z/V�U��ګ��umF����_ek�B1!]�*1����}��u]���
��F[�*��ݯ��
m��U�
}��qIv���E���Uz������x��e�
�L��f�%vRB�/��ٓ����$��2�ȕ��d�ۿ�V��Y��n�g�i큛X*�r)S[r��������Y!3U���f�ѯ.%��0�SC��LgR!_\մ�q7� ��as��f�o/2��!�[�`2�0`Y`*?a�x�cES�oP��I�n��QO!aW�f�{w҅-a���v��J>Qe�_�-��Xs�w�϶���Z�s��<�N���[1����()��7��7����]v$�%<��N]�ұ�|����-�2����a9�B\(k�'2���r�(a�Sw�����
��21O���� k�C��H�k���ء_R�M�q)�Ŭ�Rw^mr)gV���X5���Ok{*�X��Z�Tt^���4���P�x���hSs��J�|���u�t�l�l����*��Зݴ��K��q]̮�ܤL���K�c����8�v�ߚ鮶�ȹSΪژ�Jm��3{�t�.����&&Un�k ڮ��;����'���Zw��sv�yY)g`ph)�2e�2qf3���4�,�Q aR�*�U�54ְ��Jm�|��7]4��g[�MŜY�n��cs���|n���-#�3�8���T�3���N��8��^<��G��q�c)���Z�ˣ����Yy��r�Z��-��M�z8_0 
H�5�;0M+�t����])B��,Hř]��]K��]|5d��H�u��S�s�*+��E�}�k�hZ����:-�l	���3��6`��6�Lyfn\3�K�/f������l�W�4!��!���飀�7�P�Ɋ�9��r|^��H�t�݌mo]��/���@�[�yv£z���O�f,����t9|�䊝N��U9i��>:�9ɹ���;�G:hG��v���ޚ�ur칙4s�1�ݵL��H �̕�Q]<D�z��:�E��R�;ٽ�5��V�"#�c�P_7}��:>��G��W��H�)\l������)�(�
m�f[TX��S�й[��s��� C+VU�j9ϻlr�̓v2.�(V}m����(�U���*0�8�
��T�o�cX)��ս��FAW�x�o� ����a���I+\�{��5�Z�m�U��M�[�M�|���L���`�K��;���o�U�����]��5S��G����u�E =sU͔`�켡:�}6��7���T�<QP�c���5�{M�n�����]����zۊ�2�yխSRνyO,�{ݡ)��j�.q���Q���#L{��K���!�K�Zɷv7ˬ�RQn�&
�eB�5ީZp7��}i�1�������FjWC �ql���<m�df o��֍�WD�Y�s泳1:���]�B &�f=��e�p��[ӝ��n���������m�HɅ���Wm�k�����- ��I��FC%I@� ._�I7���n�"@���U�j�����M�Aq ��B"#`�R�h6�@�C� �ߴ�&��N�g#�6��X��6`�+�G�Am��f
���^� �k-k����`xFbʐW%Q�&6�`�h�wŷ�
L��>J�0:�������AZr�Y�W^â�f��am]WZZ�7�!yCv��̂&n�Gfv��ꔕ\{�͍��]j�
Ka�����0�\�;�R��nt�z��q�ڢ!u^��s ����CD��ow�Vz���M�2���쩁>=�f+��0�N��WQGF\m�h!޹(⼆T���ii�q�T,�d�4���)��t�ǂ�	�c��p��N�֝&���.���z��e��y�>}�������ˆ�x�EH|^^�-L�Huk��ꉜ̩q�e���q�Rw)��8��ϻ��1�>w��|�{��������|U�Z���6��\��\�b��\�v�mz'���t��<�x�n��/�m�}�>:��Z���ս^=������k�o7�[s��[�x�{[٩�|�睫�:��|������ɾ�����0	I,�\ǯ|���I�/��ǝ�;��c�)����J2����;x��%_��K{ݟ;_�uӻ����Q�9}W|�n�)65]ݱ����X�7wQh�cQI��O��.�Rm%�\ە%F��ۘ�˸�W�nhM&��^�rlR�%���\׉����>�r�yۚ>�ğ:��^�R�n�պZ���)$��:��Y-2�nW.��f��b�O]D�PIo��̾=��5;��u9�K<�κ6~�׾�}v����0IFE�n���l�w.�ܺnq�9u�|xyܛ�����ě�;~���_�;}Q_<Ux��G-�;^1x��ޯ2��wh4�V�e�6�F�)/���|��̮�(�V���g��/N+�z�ɽ֨���[���ߤ(�Һ$�U*��V�b��}+�U\ce�m[����e����)�&��@K����{�?4�)vsJ���c�y5c�6��t��J<@>�����o?�����y���.�8{������
�=bCZ��z�W��y��C<d8�w`�׺����|aČ�x���~Z�剺����t�NyJ$2��8�e�z�w�93�{�Ra)��}�e-���$�4j�`��\2�j�G	���T�kvz!�C񂐯�+��ޥ�/��I�`�cҺx�c�]�'ߠ����y�1^��;��s�D���;ɫ�r9m��r����#�ZgO�2r�<�y�-_�&eܢ�	�ܨ񣻎ρ��a����:q5�h㰛���vF��ʣPg�;��\:�f#[�~�6��c#�We��u��6_���J�l>��3���wf�5��r��We�]o2����u�GJf�hv��_b�.��]7���G��)���L�m<$��r��q=ޮiKo�W|��.�ř���c
Bj^�Q�/�R���6~>�=�5Ҽhyv]��(�iI�j�t��
�K�ب�!�::hM|`���g���e�Oٱ�z�g�i�`�m�y��%O����1�<����E��\��mێW��2��4�&
wW��̫�E�h��
ǋ����脲�yا����/��?0R���>{�Hq�_��8�l%�6}Rڶ�XJ����q��4�Q2"6���`Cb��o �3��]ؽ�	���^nv�.��s���9���0�KAc��y��@>z`,���NYfu�{{H|�����KMy(_�fw�G�ZB��	c���Pɒ��u~�錖(-�)�Wh9=�ʪ��}�T�;S3L��ҭC5%���8�dL�5�G�1KE��/G1��CޠJ����q	ei�+���og��<\�x����g!�w �iz���-\]yT�7�Ն��C7���
{c�W!|��Ok�̌�:������2�]���Ӝ:������"�Ύ�L�s�����9����&2S����-y76�S�)0b��Bb�����IM	>@7X�v�[zZ�E��M2gg��Ff��rVB��B�KY�A�L[���;��O
#3	$�X�)���W��`��Q�{*�x�,\��y�ƦJ��_<��^f��s�y��)�b]5/j�7ɽBRb�Z�%ܯm]
k�O-[�B�w͗�����M�eX�yM��R�
Z��Z��h7CA��(s3�GW��G��n���+�l-��?|�\��}���2/\G'�W��T�s*��_(���5�����e��}'��*�W.����%���@5J�{4��V����fꄎe�Υ���z�ݸ,��oI ��T��Ġ��+j`&w253.�|ʐ靦�^7ǔ�X�o_ױ��{�XQHkf?���6���RG��vv��u$\�:vW�kMΫ��6x��*
]�|3�rЛ�I��w�.�[�����&�/��������^�F����+�?=�/)�=�.�/9��N_�Pb?!�JB`L���;A`\နYm!��l�ck�_x��H���b�d?W��O>�J1�]ii�il�x@��@ěr�O)z�����r�,�|{g��(Y9�i�) �zc&����X5Af6$�΀gϜ�Z/L�fz������HQ�p��
mւ�M��p���o6�-��ŇX�&d���P����L��5r���7����{ֺZׂ�l��Q�s�;���4_�Erb���Nȥ�H�N��.��؛���e��})���fYq�ξ��E� �i5�K�r�nm`�$��4oc�w�3�}7(/l|�5�5���T���ޛ�K�ޝ��t�������vv�y:��R���3Xq����T�����r��iƢ$,d5)h"HVۘU�:p����L2G(��dh��S��qM�)g����kyg������wsRQS;�����6�X���ZA;=Ƽ3b7L�j��ڙ�ˑ��Tۇc���������T}m�k�e���KjbŰ�I,e�`�gֆ$�zU�mE�ǈ�4XBhP���x�lh��thSі`ӈJSb7.a8IAF�n�)��b3a�M�Θ|�i��<��=x���s'RW!���Ρ�r�2Ι�o����^42ΰ�s���&���7�Z↰��x��ђ풌$g)j.��y�&�\x��8>��G��i:��MNV����84%�����u-�M(��A�5��+���0��+ݴzo����τ�ڞ���K(��"�Qа�O��S�*c�[j�o�U��O�p��� ��D��4�B��q�T�Y�r�m��MLcg,�V�LM�9}�S�L)q��پ�1��>O�=���,��/ݮty9�w��>f�἞��[s޽����){� �s������^�^��W]J"O=]��գ���:f�����t�n���r;��m��(%0IP+I��6u�� W��4*q��zq)9I���W���T�.�d�t/���;;#��a�O	�R�]�����=Y٢M"�@:�U5v�?9k��A��o$��Y�a�\#���r��AR�Ns�w��shĮv��G�nb&��O��Ͳ%��e'&:�lh�L"ȟ9�^XY�X�V�Vf���B"��N�+���\݋k�j�A�)�q���J�l��k7�������4P8�l<x.�aj�Z���B�:�����_�R�v��Dv�3˻���s��Kԛm]N-J�U��M=l鸹��,�KZ=��51JL�w�;V��4�쿊,Y������y��Ԟ��g���Y庇���u3\�jG�M9M���m�M0f��^�ԎD��]H9~y���*�t�}8Bk���X��d�v�Ȅ6� ��N���^��-}�YMU���F�wo?(�5��=�*�?e"ξ���gu_��Ʈri�5��.p$w��;���(-�Cxx��{�azd
ϐ,kr�6ԡF��|v��E�T'�62��Kt�n_X�uW[ȝ�
M�l]�k���(��\�p�°��#yܾ/f�v������J�w\��o�i�0��}�����T�])=�*C�J��4�F�L׋�M�vR �k�-��P��A�Z9;Z�G���sWf'�9/�d�� ���3@��DNFb�*g!�P��^�T�ޱ=�x�6�������Ɨen#W�v}�FG��#������)�����ϙ�z�L�n�<'��lM�S\��x��ũkKM:�PBH{|,�|Uu��\[����}<}���w#t�>�ipeܖ%�$L�N�fV�Y�E������fM�iD�@�ak�B���4�����k�����l-�e�Z�k�u�^�)�j�j{ݫ3��7y��_�{�S�d��kYsC�'˅�n�u0�2��+�uf�f��ڕD0r�-M��� �sO@8,��������|m����wa�����q���j��kB
ղ�M�ɳ�EVTA�jAL��Ll���^*��dވuhc<��֕$�/S���JԱ�4��E@�q\/��Y켿w{���nl���Kj-Crh�鼤�\3�o���FCP?S��5����{k�+g����k��#U�t�s}�?��moST֮ɸ>P�}�3Y�?3k�Ζ�y����N�«o��~���.�{^��čd����c��Ay
�>{m���2�7z5����4�/��1�p���u2�Q�FC����AĒ���d&�PkhӪ�B�^��6֖Y��o�o%$��Y�"Oo�"-�����BZ����uv���Z5c�X򄢻38�Q���7��[R��_oc�<�07�PǛ�����QN�0qJ�\���Y�J�2��]�,"��k{�ך%��` ��`4Ķ�jE��e�͙%�Aݿl�CάK	/�����Zk.��&��C]-��3q�wL�f tjѕw�qE@܇ ��(����$���q�=�h[5�S��,�ʀ�d���9�)����I&f�yeHʹ�qe�Oz�	�ÝB��H;� �cW�'-��K�	��QlZZ��hS[n��p��l�@�KLXqt02!��g!��cWt/g�7\RM��e�i������2��~%�ӛ��3���u.���0>.�<��W�H|d�rq]!<���ݚ�seo_�$��yS�k)��V�=�:u��jⰚRbfCfv5�6S��������
|?x�-���TƟ]ꂀ\�M��o��l�0��k�9d�lb;�������`l苶)�Z^P�7�2Ī\B�H��73W���2�ۭO��x�̷{0�+A�×s >�6� F�:�.�u�����SR�
Q�B�>��Q�{636�-�l����u���e>�vl(�Ju���]:��(��8�f���
94���9��xn��c�ұ�yJ�͵����K-<�뜭uZ{�Z���vNttZ�V�� �����õ#�C��71�X��6�F��Տ�>�P�t9�{��}��i����q,I��w%!�h��EЮw ����ռ�A7:fmF�P��<����<��"�z��>�6���:�r�/t�x�`?�NP�P/�����X��=��_�Q��9�پ�#d3[�e*S�j����Z�;�o��J�@����@Ǳ_l]�v�Cѹ�BmQ����b�ϟ;[�Wq\�:�b���%�=��%Z�&Jξ�{2
��nS�a_����u���P ��[�����U��i�y�vj�Et� ����!���>���3m�v��Or������](֤v������#g��1�!�Ò�m�ݛq��7���i�D}R�uk��Kz�o��s�ʁ��.�����B�z�oc��0H��E��Zm�@N���Zv|���U�͘h���N��� U,��JP�4'�n�&m1XB�r�O3S5�kK��Y7e�!d��h�d��i�*���>��\�G�Q�G�Yҭ�$<p�W8t�u��%��!��+.�'���b�7/R:蜏�M�f�.��q��7f�L�]��#R��L�RW�-m���d1b�����o0�#��:��y>dh��Icǝ�&�k	4t�ז���ڥ�vڏfQ2�m�����������-x�v�sS�'KR�[�>�49�5�]t�E���/�w�a«p�0Np�T�ŭأ{�Y��,ӻN{IV��h.xs����Iܧwt�sW0MD�eV�Ӯr��aKw��ڛ봼�>��C �������_�Q���?���9~7���U�N��y^7�[�o��޹�[�(�ڷ�:�k���m���罱��k�k�_����6��5�p��ƍk���kx�f�z׫z�#zM\�5�J4|k�x�����<^+�~{W�4b��v9�G���m��+��U�n$W+�κ�W���1|\�1�9�Q_��Ag������W��>w�m��;��n\����+�uw�Z�v�u�o'�mH�w&ǩ�j65��-4�\[Um	x1 g
�۔��/�[����;_�Fߋ��Z�_<��o�Ž�:�j�[]��-�M~+���=�b���:[�����=����觎�̱����k�k�!�-�lF�):iD��k�n[��j�_{[���~�����Z�l��[��=�3[Dx���7Fv%U�_���6�1�[b�v��g�)� C'!����[�c�Ti���[YT(Cވ��N6.�B�S;��vx�&��D2eu`N3Ħ���`���b�5-��dE�m�T�@'�^2.���.ݚ�!�ykm�anL�� 	iH��m퉥���+��&]�t������������g/��Z�{�j�nz�<ES�7�C ��Q��G���]5��6����B��Ef�����W�hlL񐜲+L�jEk��<���z�ϯ~��W(�j/�5�]Ɓk�Lè�@���&^�tQh�y|�<U���t� ����S�6Z���+�M�1�g<"�#��:�TX)v_X�c�����T�:��wλ�40\�y��׍�8�@8<	�����������k_����ZAN�kp#[�t��k4!��	�y��G�R����kZk�Ҽ>�2A���;z5J�����ܰ+d�y��\�^�m�tt��Ջ�V�eU_E�v<�,����������r�ɐ���\�������2w4���(d���-����A���e�s��R���`*�(+泓��㤭b��46ft��p��<�,�}��w�z�����`���w*�p:�vL��Ѭ���Hn�m��79S*͂���&�2�jݕ[���=m�h
���裎�ï�.Y���E���om�8��%��t��Y�N[X�3pŬRR����bd�n
�Јr���4ڰU_;�b[�²���T$�.�f�g1S�Yh��:;lo��*4j`��ʪMa�͌������yC=~�Vp%·�ԙ̽r�,
9��a�-\��s�����Ɔ�	K�x�S�X��I����o0��F�9�ޞ�c�S�X'2`O)��"Sl��4�H��]8��֬��8��u���
�R��E�4f���K��5�t�ҏ`j�W���4yX�{��	n�r��`R(3gE�M`���l,1�_���=����D����m	\��W�xU�C`T��2��u�IA�	�L����e:/���M$	�SCn�f]��l]حx���[�Uhc��m ���v'H�\�-��*���J}��	z�4�޸K��q�mg��{ol	_.Xj���J�~��*ä�ե[�"����b�p�t-��l�2g
��ڊ�Ӽ�*����9�?SB���U��D��v�/2Q���MG�S�V�@��%�����7��j�R(������4��A�k?
���-DƢ���L1Nǝ���Q�Q�����7n���i�a�D�ñz[������MVs��n��O]&���o{�]�@�����睃�PF��-z� ��$�oe��ުr�t;��ʝ���'�<ɺ=��<���L�e�6��Aoy����ݕ�R�u�<���|�kQ4�������05�5{Iw�vJO�l�����Y����{!�)�p�������R�aы:�����`�f�a&��e���|ZbAф.Sn\lF���U ����5Q�S\e�ְo��C,q���eS�H�⼼�z�����W�G[���kc2���?����Vb�/y�y�O���6�Fk�OL�[��JLf�+�T�yT�@���z��G��P�9�w��j��XC]]6R����[٨ж$���W��7��R�J������=�8�����^K^F�,��P`����2���\��	�	�_�iь��a�,U�a�A���@č]��6n�r���H�����3�Q��j����a���)��|��|z��W_��=G��aLד
v]8��B�s٩nO���k1y��o�k͍��9��͞�K
�"�?cMl��CeN<¸:G�����}�\V�X:���nU�%I�!�m�'͋<��d�ڢx��8s�O��ķ\=�m���0�0 ��?vu��o�N��1S�e��h��F��@������Me�+��ҖZ�g�U�ƞx�vMag�w������i����Oϱq���E�S(�;��M��i�Μ9���+���F����t��9�����Y�ܷ���KǬ[~v�u��v��:�(�C�㮚>۳���͓{���<��y���Wk���P��5�GPj�n.���mr�mJ�!]��y�L�8mˈ[�e,f��N�k�]s�ֽn��D���m<��O�x�Ru���[�U��F�m�W1�)�����ez����-�����AeO-��f����Zv����	�fפ��k5�8��a\�H�6�\l���i7|4'��T
`�ʜM�n�uy��P���-v0m����;8�c����-P5���t�u�6�Ryq"Oy���f��b��S^��:i��-(����u<Ś��ѵD�5��"Zk�֧)$ۓ�"[a	�j��F�Rv������{eXM��+=���vR�_���<YP��	�s̙����۾�vY�����I�h�H���YLt|��q�Q�]:�����Kyܖv�xi�T�jz��R�	XU�Nk�̗��Έ0��ɘ��K(!�Ǘn��;�P�yI�*�����ꯨͻ�Xqo������kɯ�A�o���4��ݺgn1�f��k=�è��:{}[HM��4zv7S6��h,g@�c)'�����(;�����z�X<�x��=�l%�>��\�C)��a�x-ʴ�*M��P��[+�*��2�`�A�M@�Px�f��dfT@��D��{���w:�\�<�zxl ��."m��;�L��Ȉ��Z�K�p�]u7I��L6��B�y�fsp����J&��N`a[�zn+�]oI�
"[M�Om����(ᬦ�%�]���{+C)=a?��xL�5e�@��UhWO�`��t����&�)c��R���b���D�=��}&/�qᐬ�)SyB#69��T�\�A�s����8�����~���t)�ōo���%ӳ�]���B\"P����-��3q/�r]�? ? ?��Z>k6���4�m�:SUe��p
MX���p3*���no e��Ѹ텧�Т6�H|߹��ssqe�y��\?o=���ٍf��w�s�=��Q��Y���cm������>�������<�j�)�m-�p��G-��Q����Q͘E[m�y�T��tuAh9nC �\a������N���}C����[DI8�{}Bp�p�W]F�6@ʆ@̯?m;h.�g�q�:���\��4�0ҷ�1jA>>�Ͱ�N�C�4 �j��gi�`%���bӉ����u4����nv� ����M�Y�Ddϥ�[�)j��w]oy�'[���h����.�����J��`��w�Pe
d�X��װ��*�9�^W-�oxj���I��Z��_0�'Y�X�2�	[�@�᭓i���k��e����`!���y��f���S����3\
~T�k�q�><��ߺ��0�g��bC6�q[������f�2�h]�Kt�hpZu��(�4n%�.%�Ω��a��ւ�e�iyۡ������N7��3`�I���"����1���b3r����Q�'�%��[�WTl�2�3\DHY-�".�f�*�:k ��=��Wc�[��p(�Ղˤ��e�#w��m&|:��&g;{}���i͓�{��B�����g�wF*s���Rm�'�-���Rv�nIRk�;T����@��m�����8����l�8�'^öO�["=����f�.�3��i8I�6;)��]����Me�ԷE�>��0o��_��]{���#Y���W��vC7�#�c��v{��X�מּ뛬��y���{Ε��z)����۞Ak��~��0d;�ݵ�=7N��9]L.�n>{2�H8�ڃ[�b2���]�w�ϾՆG�d��&����ǭvZjm�#9UW+�A�$v��κ|��{:�da才4w���2Λ�1���=[M��ڈ}.;�XCd�:�nyu�|��eS:�%�Oe�#ul��5u��w��08���U٢9c�	�20������Å�@�*ﮆN�(��F��ٲ�r+ɪv��r�����i�g-d�v��ܰ[��6�9�Њ�&w�m��L�h�GU�Ɓ���zޱ�b�Z*��a��m�F�l4�o�R���S���O�x�B`�;�v
A�����g,KA!�t�lu�fn�)4�m�Z���YM��ף�����m��,�WpY*�vӦ0���\d-��� X�s����Pj���T��ޔ��^�C;<Q\h�z�+�%��
]�鉅T�;��
�Q�z�V�V~"R��e3J�ܝO���p���KU���jŵ]hj�{H�E �׭��e���'{�r�\�t�z�y�ɡ=+n�kɮ�\���ݨn��:u� �W��e	\�9E�n�w2�f�.�,O���XeՉ��#��^�J��.a�U$u��ܙ���M>`���f���k_B�' �B��C��u�{�4�7�|�W{F8w�.4�E�\�Js�f�Y���&�q�FӨ����x9�\p��`�2ch��N����:
��}yʞ#�Ϲ<�v=������g˫d�	c��9՗En��'���4��u�U��z�H��+nX�+�$��2�k�1*��W�@�\q �M�L�I�)�L�G��% Z4��^���^k�+7�8�db����tbWk�bPU�x�#+Cn��"�8��;?J�4q�	¯r�/͋�)�5�8�@�諺)fq�U/'��&C"=��fd����_t�}�����X�_L�a[�*��*�VH��mEZ��h:i�k��6��o"\lw��[qQ�R�z��U�S�z�d;��f�H'�3��L��F����2�'�D��CM����|�-��XV�,��1.�l"6��C]8�a�(È7\A�����\�����������m.ƺN���y��]���%��!H�j"�� �@d��wI�j⏲�'3^]���mj�n����K#{��F���ä�)Op8�2���Z�[�݄��̛9d�j7M+�\�Vm���1�2�sѼ��%'s����N���sR��A�f=�˂ӳ��G�j���;��U_���1�Q^/�S����W���g:�j���l�gu͏�r��[Ɋ��H�c\�Ư[ww�u�W@yѹ�{��#F1������(o��x܂�wNw���{�]�s�^8�wNj���ٞ���5�-��;-|�Ȕ)��h�@\����kּ��k��t��{��ۑ�^u\�o<����|׌�&�	�ݱ��@w7<��͹�ƛ���h�g��>w��;�3�招��w��}[�a�]���;��y��!�c���L�:�W�1z�;Y�V�M�`�9}:��tG�f��5VI;�����33y����EMQ���r���e�=]j���A��C�H�&s8�s3�F�F�x	�}�jن�FÑf#Uj �ԧ&�O�.��8�%E2cna�Nt���8�q�2w���n3l�P�z�O�ѓfv_�Z�t��@�t���i4�)�ؔg:���մh��
����:Q�[Dtg\oj�|��}ɭR�ή66)����B��g�wS�v�ޓ�,'��y�}��'�)I�5���6#�@��#y^x��њ��F�,�E��(�͖�%1�g�\�2��%z��Ǣ�=�`L	����|g��?&�.ɒ�ɬ.�|��/��-���7���V��8N�YB��)��{�s���o]���I�H���5{�y����b�w��Բ�.�G�ݬ�j�/��\N]m^1����f�UY��Ԧ��w�5fI�Մ(Ls��4�\�}�t�.���,nE��UՎ��"���a,�y�K��wxۚ$e&���p��L����P!�6nV=�tK�mK�҅ŭY�M��vR�$d4�����lfB���<]�H�	����p9j'Y��&�&N���L���L�n�쪭G5�@@5��fq
��Q=��]D��Dl� ���U��i��_�ON�����ʌ��ԫס����5�cF�]b�y��i��O��k?)�C��~y���{g�4%�6�&$e\VW���~��s�Y���ӲUCg1v�֧l0�r�#�գ¸��k��5�M��D��*��xi�(U������.p�z��݋�X�޹ ��&!��ZH�h� m_��f���$� �'���cFh=	����:g(hvU��pw��U;ך��Z|S��A�hk��K-:A�����
[��8Q��#ʆS� ��
���b���ܑ�{Pzk�4�W����U��uL)�0��&r�Nퟃ�S���|�u&&��r���*&�'�����'Im*�G���6����5h�i�Ȼ�k�E��6�,$�K���M������:+��v6�Bc1�e��"�=1��<ż�fi�;�p:�A�*�-��eqf��k�1)=����S��Iƻ��b�
!v(㾼�/:���w�pg��?(EU�c����9;�f�dǛ����7�X�yZ;�\P�<}�1x��}$��k�]s;�:���l?��yܶv�n4�ߛ��ff�;�����3�Y,ƽA�n�T�Q�ωB_A^���ˎ�����F��M�큡��6�I=�{��K���B�/�J�X��������ojĬU�2ݴ�M�t)��;�iƬ�R�3�Ꝥ0�ن������L�@O4�ɮm_CM	�@P�q��`h��j��m^`�=�Ը^��*z��K{��\�
�_ed�j��,ږ��^�F�rɆx9 �S�p�8�P�jQ�uP	�n�C8ވ4'��=8��B������K�%�K��Vg�O�i
|�}��'�	�2�LI�T��ZS(�ܞW"�zv&a���=Q^koSwV�~z��=�?
�=���k��@k �5R�A4J7�c���|_7�㷮�H�A��͆�u�5����V�8#«+�j��h�"Nº�t70�]�_pj�'�L��Ɵ�꯾�op \�((��W͋a�R#��\s�����GO�S�_?�a`�N������֪�t�`�i�ړOdZ���p�u�Y^�5z����P}o���>�w��!f� ��0���4XM��*v�!�����[�X��� v��0M�X�Z�s^&v�Z��eE�݅+D�L����*e ��9V�z��� 3�F��ݽ�H�{#Md�6cuB�m�nq��j�8�����ԭ���6֠ɡ�]R�>�0!�F���f�����ǫ4S��j��N%��1�iSvج`6����0�l5E�tت�g��}T�w�{�����2�7��*�QK�E����qM+�����;_$%$��"�RQ��2��w�yLWNj�ǉ���ُ�ª:���Џ�����*lU�5rf�+i�Q�_��f���,�A@�v|�s�j	�{�T8��7���KL�+�X��jdϩ }�g��L�%A�<sɉy�Ff���Ȥ�c��^�����,���c0�c)�7k�u����(��L�:Iw��2i�F������u�5�F���c�̱�Z,{%���F_$�SۦP��>���T4�Xha*o��h㠦SϹTlvLC���E,�u�[��?m�mĨ%�W���u&���yn%U���u7���E��B��OR����=�аz�eGN�L����e'�`8��s2I�;��*Y���F>�N��MQ��Fq萦F��ٱw^��}�lȃdWcf�!&�'�|�)��j�ھ��Y�;4�era
��G�v���Sw2�B�<���rc���җ�.��[c�)�����7۝�,h�����I�[�x���<!��7��oTU���~}5W{�W�>��l^�Պ���~��!������"I)-�4HQ���N6�	S�n�zk�������S�5�EcE��s��V��~DTm,Q#U'� Y�K�({-2�3�K����w�|;kU�]f��fd�omь��:O(�g�`\9����	� k\6��u[L�2�jz�d��ظ�|B�	:iK;A�±��;;ըA
r�ɓzf��}
�f�'Dѹ'�m�"�bzbω�2�=��u��iY�=� ;��Gn�Ʈ�*eս�[���ۍ���y��Iw0���7�m5�`߇����RZ�C	���X�-�.��\��g�|�o�MV��C�]��~��*�_5�t��@�լ)��re���8]��X".�຦���U�6�{�N�_���{���V�<��� �˝K"���,�a�m�Tō�p��c�B֢�|�U�l�ب�"��zP��u�A;u�=Ɔ�S7|Q�w
�A�,Kc+�M�tD��>�Ƨk-�pV��Ա�a*6v^���M̕`��xni	SM��}4o{O*��zX��!��P�G^Q��q;o�QPW��H�����,�c��K
hiHՁ3���������ݴ�uRn�pn"|���*�Ŵ�1Pu��:���^�M5�]u ��W"�Z�1av�g%��H��4U4�@���D��
��Pw�׈�Mް�W�Sr5T�J�:�mMđ��*��7^�X�pX���H�1�In���sj�n�������I5@�,}��JدU$��ɝ�Hsܫ#��(u
�Ry�N�<�zqj��Q�o���ս��H8C7R4EC�����5���{���5���^��XY���)�n;}r��[m6�a��L�a��wo7�J��|�mq���bg�t���;q~ٙ{�:��g��HB� �j`L�Uȳ5�
�Bc���:0Y�z��ǭ�O�r瞜c�LΛA��z74ŊP�QǕ)�Bi�N��9�I�3�ɧvޖ��A�f
$T�{���;�u�j�����j��4c*V=UT=7�_�abQ�Yߋ�;6��n-�m��5X")����wlH��nӬZi��i�c�~���=/�����eڄV��7v2Q]QZ.�R�>�[���KY�~�^
�X�f���T�Y_m���`��ߋ*�"v͛�J]�/�J]u9�ݪ*[�Pv���px]�(v�Nx����罜�B3�QK3��U�g�M։%�w}a��T�İ%��	�׻�̏~fff�� &s�ڿҾ��bڌ탶��N�����*�;�B�zL6rZ�GU����ձ����]G����;^/(Ͷ�
wnT�T+�`O�ܤ(�k/~\{[���W�.J'?1���zR�Q@�M5���g�"�BK�P�:�p5�`i��:jMpA8���':@��u�vsQ�
�X�hkDe�d�U��#i�@�e6�sI�@�=��f�n`�{��\CD��*6�����y�Pe<W6����z��;1��b�nk*�����ށB�S�5�tKU�
s^ٔ��Q�V#_NP�C�)�K:��([u#��bn��Pm������߀�$#}�O�3����c����Lr��޾]�>&���/�3ӎ�d��byƃ#
t��(]�u��1 o{h
g8�� lP��*��8͆�q��I�����X��!Ԓi`ӈ�vOn��W�����P/�?��q���V(𞦃�t�{��t)���3ʡÎ��]՞zLi`�it�`�gi�^�W؂|Wk�sS*�u�3}=}��t��E*�ݮ��˝��̡���ɣ*A3��s�tI�rh�wڡ����r�93;g&��_,GB-Ҙg;���È�Rs�P�>�&� ���+r)7�u�N�w��giM6��U�s��7#�"C\/#��]��G����>��b}�˕D:)jVY���c˝F���g.{�3W:�*���<xpj���ʚ՚�r7�����]��Y�^���k�}��pvYЩ�C�gp_��n�K1!u��	q�5�^�o�xc#�tX���*̒�N�N'���y�znW%���X��zh�ݍ�<��ԭ�����+��å��a�ؼEB�<��5�S�L(w
�YeQn8I��3,1a9M�d� ���Д���gR�ۃ9-�/�<�rR)����d՜M�]w/l�U���E�f��/��1�Xꃭ�8tm]�y[z/O
t�;��]��S*j6;>/��^�;�EV1k�H�n�݊6 �ss�S�8t#����{g.����M�J�ܦ��v<�Oj�=GmAZ��V�;_Cm쒅�^����!K��H9�t���9ۺ��y���nL8�osLK+>�j�Ji�wR�f�[�
���<�kd��gKcP��+,t'.*�� #)�:��[��Gxw�-N��і:]�%r�bH[f��\�Y��`������jkoIXA��$h$�f��t�[+m$�')Z�'�Bڋg�n�w=.V����J����ĒI�	$�
�D��u�;�~��_W1��.��G�䌒c���xκ���M|��X���럥vIi���4��Q���w\���}�/�^��2N�qҝ�RHB�Є��i
{��x�W��N������S|��
%	]%�|���H��@�f}n̜��3D�D�ň���޹{ܿ:��(R��ۍ|�e	�10L{܍�43'�|�RA}W0��q�1��)]�]]��US���U��3��'�G�a�����;�wS3ZEަa��������P�	�<�ޓu����~�PL�j%���:L���U�'d"���Q�Z�]��\:�B*�2���,<�j�����Ʋj�е��n���h�]�34�թQ��O�n���,����Nh���뫝��y��k�n��6�����ܽ���
}�{}ۄaBQ=t�{���Չg��^��9��&w�=z	�����7b��)z��1ˋً��1�^���3���e�q]�bF���r�7V[E�f��َvۼp���m�Oڭ,Q�឴��^�;
g�=�Aˠ�g9�~�L���Z������[�U� ���C�fd/3'>��Gfⵜ�"��Ϸ^�e4��I�FR��ݻ�KP��Y>���ഫ��#��Khmu���ي�}:��+b{U�g9�D�7`���̮l��;�Mn1S��4D�j#�a��;%�y�����as�.Ih!�6e:���)�xUK�XQ�����Kr}��,\�b�X�4����;I٬�2�����r�^�P��,B*Z1l"�ju�&:n�d��z�V�����YT6w7�����[<%6�Al4�V�Ahؤ���L.0U��h�F���\��}�b(^�+V5Sۻ!���O���&��յW�yDf�C4�U@ʣ�]��T������v�)����s��0��b��Rϫ��Ƒ<x����۾�H�Գ1b�.=�z����h,a�|�0��LI~!��3��T����^j�D�)��4Nԣ�>�s�ޥ����΅�z�͝��$�� �߸��=�V�ѣ�9~��e.pj2�] L��a��̭0��O1�Hq[3,Zw�N�t�C`'+gS����@'G����Pϻ@�H���ud����LZ���K'�':_uz�M@f��C��M mz�w뱸
����˛m���C��Cj�b�T�4�ʬcGgY�M�|�;���N�H㪺�Ȩ�>b�;J�[7�I������Ux��DrjKKQ[^����6]�EO��ε�n��1���Y7"
,�5���O���.w�G�żnMp�N���-�ډ,ጵ����׷4j3=��M�oX�LX�tҶQ���L��؞�Sڥ���雒�:�4�Z&��m�o:�Z�(�wK����'{�)�ԃI��JZ�g�nml!��=��o/S�/�.n)������c�׌�L�ơ����҆Q��s��7Z=��勯#�-�O*Y}��������Ĉ���V�)V?�9%�6c���k-\/;x�S{VB����@�]�v]�AA��[DLnp�wa��5z(��z:@1�%%[{6̱���2��ݩ�,^ݖ�}�6
_�dnJ�Q��R���ơ�7�+Y�D�[1:{����K���`�o����Rr�1G�����9�q��[WT�K�2��[5���s�;�`�$��m֒�eL�T�a�j�����~�-/�����{3�n⽳���a�@��7O�c�g�Rq�3�㽼�cX��.S��7�h�ރ۷8�(^/Fq���#Ҋg�,Q��������eT��uoV93��ކ�*!�Z9t�Az��^s�,��tR�)hi];�0�pd������[6��1�'\�n�r��n���}���>�&Dy��k��S���k�����oF��1r�h}��UV,Qt�ܼsIٹM�j<Ko����pb[y�-��|�M�..x�w��`4&�:e">D��z.�0 ��	G_����m�gQ�O�S1'gm�H������W�ɲ���T�f��`�3F��\tD+�Y�עa��A\��t�Rɲ<�0	�1O79 p���І�ع�r�Ru�L�֩Cj�V�b�=GBQ�z������w`<�´uz,��Xݽ�^������|��t�y~���N�`ѡcm؂ܺ߱��v�h0#s��:Y�r�ȫ�ջz+�i� 3�FY(��=�j����U촓�z;dv�cwq�ڏ2\U�gW�@���n)�ɢ�z��y��%�Q^z�ۣ��h@r+$��kNH6j�ݿ|��+� %F�iWL*-��ۍ}5���th�c�)qGwĥ\
����D��U�3sy}5�o;�X�����fI�7+TTIc,cKSqE�"��ɝ���v'�g�����-C��ܤ��ϸd_q�S�G8��!��ig���u��cm��.�j�>:�pq�d-�K�fM=�1)����)㝦q6��X8����F�^Q�x�d�
�9�<ќ�mU��U�F��:�9�K��t��g�e	7��[:ں��e���Y������-2��MOw5n��g�ב�6�KD�V�y��I�{��̟j��F���$/�ު
�F��/���%�|]v���R��E�t޹$}}���v��7 
���)Vkw�aAbf�Q��(˫ս���]*��z���OypV���WE��� �E�i9��nƛ�AY�բ��[��ڻ,�yor��X�<��l�ޤ�$���Y3+�m�6!��7�?d���b������G�t�'�YW��G-U�X�@�����/��I,&U0�֖�hh�n��A\l�M%�mKm[m{R�jm�:F]Am�il.:�d���RM��9��ӭ>�g�&��Ľt�voM�V����ް�d��`7�� �;w3�mR����L�����T���u�+؂�y4���	�jsZ#�������깸Mv�]��l�Ψ�(��כw.�oŜ�f|�ͻY��1��l�-�Ӓ���D�2�X ���g��uO��v.�f�!P�{�u�,ҋTMt���k�3 ��LG
�נ���4'�{i��/ڰ�f1����e���Q���^�$x�d�Xz��6�TN�y�ո7��4�XD��_y���� ����W'�_\��e�AD���:�h����ͽ�$�;��u3!���&��1�.�Y��8�1�e+��IGY%�E�V��6��2�#;e�im���^D�L��f��Ҙ�۾��0���a�;�o�W6ii�a�c����Ò�W��kY6j�4e(��JKT6�f6ϬZ�Y�C]��8B��J�s�����˧����lύi�r&TK�˓x��T���v�lS>�ߘ,ԟ�N*����u$0�[H�i)�8+�F�hʂqNp��ލ�Ҹ)�n������[m]۶v[oX�V����P�_�����	�wgc�1��{oe;��F��[��~��d��j^����Q�\, �e�wd�.��:����R��J��!���s�\N�ے��D���xw�>����J��+�0o��*��cY�3�Z;����[���˔�+f�ob�v`s�=ާ[WS,�^tJ�-U7�;��sp��k��7z��	�H�g��S��v�6e���l�^��PRgI�m' ��[<m5�p8����ca�N�6�ȩ!�BM������o���u�������ֳ���9GS�ed���g�"+.+b�%���}�Ñ�(��g����0Ӥ%Ӄ|�o�+}�f5�
�������#9�U�M��N1�	��űC n�:c8��q�u+�����[mhүu���� I�e4��t���������5 ;nUn��1��<����UҘrC6�_=֦0�]i�"�/T��="��4;����t/��\2��e���eh�	mjp���Q��=��Y�R��x�"n����81��1#���p���Ufg7Z�H:+ N�=F3[0�O�X6����JvkV����Wyb� J��ښD׮
���	62]5.�5`����5�R��5�e0[^�5�����W��/;yܢ���A�ջ#���s��������7��K���U����Mi弧����=��Ā�*}��ӓ>pe�2���6A�\dŖ��amQD�=sxE~�@2�g:��ז)��ం�,D^vr ��m��Ha[R�v�X����=�g��Ț���=��>�[U�Ͻ�O��ӽ��)��5�+Ѥ�$6�j1~m������YN50��(�}�/�V*�.�_GF��j�TW��i�O&��8Nсu�)��7�Q���V��V��i�xۻ��o6�7��@��Ȫ;;g�L�1�o��]�����71;5;I��j�=�g?h��Ea���$ԧ8�`kf|�mf[�1��z��I5��T�N)b��#���4rm��:�`�7�����+i��"m�+��:��Bv�s���<���S�]��q�4��Q���;�{�wܪ$z��JZ����4!\�'C��fL,��.e�u��jO�g\�@��WȨ�%��0r,�kC"M�H�we�]�`{�c@c��t�w]�hm�`��6�Xv�N���?����u���~J�q�L�V]�;�F�!��\x7�{���l̗'4W!qY�����Ү%K-�4n�L����2ﳣz�C�;���U��)WA-I�����P���(Zg�����ڐ�[�z�Sjm�z!�IWϠ��6���n=v�������<󁂦ydYj)w;�3}���&=�)m'�Af۸!	�BC_�d4"��%�D���_�$dX���E������?WXf�6���vVn���8e,ҹG(�T�IVњ�3j5�VQ}�Am�>�&j��Cv�r
��+�6u�����u\T�eL��h%���W�R��;��$ݾY�֥7��z&��v�}Sb�%
U������ќ�T���p�Z����2�"^���Q��}�vڣ�7�ԫ��np����5���R� .�7s^�~�v��>�W<��(�νY�k��fب㹓��l���Gp� @�LY��6W�^.�,F�t�mh��-^��f77�a����= V_0�jWS{���.-k��XiX����v*�Z��h���Z\���!�݇���$ӵ[��t����D�����+DE�>#6�����e�<��-lՁ�`.Ψ�[��Ġ��م��e��qwھA�����e���+�T�61��Xt���L��,�KC�Z�8j>���<�d2o9�U$#�ŮNO��������V���d�iws%b珻��ڽ�ڗ�Zk�,a�:��>w�w꘰T��3��`������� �|nGy��07�d��W�y܏���w(�����^�ҕ㏮������I�x�ޮ~.z�_z�&e">v�4!O[���!�=��2H!%B�(�/W^.F|\���~=��@C2eB�<�κ_z��$���т�wǙL��Ѳ�2$)0g�׽qI�&P����RDI2z� 14�'�Ē��H!����C1�d��@0��pc1량 ��K�B��e�
x*���E�vK;��8���[[Դ�͝`ۢ>=A\n+�����?��)��oA
��7N�~}m�T����'��1�����f�Լ�g��ڊ9U<�l��2+!,u�.���	��ó��%�ޢ��N&U3Ce��z��ZJpS���&��:؈��3Gm��Zu=�)��՚�����/�� ۅA$�#"��t�z��Q����]���i�� 4��4�ͥ��2)�^����H�盤4��D��k(�fƣ=>8��yl��|=ۑ����'A{�E�^���w�7w?%Mi���we�x!�\��^����>�1Ù���}�s�M-�'2O{n�OB�(���l�������^^5��܏����e�4{:������GFC=�Ҋ��MY�\VL�Kqތ�Y;n��澕�LK�y{�U�7�¯d*ᬷ����]�L�YU�W�Z�6唵�3��7�_MMw�f���q.��ԯ��C�Ȭ�:qeS�5�{��o��
��7K��p�D0Y>��F�Ǥ�6l���5k�A�y�&
X������l��Tg&���:2+p���t�IQ��{�4�Ĺi�gN��βQܻ�����x�Z�mu��-0���$ɮ��Z���G�f�QBs8;c�\)ao!Էi��Ȧ�T��M̤ՠ�O�=Λ�L�dI���j�٪o�Q�)���
:]���*��Rs�@S}ݕ%��)4�]Nm�cvW����<&����LT����*�+�h4� ���k�GCJ^�lR�1qu��-ׇd��`df��rƁ���d�^t�����3�$�6�=W ��������OChr�nq��'����}���{|=׻uz��k�r�B(wp0�9SL���Tz �v���5�y��IA��kBZ���Z��$Y����=��'w
��L���6 h����R�48.Лd�l�f�yh��ث���8,:6�����=wNh���A�EG�3|��M��)���C;_dn~|���7ߤ��Ķ�L�gwPB���~\%h��'.T�]���b7�[6�W�=��ާ�3����8�q�>����u��ƺt���訑x4��Ni�p�[,�TP��������4rAL��oj����P�j|�t�t�Ƣ��YTҭ������8�N��1_M��_�)��*��
z�����KJ@Lj��N!Dg?��e�_�d9�9�Vg8��3������)y�;�����V�/���7R����i�+z��G����䝣>�[�nXؚ���sRV9�ig7|Kɵ�,يc�{6e˅>̽\�a��F�Y ��<��o�Is*5�ƣ�S�^i����OMm<�b^���	�Je�l1�o�#j�b[��L��1a��V̦�ʼVZ�,�Ω"��Ǻ7<n��^�N��2��i�|1:�ߕ[�୤�j��R����!�. Ƥ^���2�׭����.�0R����N�������d�g�w�3D�b�b"�ZR�tF�,�Pl��F}�JZ���\��M�p�M
����0.��2m����;Y�O�_D��y����L�\�5���UM@ƾ`��隇����hh#Q�!�7jlPeu-Q���#������Re ��h�?Pj#����WZ�j]��ieM2�m_2���3'���v]eW�����z��oZ�W�Q��#/{Gd�ᮭ�ڝk���]_�4*����	�7��hz�}�gt�8�co*�1������$�aW��|�uTζ}w�a<3,8o��}f���}��&p������P�y�r�T��Q�TBv��֢:�)�(o�ʈ{�1X�N���M_���pN=�Y53�Ir1��ʉ����[I�0y�r$sh-0�Ɋ�)��Y�	Fd�i��8�
��31aQ}y���vK躱�dsv� �lI�ƪ���t�7gۏO,�4��m�0i��~��R$��v��E-�-�y�{w�}N���S>�Y˳y�w��7��ŊR7Y���V����%nhh(�r[&��N�\�D����^t�̥��-U��\��ٷ}J�xN5p*�b�P�w�u�%b��/$j��EVF�t����@_�����+��#V0�vy� @o�
s�����u�2^G�C��a�M1����xj�����w����J���@��`~�3�b��sw��jFe��jٍw���&Rn{R�~�8�ǯ�31G^�{�M���u�r�ݿ'�Y�S,ԫWD�g���n�R�$]�!gkə�����E۾nёǨI��v#�����̦���ѭi���i��K���һĿdW0;-\_P���~l�١UO;_��ZR+@|ՙ���P�����ᱼ�=�
���ʷ��y�~�l�W�`�9^N�km)��`첕vk�<A�Ξ/�-���q��=7�;�&OE�q�u�&X)IDpo�/ ���򕡮��<����ݷ��8k;M�Ph#}ի&%Ʀ�]�x�]�b�w����K�1�!����1��-�[���to)��h�b�79�e>4��
pɍwS��\NQ֙���^pG�~H�K;��m������U�)�bW��ʼ�u6eB�C&�d�j��IR�k��|}7��]zwx[�����k��CO�z����g�~��C�s��D��Q�$����S4��ā;U�5|��x�+��eg�f��7-��#��Wd�[�p�a6�K��Z��}꡺+Lt�*���!րi���Lt�~��Z�OW٧˳1#�B�m#��
�%��L�6ce�z�KU#5C)�K{�^�I��WK6�>B;�-�3/qG�Wlwb�D��2�l�0�MXÂ������ռ�8q�'{/]<c4gt�|_)L�Ɖ�����bY��Ձ����+:WP˦��:�v[�.��EM]&�,Vn��D�*(��b��:9�^.Wf���^'��瑱�o�rY�T��3�ϔ�l�ӣ�E+/
Ow:��P�b�l���b��Y4�45�.�؍�çA�m�U�(�''mZ�Aے�u��������]�l��6) �V6�0�0"Z&�c�{�w�TC{B9�!O4��T��%��J��^RكR�q5��a;/�����I
`d&��R.�����N��ʚs;����>���z���WHB�`�{+<��C�MUF�WDX(���k�U{^4�i��+��ܭ��ɿ5D���h(�,d�/b����M\��ƜPI�Bnj������:٢�$�����cu�>��\:��i?De}uc7�+��X��=��e�:AYm#���|h,߮�1�*|$���ʌ(�@����%�7zǫvи�X�|Q����t<�g7Gpɼ\ݔ+/Tm[F[&���:<���y��˄����q����~���ذz��uTj�Ev�;���Ǎ��yzy������N֮ЛIB���5��8/>��ݍs����<�zf�*�A�v1z�f���������.(�5�7zm��D��X��]l[&�K,�FV���S�R�Z�4è8g�:�ww6�����-���F���6�tօ�D�t�b�S^�aͩ�~:)O`#�!V��fYy��6�r2�����{�[��T�Oő�F���xV�'j,��1&�ba��r^xT���Ȳ� bd#EĵM�a�AxL����Z&�_�݅r�SF�f��ǘ�\K;	�ݠ������u�uN�����!��r:��������s�pp�)�K�
���y��*�Vvw4kۜ�s`��lC�{�er��ov��&&�ư4�Tzqrn��Z.��ZZ�pta)n&D�v�V e��U4[5�I��ذ � �(�\)��&m���0b�:���[�������ש?Y*�n
���;bgrb�y�	����D����IU�i��j5��r�c��RΉ�:33Q����;I
�Ȇ�r��~����od��z��T��U���w0,ե�k���'��|���U�E&ƬON��O�T�ʦ@�8ѶPU1��oϙ%H&��`��d�`�N�m�dd��j��7���p����q��=�V��xޞm�R�-�3�v�z����Or,��c�l�ʾ���Ǫ�s�`":eխKE֞��T�f+�`�n_F����2]^.oo�M�I'��Q��4>F�S��}Ȇ(A��Ҵ�U����ǌ��[�m��aN[��^n4�&�U�hwf�1�̳T�P)�7kN[�����1��u�Kz�7������4�;����tN���*Π���Ǧ�2�v��%&qU�C`j��]��IrC
bM���i�g|�t�j4�%�c⮶�)Q�n�z��W�ٌMn�$F�}��E;;f�I�x{9rΉ=}�䒂j�5Y[@��2��.��JP�^N��l.0�"�
�Y���/��2�m�d�v��>w:Z\��b��9�p�3_5��zfެ��6�+kLw�C\��F�:P��h�{i��(��r���C$�0
.ȅY���
����A�U��;���N�tRVJ���G3�tD�=MFN���t6n�^�ǪtI�ۀ�K�e��.뽹2�J������{I��eha��g'bƲT�*��b���+�l����B=���W�,Q����D�vm^*�'yQ!�ah�@I�=K���c]3:Od�q`	�b�t�Ω�eb��퇵�Ľ̠������6p�(_MǍ�����e��Y-"�&�u-2��S)��h�Rt��\�� ����长<ÍT�7}V�B��t�&�l��Ai�-\^�Ky�3g�C�R1�)ۗv]�r���J�TXZ��Z�&��u\�s|��J�'o:�b��ee-�gH���)}ӨQ��9�yO��=O	�ꔾ�(��#߬^�oT�|�uϕ9z6��KJ|�V������7����-@ԡ;U��x9�k��f[m�z��ݤ�����'��}�����S}�f5����\����v�-8�-Xpl���}������]��x������fH��2%1��h1Ρ)�'θ���ώ�؈L�ι(��n|xR���A@�7�;���;���?��7)$�H�z���1�ur�w;���<r˝����K1��>8{��.I~wb"�
��n�����r�3Lh��{���z���?;pD
'ιo�@�O�]{�H��̡M�Q;���&�O:�%!�/�z���5�m|t��HJ��QG�D�A��$"q���Z���bqT7ҽ��6I��\^�)�u��[z�ܼ�	�b�)���:.�W�U|���Y��-�`rY��Ѥl�L2��|.)!�Ì�)d�Y��^u� �b�mxT"H���hO�!�@h�P�i�!�*�{t^��
v��sw=�f���b�ج�}u��s�u�D�[��L�����O�)p�?~T/=4n�)�-�1r��� �L��Ǉ��s�,/d�B^�?�r�P�wR�y0�w{�6#����а���VB�m	���Z�� l+'�V�f<�C�*����R�U���5'�����n&��6�i�ܹ�(�UcY�����Δ����|9x���U�un:>�{��$�E�I�~�r�l�~���"���Mi�%�;��_�]��wt'��4tm���Ƽu�d!l�H�AKg^��pP�gE��[�Awũ��y�&�\�c���ٷ6w���bM���b,֗E;|���~�����c��R�A��ʶ���������K���]�ΙGa�*�CG�=q�.唫��82���(��aT'��E
���k�9 ��}g��`�c5��]=�-��]�GA����K��eQ����
ܚ�B(�3���2䤴ۄ��3�o.&��YաM��޽����YP��z�J �`b
5�y�3ZjZ%=e<z���֗d�6R
ſ�Cp\�����ɇ]�K6G=ʹ߳�T��1Ï1�o���.��i�~)��H~"\����֜�L��[��*�vG�lF�E���=��uz]�/bvv��@r[����-�ώY�d��ӷ�"��l�Z�m��7�_p���s�p�K������]�̅��?/��lY{
V��麛حhm�>�ea�$:�.�nH���M��޼��q��	��!����E-�F��_t����H�1I���Z�V�7�k]3�}SE{��\�޴�ܘLY�pwM��^�ugtf{�5�V�\�����e��ReT�c7T5�EQu���*�Yѩ�^�,��R��5�o��al�g�67Z���'{�e#'���4�s�SP�n�)fV{hz���/���;]k �-9=�DoT(�n�=���[�7^�	�~�����Ǟ�D24���������^��#��dn�t��am�dw͙�_L�-�=�T	�:��o�u
�H�A��"�d���o�z�\}�gU����ۧ��L0M��DhfG��k,��T��� ��K�v"f:��W5�4��u�rC���CĂwt�7���1 �n�鐵��������'� -Y�7����T�Մ�^fS2��jbLӖ��r��7���ݬ`�R���:Q� :l�H���xE�I�-�Kq��<��@Չ�� ��随�Gz�z��V3փy��i-���ax��2��t��Q4�O���O�H�����O}����I�½��5�f��-���ń����ڛS�s��t�
���9�Y�=�m��؇�в��Y�3R��_<ffL��k�T�e*�wAF-���m@�@e^t��|�5���v�%���׻ԫڃ����P��3����D/���(ʸ�^�ߝt܎b��ʃo���T�`���Ƭ�/4<=���4�[4�������2��a�jj�f��H5���:��#��nm�}p.��6����3't$����sd�4�W��7't@U��`�|�g<�{�TpV�S��M�{+iee���'�]ibS'�̞�k]����.����&���ȴٳ����A�,I%�h�^m�>����`���S�ݵ:v�����[��ų������3��^��\Ɯ����έn̕;V  ƥ5�M�5�>bMI�e5���ZZ��8�$f��de3'h׌JlT�g��y�M��[e	
J[��
��-J7,|\5�+�t���c��[�v�W���I���N�U�ƽ�G��D�d#��gϞ����z{�e/u1ن���Tct�D�͡����)�x�²�+6՞����bu�G�l<�����^~���FA
N�;+ƹ�k���\6ŝ�7m��1)�������m]m����Z��Bc�����E��FZI��Rũ4"S=�KH��ʰ��V�����)�����!��P�t��R������a�7��xVn�v�5lZ�����N��9E5�������/���.�=NNB:�V��R��c�$�}[�B���T&�+:+Y���;~l���T�e}���+'q���~����N���^����E{����W�x�̾X:�F�>^���C7�}���8���p}V{�j����V����"�J��3)� �m�L(ۖ���+|�FuyftT�)�nǃ��WZ�Tw�f"S�9�X��<\��z+�`yu�R��d�]��c�Ǽ=�.W�U�t���X&<u#f�J��sJ��T#�6
7w�\{���Kv9t�n������k�e�1ܬ����f��s��9 �K��y�1���{���@vP�x��R�NV�0���T�������ӝ֪t�;��a���2��49��,�4�B,C��9i��:T妛m��J�.*&��%$l�tf�6M1�)IO~-��W�b�u� 3�`iSU-�(4l�kV�$�_q��#'p�D���l�_g�cB�R�-SJ+5����(�-�f]愩6���:���ت��mC��;�$��W�Z��ڦ������;��E�Y"��x٢Z���R��]H��|jw3_?yH�!ޫ��/�X&ڕ���M��6�S�, �7��6�?J|/�?v��5��^t�
�+ :z]=*\1�z:���]k���'��(�vQ��X�n��C;�������^ѻ�W~�E�+��֫
lHn�d���U�e�6ݞL�cK������?�����ۂ$��CdY�jj�!�y��qjI꡾�E�C`���U\��a�QF�b���.����}M�
��1x��^��N|���ب�mZ9����к��;��jkm�M����i�tH`���pR���������eM��q�=O�^L�1
.�w~}�i��h�t�������If�%-��ݒC��e�CU���਎��#��lÿLk���~�7�A��e
�}熹0��!?�BQ�yK��*�G��yU<��f�@��k}��~����F<?��L���]�>y�(���0�������0�D{btXv�����bDl��dl��R���ʤ��B�0�y�˗T{����ݧܻ���A�M6G�+�L����"p8ï>'�߮O�D&�{����W�ر&��0yic�NR���e?1�i�.�~�dZ,p�-\���I�û�����-��G.���j�l�DE{�O[�F�y�����2���W`ѫ'w�0�7�4>w�`�r�u0��WG��r��ǥ��~ ���>���`+�"Ƥ�c��;*��OtA�U�ry��5N�|�8�ޫ�\#z���sK�̣�\'�����i!ͱ��VC�*�K����o�U�&U�?~�b� ��0kzw�� �Y�'G;j��F;BXMD�m��DY��lCZ��?���F��l�"_�{�G��hi�M6$���+�r�Y:{{�"�1�	t��\�m[��t��ɻ�&[;�b��=l�P���˥�)cq���%��m�T�m3o5�����w�~�1{��'��˼�.%��s�W3�w=T�w�x[�v��v5U��tP��I�[�֚�a䩨x�ϐ�C�O�?l#���u�c���q�ӆ����v�/�ؤ�4B�]�SO��~pÓ}&�+�Ѕ`�Q���H:Ti�� )e%��1���I[Ռ˃��MVr�λ�J�F��Қ>݋3����Wa��c�Jz�R�9�evMo[V�y�;��Y�-Z=ʢ����yC`��7��p����#r>5,��׊�Ԍ��%�4kB<���J�|}�gn}��ܾ�C<q/s��������o+.+�@�x���/�o C����̳S7Ok\*d�1�:[^L'��Qw�����e=E�S{D�w{e����t;���B��/σ)��ǝ������T�^}�}��;K�S!�����,�z=>��oD���g֔ӗ|��¢ry!���*1�5)l�w�r�8QQK���r�䩷j�=������]1��	I��韛xl�w-����������,s��L��M5�IzM3�������?�X�ؤ��o���bs�BBT��#z�3���5հ^�FKsd5kV][C��,*����4�ѷ��{�����nr~WB-��ӗ��<�Ju}(�>�N�l�#+�����?��9��P(�	!lƀQ�с��A?��qn���w�y<�|��}�_����g�}��*�S���i@-���(V�l��X@��T��c�WL�L=�'	PFj��L�l;�nHqwk���M��ŝ�9��u��;�b\c�u��ms���wVP�%�;�S(������Wq�v����Mi����87�%�� ����Р8s����؇%B\״�P�lc��W�
W')��~�<�K͛P=��ʆ�iƳ:�[�f��%>B�����md��b���=n]�tm���]�lv�6ۇv��qɅ��e,Vj9�-��ˉ
Y��ܣ�+�����\98vᭈ��z�RF���M�`��b]�#��Cl�ƽ\)|D����2�^d�-�8W]�Ep�Ut� ryt`Xf�Q-�,�f�]�u�f����<4��3,�C�8�����]�u�L˚��ξ9Mܙ���m=�+
� ���K� ��j�3�ܖ�y������%�1Î�Kr�����[ⱶ���]p����ԯ
����j?)�'������Vx����3�j�ճۘ,���%$�!-��iF�Q�S�$$Q��1X� ���*�fs�h�B��^u<]�"\s4
ÝE&����gX٧���0ĳn�&nYۊDu&3Z�H���_;�H��,��	���se2Uwr}S=� �i!����;cMm�`�v�Y(vs������+��c<���Zj7(n���I?S�vQ�r����ڙ�M9o\\^jtt��N����4⒞U�y���q��m�VƬ�;^꩷�X"ይd�͌�3�2�EA�}%۰AxiZzQ�Y<�ݺ�{�Ys�2�[�����˼<k�j����<����,9�t�*�,��e"mv�\lu,�CY�!���Wvxop�R�XiUA˵S������6�(�*vDt��wH�y����PFL8Д"�xU�L�����İB��1���A�)����-�l!!5�#6ٛwܚP��{���4'e�3�`i[�A�6E\�*.y�a��݇s�㽊ʎZ�]v0i�����7�F���37S�NsI�'�I����0�x��Jvd���T�GwQ�a_v˭�t�Ç:�%�h����A!$I�J+����ۜ�^���nn)]�~y眝���\�9�.%]�A͹tݔk���u�w��:�?]��O�t�ߋ��WLE��#��D4.	��Ѣ�\)&E�"ޫt�[��+t�4{�h��<�E~.�b{��ơ�Ш�wk⹌c�n/{w;��^5@X�,3���e�u�>�i5�~/�E����y����%�EKy�L��v��o�x�0�$�R����0HLP�A(U���u�Q�DNn5�a���ؒT0$E����6�}��-�p��YMW���`����C�0�ȿlO5�ޢzz޹���_s�z-��a�m���~U˅-=K�0"�l��\�iG��?1��7���*�$�)`.<ǝ��*a���܇��z���.�X(�<9�ߙe4�)�3ÌH\�?|����||r����O̧�U�X����D��%ߦK�j�>җ��27�M�,��'��m�e�&�t=m�K����)w�i���L5��0�g����V}�d�i|1|zz[]D5�Ҝ\�t�<������0��^�;En��B/���QyL{͏\�r��ɞ��"xk����3��:_[���Le��0|e(k#�n��]_+��L�w��~�gu�2Nr]x_�^]��t~�O䁅g����N��-�;�Ql�͗c}7}�/�`��DjT�ۤLʡwW"���{]�KЪ���i���Օ��s<���B9!é�V+�c�\�o�;s��JRP�՜V1up���5R{��cm{<�fٞc�0vΘn��h��UC���f��C}&Z���|�<!��4:ط�� ��^>̟��l:��F�	��tJx�)�G9}[8���D7�5ʆ��aM��ZØ4ZDV�BSÃ��5f��/)��b��e�����;&���n��BҚq����S�q�q��#��6�i��b)�<��q������U�E,�m;�x�X�QF;����퍢Z�s�3	���,P4�WY�M������S���pd��^�&/��co+w=tc<�M��.�k`�2���U�����;�>�m┆�mt���$�����p��K;���Z̦�8�Xռ�ղ�_1�#V��8��˷.�.7�������=���R����*7����4'n)���<����׉�ܼԵ�\�y���TH�'{��'��6��ݨ���-LdO??_�eEx;0v��p��l5�;��ؽ�Tn��u����3C��҅A���1�_re�2[}#�qY�/��w��Ȗ��}'Ҕy�}8Nfݚ��ӘlU�ygʛf��=�S�G"E�P���/,V�}G��l���vw���~�*v-�2M[�SZ�zfi�����¦i.����jo�p%�Q����|��a?S��Pq3��gK��n�-6�28�C�,�zR����.6Y�ǩ��cr��NC֏�ܪ*�r�'yXs,{���B���d�Q����`�0��l����<a�D�1����z�ބ�D`�<\q�kP�9����P/���#?yV���vD�>���Ex��#�$�sk�/-S+�\TEL�5O�b �&S�,�[>zÕ\r�U�>3�O����N%��-��;�ߝ����Q�*ߺ�o@AcӐe��n��#5�,N}�-~_����t2i�Ղ\��9��������k�	箎�<��S#+��0R�>m�����=�i��YƵȋ�W{��R�`
hq��g$el�&n��3)U Dk���S����U�~�*��Od��M|�}�.n2;�����e!t:F�O��iʶ����w��zA)����j���t`��;�m�g1W�}��4���t���݋��"1�1��p�6Y=9}}�. �@� W�.yؼ$vݳ;��z��޿�Z���s�OO;-*�1K��Q�B��ʞ����%�՛�3q��"g��	�P���ilEx�t!��	xED~�&��Db�|i�;��a��c��T�1�����R��+�ƏCT5�������<7�R��!Jz��Խ@y�c��J�4SC���5�E�����s�~ݑ�/���@��;��P,c��MvX��w{��K����8~�c�KOĘ��)����j�͞�.������2�j�5&
1���Ft'}:��JY�z�E�5ψ��/�f������Z��5����X�dר\d�q ���g���S~:!�&Cn����<\��-��a�:ܫ�m��n���EӬqgo
J�x�VIk8зO�ea8N=+{2$ي�j��+z�Qs�]F�i����h�&˽�N�b��F�y���Rcw7�k*9;k7�������J�xĴլ;�|o�1��o�R�|v��^"{�{�2r���s�M�nz=W{L*�C�̗��V��ZΛ@�����@}r��&bzL6�e���f���{5M��=�j���A��ٝ��]:�/4/�W]b�yC'�yP:f|���L��w<)�+�f`��x��0�p���|����	ID����8�\~�Z���=k�I�w��L��L�CSY�O7���Ls�f��_!��m<"i�;��t��7ͼ��X��ت�=��fK�@ثZ}��4���x���AnUN�<��ovx{��-[��}�g�Pa� ��2�Q]	̻[��<����9;<������'(c����Ƿ�ϊ��$l��]7c������-qH�'�hae����x�����=7���w��W)�����}����k�/�� nL.�Zۦ�^�a�������1���Esy��g>U�X���='X6�{y�o-Be�X��-��E�H�e�\~������f��3HI��C\G���1�l(��M)�L�LT��O�!À�>urVw���K�Gl;YS�7�nz�N6z���:�$�wM;j1��SL�["������WKޱ�qKX|hȖ)�/b�.��<��v��{I��F�1�X�<�^��A[r&
�񙬚_#��jr/j�h�3�c�n��6�0�WT�i���L����-h:k�c~��|�����i��;W�L_r�����g�(t�k����9�}�/n�k:e��3��aZ�5�G��qaȇ\r��Cz�c���{k������>E�8V\U�Qר��m3P�/����xd���4���8g絵�����u��rx�	}���diW����c0r��!���:��ٟ���WoyP�ߛf�~��lL_�ڃK��g ����B���H�絕�kGI��=���}�S�Э�VN�!o%�$y��5��.-Q��Rd�yǷ)ovoF�S0gY��v���@C�{����m��/����o��`}����FƵ�i#��d���ݽ���EX��Φ���e`�'�;ޛBVz1��������.=� �P�c_C�-���==��8�db�6\'Xj�CW��w~�%޼�:�PT�;^�7øχ;�7F;N)/l�b�����s�ltE���e�(J��6$����Y�� ;�\^UK,��R�)���߮�c.���C��e2q�6�gAr���9��2��\�VŻ
�g�/�^����c�D̘�j�.�'�À��ɗ�_���pZ_���c�V �pٜ��k�ܒT��� ���i0��x1ϑ��}X���!���u�]b�s�l64�uʄ�
�%P橎���k�ߞT���_��{�#���$�o�6�'�4zN��\�>=�n
_���+gz!�E��a�����؋��M��O
�`ϖ챢�iX�	���dp}⌍ye���,��{�Tv�����)�_|��wcB�x�����h�����殧+��}�K���u��<�1���yDTκ�>��Ƚ[k^���z�fϼ����hJG��a��wg	~�A��BP�����9�~B�'���v��鸋���si=�щQ��s�9��1�;���~P��{'����F�k����;]wHv��M���S1�&�.k�!gO���3���U������g��W|ś3�:|h���I��7L��3�1����$n��o�	�B�.u�/����tg�c��k��b�Y�uL����1������`8r������:����4|lb�R��- ����7�"���EՉON�\�%�Y>�LLh�x�/�V�_z��g��'�_�/{7�I�}纨yq��!�/��CE�b�S�@!�M�Ƴ��b��⯋�,�H&������ϣ"kA���4��,욪Ďr����j�ner�S�}�|��.?��3m����MRu]y!� /ߨ{�l4��+H�/�y�S��vg_I]+n9��/��m�_WK��{s�K9��*�T��d��P!�mާ� �4�섭�#�4{Ix~�[�e�(m��P�[+��x����� �vw���i����[�`c�uFBz)պ�)�<�.������:6�KZ��$�_)��lz緼�j�c�w|
aF,j3p��4��\o-y��'X�e����w�߱����4`Ŷ����Mn�K?B�,�YM@�C%��y�c�yG����F�?Z����b�'y�{W�F������5�p���FU�k�!Z�ޑ����(~��O
ңxl���[<��Y]�,=s��g��y�n��b��/ܨ� ��
��)=0c|w����_y�e���t���ri��B}r�d��j*x��n�#�D�b��vщn//���~bg�*� ڽ����y�|����]��f�T���{H��T���r~\���>7�����d1��PR��e����1���5-���!��U>D+��������|~{P��^��U�>��Ԭ�2A�6KN�}�=˅Z���t �M�y2E(p��K��v;�%��jp%�Ӭ��r�����×-L���
�����VY��mY��1���jI
��&>m�KcM#���r�a���[�K�/���=�C�Ǹ��=/������3����G�c6{ ��vP�)_RC�~�~���\_��Cע�.��T���%OV;���1�kg׾ϻ'�!���Qc܅g�(�7���G�Ԩ5�Zi�+�퍰k�N�D�k[-Qp\R���H9��`���~��_���<Q�ʥH��u������{��ʋv�l2i�[����h�ml���y��N���P�uo�X�P�P6��&{]�ݬ���ƥ�vF�9��'S��|M�<U}�S���D�����f�iT%�ь{�6��>Ĩjs�f�gK�z79ϳ��3���N�"�w�ˤ�<�P�������ަ͋{{�0v3�t��8��)g��3%��7P�~l��B�_|���r������/7ޞR��|����p�ౘco�[�o�f�9MV=L��خA6jއ��iwD�X�L�WXegr�L$�a�t��_6:̒������U��ٛ�y���#,��N� r��n}��Z�;���oQ퍑8͵]�ݏ�.�&<�#��R;����-b�)�=C*4�=�˼�L=���[�nCz]���'
f�9=N>�P�Ywr�����׸�[aV18��T�qg>�+t]h�8X >ee�3&0��w.����sm=܊��^�)��!��s�m���U�2�n��[	��௜���	K0XUP�s�5杩�C�!�gJ�Q���l^t�^s:;�����nWo�B�����e�G�֙�0b=�[�f�z�v̷� �p��5hu0�w>:�� �Tu]o|�="I���9�O�fA�eC�xܾ3�m�>�g0Pں��SB�ݛ����^9z�L�A6{�Il��P��z����t|[��u	�/��9$~:��<h�����Aq���H:�[��[[M[N�xJ��2bR�M���`4����e�4s(�^�s-���M��8D�j�嶏R����C	��
):9����	��4+-&���b�8ou
3,�Uy/�=QGk�E|�b��20�l
���T�%�u�#&X�b�p�n<�A��[@��p�5J�t�-@Ma@Վ#E�bj�/uom5N5�ԑ�k'��%|�VܘNH7��__Mw]N_:һk� 	s1�:��;]X�f�穉$���<��w]�q�2eNF[5� J�u�)���ؠYU��5��,��mm������J�묫إC���e�k<���M��+�z��(]}G�TQ�O$�e���Ǚ�\Vu#�k�f�,Wn�^[o�c;'�T����FY:����m%��t�F��!� p�>������I*,�}[on!�s3u���$�r}�ę���$�Td��d���;�����+�
�d�6��"ǳM�Zt��ߒ~�v�����v����y��b�5���׈��H���I�yۭ��ƹEd�}�7$��K�^3���,[���wXѓ뚌j��F�c;�?=��(f�ҬQ��0��4%���4�E����;�͋㑴D$b�И��ɮX���w~y�o�:��;�%��뛞�u|���k޻wv5��\ܷws�+�9���76��b�����wy�����W<U��Gww]I��� H�g��Z�ܽ|�>��wu͞�Ϥ=:3���le�S��}��K� ��l��f~o980"����6������ ��R��H��K��S����N�Q��qԺ�>;�
�����ɞ~��a9!˅�cTq�L�L�ң2�@գ�JH���Ce�þ�5F�z�c����ϕZ�/�]09�15��SM�i�Y��O��أ�Ӡ�j����F�lºؙ�.X/5��gx����7+�Xd����Z��������:��PR���������y��XW��<��m������}�ϫ��`E��̾��|� 8h����_��a�)��4���8�ߕ|��|g��M�''�>\M��:e��������/�<WT���S�&{��C��g�}��_�_y@������b#j�~g���!ߚvu�KvY�Z)����=0b�D�}�����9WU�GH���8(�b{ϔ��@�t�Fʖ��z�bo;.�/:��ԪÜeZ���Bl��,n��~Sj�δy�.<�޸�^�
�s5����q��̵]-VQ�<$���9���$%bs*^��T0��&A#~ozbT�ދ���о�͞�*_1���+9���__$6V�ׄwX�P於����]߻n�ߡq/��^:���<�pש�_1���Lϭ.�mGd2���~0���t��U-�Sa�o�Z.|і���G-];��ǧJ4K�m�[\���]�B���sI��ia�@�S���snkY6�,F��w~�ϳ_�`�|׼���<�L�����W��zaz�A�o�j���/�@�L�\�y]�����k
v�vX��~o#8��/����.����Ի�kڣ�!�⯆Z��w���<3�X�j��>���7z�!A@w��7�ز�� ��1Oq@V�Gz�/��r��3���o�1C�y���<�e�Ũ*;���$�[�9���X����m�r�����Y�Gy`� �rZa���Ȓ�H��ĸ>�x��kXvr�ft�k~z�W/��vH!�wC:p��az�Ӡ����9���]]1[2�7tž�3�]���q.��}�@�1]�)�ꈚT5�4i�p:$�f�-��Y��	q��湝u�-y]E��.zh��|��VЮ^򟹶��.��}w��}��C��d�9��Y�l������P+�O������A�q�=������m����'���j�я��?�?4q���Oo T1�qq�m�:�l/��URN�c�-_2}���ѣ�/���W��]l29�1P<׺^;�-�)Aq^J]�A����c���4��=L'��� ��X�!p����8��l�2��W�%�%_���}��(�y�B�����כÌ ��N>_�u��q��u�-�p���h���bz��gAm�h�Y�µ�87~����#�s����><k�3�3�mɴQg��㼡�� �j�����k�z_��Us�3�ϩ
��.1,7Z��T�kk����g��u5CH��)�d��t�n���*q���a8�[_7E1��g�}_Y�9vެ����5<|��k#��v�h�nVo;���J�Q������x��N��qQ�4�)���L�v�.�:qp�a�P]�SP����Z�_#ta����f���E������ߟ㗟@��%��6��k_��h�8w�n��Ȉ��iq���y:#���&%�6
������rS岒�<|��Q�w���K�/>�\�	�Oz �c�	�خyqښ�V9ط֥,'�x9��u��Mn�g�.�;3��עy�6�q�,�S��ډU��l4��[hI�ѽ�3�'�Eރ�ZxX�&���T8T��O6*�?tc�쵱\�z�z�*y�����Pqq�P��{�L�$��;kM(�)�/�X2����e�Y�y�ƨ/n���E��wq�-�}]�0z/[����L9���uwmsC��1�~������R�p���۔��	D=9P<:?T�P�}-�f��^T�Q�)��ːZZT��(xN"��]�})�:��hU�i3��T��D���z~�����ˤ>��q1������n�^3��m.��*f��7��-�u��d��jf��n��]�ͮ��KJ
�u��2n���,(��.�p�r�;���c��	{Qm��=Q�Y��;��9�d��ǧ�M�:AS_;�ݵN�XIzd�!�Yo���-�)笄�&��2@νu[�����~'��Cc�q�����s��얷
o����z���tţf�#����d��6a?dp���(���} a$��B|�w�7�b��t�gqq�c�����&y�t���D=Y�-q���0����3���m�8���9�S�����P|"]P�{c ��'�9�ZG[leC�&PD���uQ���q��I��W�YKf�~r���r�D�l�O7\�#]�w:m��W1։���^R&W>�Y�<~��`e��wS��_g]k�2���yd�ؘ7�Agܳ��$��>�H�_���XQ�ULvf����=4Z���{���K(����rx�ʷV�t.3��}Iv!�n7�K'��aLҩ���m�*K����B�u�_"F�z�;�(���g��^��lˑ��V��.��҇+�pU���lh��;�;ZJ}�5U����Afqc�c@��-���4v�1m�>������ms9Qm��M&uI��3Z#t���lS�����B��mq�oQC�N�ӫ����wE	�g�������/ymFK�g��gx!����"Ag���69�\׶���N���a�z��M/��?=cם���]���˶s�}c'fP�w�������
�@�y#~��먅l�����{�˟��liL6������&�?yL��1�z!�F�Ks8�~�~�ep|6Z�)�LgTF���w�!��_8��}e)㢛�D�M�$�^��p��!����D^��uj����+g�kV��H�L�*]�͡{����(L���z��pp�L��K����>���3兝�/Qφ/�A��yc+�=<��[.�
��l��1{{�,��Y�L���!&��WܽZ��(0��$Iu�du
殧	��(��Xk]���Y��|a4)��Ii�o���w/,�A! i�nW7['�^V��v�h�gIe^᳇�*��WϺ�mE��r�I��ʇS�^r6�,rH3�3�}�U���M���SPǼ79$ں�/�l��]��v��6%V[�^>���>�����#��O�:�8�'>���IQF�4��>�ޡ�JQ���q��%vnO\��ܩ�����j߭Hj��<��ߺ#�B�s�l.e��ygGE��t���R*��W���&=�L��凼��m�!�B�C2O 9���9�+_�y˫�l����7'���81�	���t	�@hZV�~�{���ڪl����Θ/����;&�<��sʱS�Ȏ[�G*a5��D!���eݡ������x����2yn~g��֧�yA�[�P�M�g�'ޠi�ڼ����!�4�L�s$y>���/aVU�L�:g/����.�%�����.��F5G;f�On2e�x扪�*�/�vn�Q.gOC��_S������D��7�,0���f�yä�ѯ�+A����xIz{��$�=�c�3�"N�{W���E
�W0W�vy�e,o&�~�M�)���U>�I���nANH�x{&^�D��5AW�M�,v;:rI����s� ��c���:Q�Ж\�K]�����;Yc:�3Dq5�3�}n�{��f����h>
���X��C�_f:��w^�Aթg+�[4�˓L�v�+9���N�����u?"g/�8s�5�dd8��[�(����\�kev�1�0X���ً"�],��g0n��7U'��������Ks;x�c���� ��юd*b������t�Z4��1�e��UV� �l[��p*d���关(K�9�x�_E��m��{:"�a��9�]���ڮ~;H�EM����q�\�W.~G��xٴ���~���vϬ�b&o��O���~��������k�@�'�Q�HW��,r~o��]��K��^1��#"&{����B�a��1��Z��.4١��c��)����W���GNa�����*�Ҝp��p�2��'_���(��\���<�k��?R�Pqq�P������bA��=7���So���m;���vg��>�&7Z��u�P9��ͮ�\��PX̧D�:�(8�|�ϱ�o�ٰwB�����P�ܒ���|�V�ÖY���wX\�n��v����V��[�F[��Q�X�~1y��^$��2l}_)����&Cs�n1���E��g��}?R��4� 诂��~�'L\��C�0�^�9����Ҷ`�,��������s\W��f`T#�ּ�ؾHw��	�4�����5��)��B)���߿_�a�5x6ſ�f3�}��ߟ:���h1/N�f�|U���u@U;Ss	O]���Yv�d�p.�|t��xH�m�wFz!St��!<��M��������vm��)n�m��i�>��eJw�2�{��(Tڋn��֦�koB��1~S�4���y瞍����|q/�}�����Bj�TX�g���xxz�ꇾ��}H��w��>VaW2��EHxQc����N�!SC�d��;�'�|27NѼ��g�s��}�E��5��U�0_�Q�̺����L��1cp�83�7�\a���+�3a��kz��v��0��42�c��!�!�W���M�YNl�+1%{��w�mw�,��N��phYV��c���j�ʮ<���Hc���@��4�C�G�ރ#sIY�c��-־"����օ�m�tK�	.s���ۇӼʛt�U�T��h�9�ԧ�i��4�}���A��!�C���X�+��;B�)�}`�����!mNsi��`sU���:a��Ǡ�A���);����TK��s����z�];��� A�n}j�aS�����1�Uu���2M��yl�lɵس@�n7�Z'd��xקs#ЫTY�o�w�>y��X���_�ܚ�;[ƛGc�7Jrc�@�{���t�ݼ5�z�[�a�6TB'uK��(���nD��[��������k�yQ�g���)w�wF�1�
*q���)r��ޏs�]D3,gt�����Pձn�Z��gm51���B_�9�*��~��,��o��A��[F�u�!�E4Q`�H\����}�7�~��Vt�}�o��2���y*��Fx-/��8W��YT4�	(�d��K�!!_�RB mD%��k�\?}��Qd���2��
$n��� ���m�/�dsx��o.�ot�ɿ�0��77t��N6q#��w3Miu�q
��g��,�P�P�{4��!2�2]FeK�W6���;��^��Ws���R��	8N/��:'|8h�:�`�r���C���vl������� ��~���צ�e���ܶBu�֕Df�a�'>�]��`�t�󱩷y���>������[��i��-Y�g�^�k�TCFA��%\�t�C�&���4��ȑ�X�Ի�B�)+���;:N瘮��C��n�d�ǯ8r��! ���4t�a+�/�W:���A�$��Ӽ��12����MG��@K	�XlY�Q�'��u��C;s��O1T��npma[I�+�p����Z�֭��Q��f��h=/sjol/F�Ö_Lp�9����㔛;��f��<���zޓM��]��n�l��rbhr�B񩙝�4a�R=�Yap���@��z��4mʈ��ڲjm���Ѽ��o"QnS[�\K��wL�L�"�H\AȋE�C!((KZ#��[Mw�i��c:�Gee+s�z{)H���L�� �ѡ� q[3A�YS�aԟ�C� �QὛfN�'J6��5n�8��ͦ��:E=;�f-w�VeaM�`�[u0�8��U�{��+�"�*��L�@�f_AquT�D��\e�tԉ�{j胬���ԋӹ�*�:%i�@��Vhݫ���sӱ�Yۡ۵��mӡ������J���cq<{�S7�te٢���X�C���m̈́�hf���4-a�d��1]��[�$�Ǎ�y�&���c���(fU�2�L�h�=JW5JċѧDc�W�𴷲�&&�oX�N��'�T���)��ܶ��G����ói�v�u��kWש����sS�S�>���۩>���ݛ���ǋ��%1�;.��>����5p��!tb�?wk���(��<k�h���}�{ݶ.���^{ڸkx�s����ׯ^͹�v��^+�b�sx��ח�}�U�ι���y�wv�6���<�;�nE�\��|�s�Vwcn�u^wc\�s��+x���*��|��kr���;x�$�o�F3��/<�x��gwW��t�ͷ8��^�ׯ���ζ�Rj���W����R�v+x����[x���m{�e5�Qmй��o/�{���M�u���$��˭�%C�Il�D�D�I��nY��x]R��t��[?gp5�����PBU�{mĮL��z�.c�3w[W���l��-�2����-�q����~�d��:��<G��{���5][��7c��i�i|����6XzK7���Ͼ��?�m���jH�枣園W|�q������9C�n��T�{A�/�cMs�3�L�#�oc��L^�!mv8�R�wa0����&1F��θ{����z�T����;���11���±�G8�=����SoAeCL���þ��Qۭ���+���̇O{Q�a��j�3�0�����^�ɼ|4�������QƤ��ko�q��,%��5V)la���z�ͽ6�F-�K-�r�i�Ɖݰ���4wB0,�S�ߧ�U�>�J��Oϥ�>Vx�Ky=���e|$��v�o��Ύ�L5�+?]}T6�ц�.{������������3Z12��n���!Cx���S]1������~�C���O��7��TU�\O¬�g���I9�$*�JO�Y��
]�L���)�����;�Wrq��0ܻt�]�K���,��������t���-��'�>d�+-�M�r�ĸ�����މ������ED|�O�'{��4�g��Б��Deo��xl�~���Tk���M���f��p���:�y�G�%����Ju�,�#���o�`�qԑ��2|f���}��<�j�����Uv7�zx�~�Ǿ֝z�Uڟ�g�tTaB|vP+�=伯���a��uӺpq���\�&}sQ�-�C�Y�OR�k�������7˹��]Os7|}�X�_���+�t~'�Ș��RӦ]�Yc�D?��i�%�.x�ZI����l�ju��΄c�U��.����%�ﲪ���n���})|My#����^�UsʋrB�ʎ=!��rj֟O�{կ}�^�i~���w�����Ȑ������>�Oٷ�੡�[AY�����xUo;�ݠ��ˉzw��6�v�ȗ=�,0I}�On_Th����g=J�Ѷ���?�%���0k�կ@c,MOI�A���J��ĶޫvwzS���p����wvZyG6-���d�苮-��9�K�E�u������_)eh́�ܑ)(��.JV�뮶1��sM�DG�7����T���C��o��p!��gJ&��_���S�MvE-����-�W�ַ�/˶�/�X��̇���T�s'!�D���}7,i����$���w����c�[��]E��r�[�:c"�
�^�ni� �.��/�)���^�q*5���[L_ �,�僼O�n�ȗ!���#�Ξ.5�F�i%����5��tԧڂ�
y�w��%Pw���m��5 [*w�<AS̞��1�D[�E�b�g����M��N�۶k>������gݪ�Ƭ��W!����I�\U����ܚS�,�>8x��<M�]s�$��Q�/�@׍Mvz
vFj��S�s^WWp^�"�W���+����RTK��6C���6 �������F���ӯ��Z�߽�O,}�>�����M}��?{]�Ԅ9��X"ԯ}��g�۠�0���=N��̫ЮN8���-O���;F�س ر���lr�Z����Uy���挫"���I"�Nj&�)�ǭ{�<���A'1&*lQҘ4%m u����t�Pk�ti-����ꄿ���1Z�*;��`d|i۞���tj�$�_�-��̶Nm7=5Ď����.�ê�>�N'�\ɖ�J��?������T"���j��>������\�i�R%t',fmML]]pg�?����|?Fi��[��I�6vQ˻>�'�]��AZ���6-��2�a�S�(s��3��)��w���ن?\%C���M�de�n��M����!�eSn�0R�	@zr������d�쪐'.1Vsg;Iڍ�_W[Q��%x�����OSu3��F�	�.��7Fn�r��A_T^:�rƇ��ӹ`��$���Wŵ�{����e�.�k�/Wi���b��g1i�Y�d���CZ��C�����Bq.�+�ɣ'��8�}B�z�7!�;�n�)�m7����c:;K3�&͝��˒�Ҕ�xyPu6�2E�E4Bfz�G�!��o���Jΰ��7/\K���,�m�X��9LP�zY:X"�7������KCȘ�fB8�ë]��ɗ؄?�����w�ݾ���D�?��Or��+���_1^��#T�㗪m373�ڕ�vů-�!ɘr�����US�!C]Ż]L�K����P ���y�t������
!�J6��h��[�=��!&�\�;A���ά{������� ���*-���덖����[�pi.���0�ܠ�S��#�Tx�Ogμ�}'�ƽR���X��n��6�{�ٗ��=8P�\��]�L�o�>�z�b�{�;5�����`���\���?F��������,^jg^����u�x����]�¡�2y�G>��[q��?av[�Ђb��6Pr��2]F��|ki�n�D؅��K�5:6t�9��f;�<{� �7��g��듌�� S�ߪ��ɔ����:
��3��>8te�3�˹{�%�ꋀ�_LCaG��2���h�d�ov^��w�Jy/�-<�EXy��Y$E��8n�b�Y�"~�7��7~�z}��������s�>Ġ�7�a�N=\�P������G��U�t��Ə�W�l��<t��x\�5|����|��ڄU3�wGޥ���g�9��8)�=�H/t�h��@)���GH�-Vb�cc�F�nh
��Y�n,`��$��^�<ޞ�͒�g?�L$�f��g���ծ��X<��iOM�C�&��P�+ހ��r^hz�a!����>�5�B�Ѽ`�Cӡ�������7tT@Ly祆�	�.8=k ��c��+����=��O�j��V�Dg��~Tjx��������̟����s@φ����S�������:f*?ET����T��zc�&�k˞,�q�}7x����� ͟��]��N͝=K�YD�aJ�H���YmP�|���}Sr� �X���z��Os��q_�D��5�3�1W
8���J	�t��B{O`�* we����NHYӝU�<�Ҩц�b�OU=�n�W�rgl���6_j��]�ϝ_1��x��ew>q�u	���xZ����Z���t$��r�%�`���:*�+mZ�������0���;���\��c�3ϴ�ֻ*So�q�`�E�L��\�����`�"��O�e�i�e���m`Msͩ�*���N=����*&�\a�^���q:�\$�d�f|៵f��O6ݞ�)~>V}���e�.4ޮ��,v(C[��w,����Ĺ趭�`!>�'��C�c��P���]�����S�팶]�	k��V�p��8l��%<�v�͌��G�_c���2��1zْ��.�^e�}����ʤ�y)�30x��~�����vS��>(�1����7�:�s:�w�P��î"U�ߚ�5w�fo�y�Z�`�]��/l���k�/Q����� ^А�Q}c�ώg���3s������r�XKƁ|�V?<Ns���N?�)N��[a��⟦cy�X��;�����ʍ��/B紐�"x��'?}�~e!얛��z�ky龇P�&�6��:Ɩ7L�h��^P��z�ՊQ�\���r���^6��&c�]]�VDަN#l���2�{�
��(7ި�:S���YM5�\��[�XZZ7��Շ��h�+[��^�kթwF������#�\�f�.SGt������`��Wݻ�T����9r�>O���gß�|��1�e�X>�ͼ܎EX��y]o����R��^&�g��!E}�<kT/�5�ϲ|'b�P�Y�y��r�[L��\���KϝyP�{��I3���~5������o�$��\p�|̺�Z���L���N��s��P�0�q�)ν�M�p�K�4[ۚR����-��J.�uS������3��"⣼�[+6WN:z����n����{(�c�#��'ۚ���-0�;0V<ҫB��|G���l��D�v]�I���]�\�c��4�m`�]�Æ��2?���r�A���`�ܼs
��0��ђPV�FV~���3l��Y��f��TT���vTY��6�^m��F�l������g����vЛ����.�vwm�t�iΝ�+T�(lgNw�k��ΥJ��k:����W���>�f�bԍ�̔�x���A�9Y�sgii�}�'����I��:-�T�����ͪ��:�����up<`��5��+�:;ˏ��^6��|rخ�����4{_�Ќ�ɑ�3�-d;8Y���}h���/���*o^{��<>�����|s˽(?="~�?�4i�L�����{��)�l3�Q���ý�)C�ɐ��Ya�&֣\��f�]W��֭�t��yif�/�na��T�a(�]��r�E�1\goO<�<ɛ��4�9Ӆ�>0��B�:�I�:�����Ƕ�WJ���j���ю��:�=6L�za)�Bs��Վ}�*��T���2�z��
�ìa�dN�'������p��={�W=U�Oj��e�c���چ�k�1d���z�:���)�A�x�(��A6nh�zz�ώxގ�Vw&W[�o�02M_q��l�q{iyclr��es�r�3��ɳs3Cz��q:�"��N��Vn�(~܈�/b�u5�x|g��(~��f~W-�1*J�v-��>��̣���w���-��*��r^Yd�o<#?m�:f��Q,Sä5[���|�V��i[�F�o{i��6�vKр�F;a�M�r�n:fP�k�K�3�2B���22e-�R\|zeOۨ_�8��T̂�L��oua�j9@w"����?WC�T�✅��K|���ʫ�9�t<c�y��j��S�O��Ҹϔ�T�^��
��l>�������+����������+a�s)���s���Z�����d'���2��xX�{'�$ޠq_�9���I�$��S����)�C�c�W��+�Ͻ�7��8g��x�^-c�P&��W�=�@`��=R����7!^.�pwweq��DP�ƌ��|ǾD�?�x�|����O��M����umn�2d/��ɜû�% o�yt[�,�;�}�[1�T������F��ϸ���k=�x��ni]�,����9E�Cz�o�u�yB�����t�T�d�Z�VrNk��M���1�P1|e�ۘ؝%.V,�n�i�Lf\X�R��ٵ����t��Y��Y�7��u�ať���9�i��.�L�e0N���HPz��W+�z���$�|�����4�U�6�޲%#N��q���L��S�w���}fR��F�`)k��+-K����ٍtC)d�t�/�s��)v�#TF�]�f�W���~x�ụ�}X1����M�+�S{��/���U���!�V(���x��b���wpa���!,�]To��� �[ع�R�ƛK'*Qc�Wid�x����9^ڰ{?nʡ���n�r�s�2&F�-����X���;��������P�J����]�Ep�V�WsW 6��{^�5}W�x�b�K���6�CI������p�e
�Gr�7\�%h���4]�<�w��Q��̝��![��ZGnTi�SM�����v�T���^"fo۲|��mDކ��V:�����ZXE�p�9;�Նՙ���u�١�+3�q��[BfKGN�\܄2�E[m���w�����CB<�m�;b��kv�H�k��jŷO��Ȝ�s�h�h���ҁT+Cm��ǽ��|/�&�C����$�2�ݷ�w]�.f(B��nN����U���)}�b�u�������I�+{WC�c��C����6�YFw$�h�ޭ��Ҩ�D[���sF��G,X��M����<���:�-=��V)�c4�k��mO���%}o��*�ȭS�{3�B�R1t8�v\{ZΝ�S�g;	���I:�א��B�T�Ŝ��d�V�W"�N�yu���V�4byj�;�u���R&d�����k"�}e)+/�c�)r<���.ݺ]�:����+1=�����w'��8��NDhG��|�c��wg�j��ȏ��
�㽼�m!�'S��ig�k��c�;���[�9��͇p���|oW�7k��;U˖�-���W�׊�s\�\���/:���sֹnZ栵x�6�z�kx�J�;���x�"ߋsk%^*��m_Q����N����E����W��:��6���x׋��X�݌l[^-\�x�x�x�csx��k񷭫ů[^/��=��U�uz�Z����oZ�}o�V�f�L�����s?=�IeK(��ÍD}&oxT���3U���VP|�i��+4ѳ�	���3�o�(KC�����^[�T>�wO�F�3���*�lw��Ox�3��ŵ���QA��Xy�j9��X�]�C]��5��M�Rҧ�Ι�p'P���q�Ƹ�ј�Ր�-��nÊ��+������ab�~�]D������!�#�2�q�<����7�n�4u�ɮw�R�+�;���R|n�����c�+5�j-�g��n=Z�=t�e$�C�B{0�&\�_u0&y�YLd`��!>�"qGEQ|`͈|���Zi�����6R~3��V1�$A��i�T��芷���^���M4R��{��K���0^� 6����&��d�m����Ǻ�*\p\J���A�/��.�{;�j*q�Z��ه.S�U�0[�}��g��U���,+M0uP���v�䕶OAO4���|���#S!�' �e0���sz�_�Lϕv���d;Ͷ��[ݪ`[=�U�ʀ�����j���Ɠ_���\(�9���V2��QU��P�(�7�!�m�UEƑ�%�N�q�XȞ|zn����z�c���G���ƿ{����*Fg5Gr|���w��u��2���!�ڧ[N��Ϫt�s�f���H�ʺg2� G?�0�������-�<�x���{�?n�0݋/w��ߙ�@�le���'�6Pa�+4�9�|{��B���h�^4]�,�p�z����x&6`�/~q��!�@��)*#O�*w���Up��D7%�\��6�n��Y)OM���{6ӎ��u�A�y��޻�O�1|S.ۻd�J[(R��7tӵs	�t�vK,ƞ0�r���]m�QC����w��i�u�w0��w�~d&�;��t�Q�z)�7��.Ah�b��e��ly�U�q'5~���u�|<��C�/1�.�omP�Gc�f�kQB�)k�G�L\����2s��T�+U�T�_��$���A�^�g��0!�X�^�(o'g`�»�E�;�We�7.5׆�,"�Dn��W^��b�;�$=���1��7��h[�6Ŋ��2s�j�����Y��f�1T��ՀtP�.q����N>:�T�^�Lk�2zZ���.�]�6m�`��?")޲�nƵ�E���vq�vK�Gl'aZ9�m�̛ -L8|��~�C�Y�7yo�/�A���v�M���;�5���ʩov��=퀡v��N|��)缆�]L9KZ���=�R�����/oޕ��M}<�,7n�>�c��ۛ�ii(�wOyڲ2�����5�3�wO�7T��v�Ks���On�9���q�Ɋ!aG.�~�A���� ��T����KO��<x��~���S׹���w���%���ӏܾ>�f�J�g��+J�5�P��;��]
dǛ�(j�������'����ON4C���|Us����+�v�S��G=�wk��8O@h_�>��=�Dg��K�}_��A>�a^�\�;����k�;;��k�У�ţo�>�޻6��;�Ǭ��{n����oyS4�H�W'nr樮�t[�(�L_m�'����̜�܌��I��ƙ:�<����	�r�!`5N��sA~�ђZ9��`+��������T� T����VIG��f�.�s��T�{�Zל1ן}���Ȝ=HK�6/�w�C֠����NyO#��`�緐�}�ao�Ŧ�d2�=,E؄�f��~����w�������8��g��L��SwKK5��Z7��	�tv�M�ZX_Vt?Gٕ)�;~5��A~P]\5�Z�d��h?~����^�#^��ѫ�\쑡�0�W�ëEQ_X�7�����ǎ�l[�8����y�>��j]���,*]愕�!����Mb��ǯv�u�5㛅Ӆ�7x�����G,�0�̻f������6x�G?i����ZK�������c�>�ď�b���7O��:{l<2����:���G�1o��̜LIVN �����J�z|��>p|�-�����d��F,J?v>j񫧩�}ҝ�h<:V^��Icg�#���:�������iIv�Y�pf���o��0�����-������u�"��U6E
��q��T��5�yࣷ�_!K_|��n��I?j��oN$]��&�KS�]�<�G7��κ/Z���������@�s�W���}���[�=H��|�c�ou;��C��1Y���zG�����<[��Ǝ5��H)r9����g�~����рw���GMTù��/"f�tG<&j�R���h���\�%�xO+����}q0��ݓyeؘ�S�'�n�`���̒Gmn5�����~T���&k��u>7�n~��Z����w�M�}��xh!g~n�m^�8X5���������~��f�8����O�/bt='k�]��/�	������P����{/��ư5�B1��V���nYN�8݌Ž����u���̧��wU�.�;���&=o*js�S���q��f�1���?X�E6Y�K|;j5����b�.������#�ojQ5ҘF�[�
屁Yp>y�+��XY��Fg_ˉ3�����u���r�of)S[�I	�@/ې��N�'�Ǜ�U�sё	�oU\6���_m�y=*�����a��>עo��$ݵZ���ږ$������_���ȱ�:}������NZ^[��|��j'o]��1{�㿭'ɘG������S��s������X]y�Nm��۟�W�s���۫L��w�;^v5A�S�<���e�r��j�,Q�8񯾹�s�t��z�A-���柎U�!�{x�kJqչ�B�,^zB����m�m�h�8���%ҋ��٤,=�'�xc���9��\	;w��$�xN���k��}��k�R�X>ǎNd��g�U0�#o�{e~Ϧ�����&�{�x�5��<�|Ǣ?%C�h��ߧ
yK�\�^?�enj��� &��H:����`>z���O���	��m���R��nt*nb�v����]�˨�Sd��Nu>����b��n�}3p��S�F�mu�J�]��7'e��)�C�[�{��u�w���:X�:*�׭���nG��G,�b�Y��/��c���g��䤅4�*���Y�|g,��p�$w�[�����|(��?禐s��ȕ�N�%�������E{�H1}��b�L���W1}�&�x�c5��yו�-��6��:�c��V �Q\�`=,�>��e�t�ϟ���7���BX�<�9L�i�����"�[���\�ҋ{sj[3e�\��al���b]e�vq��@���~�Ύt��2Z銦��\T�}���W`�TH�=�!p��_SN����2/,-�ӶSq��0�w)ܷt�m�׺:�w~̐#(��mחy�<5�A}�3���s6=�l�=�+x��mTy�-�2��.M'��e�q�:�c^j���w@�{-V�M�S(N;��4�~i����;��8k��7J��F��T�d���`�9�����]E�}8�^l(��`>�󵭫�GF��'jJ�K�wϊ�p;���U'T�F�:o�=!#�zBިH�z�#v��W�W�5���k z��w�t����g�9���Q��S�R�z��	w�
�Ǯ�w鲄�T�����z�w�gT5�;����>5L�~��@PTj�4�����m��I�;f�(|���X�̞���~I~�z}���-�Z�k���7`������̗���H�|X��s�~�ǜ���D`�}����<(��Oc>�m�-�N<��t�ОD�<��0��](��,���D[�u����w���;����c�P�9N��g�KC���%�{_��7�4}���P:c��{.9����ˀ������S��ݑ^�,��D;b�Q�*�MJ��;��U��qq��< �W@�z>4|���2e܇l�B��t�PB@����8<���Ӽ�Vw�x���6�e��Oe��C���i��k�㭃mͽv��V;K �}���F;b�zak���嵲�G���H���+'sȻ]�w=y�S72n&��f�\2�ݨm���<s�=I�bm�ƞqʓ�Wv��Cu�:���됅3��k��wW��t�)�1�;�2�P����
���>ζ&�����7����,�[<,7ex���;~��֯��_P�5��v��OR쮩���v�f#��J�yIyP��v�Ѧ�]t��)��+�y�Vl4�]�I�AsT1ا��(cje��Q��uNNz����.�d;�-����ҥ�u�gٱ�~�D��A�q�
V~2��AK�ޝ>KSx{/ꡒ�Y4��η�����=���D_CSA���!��c�sĚ��S�������͋R�����N��t����z�sD7��픲|�.��.�M��-E+gm�m:&!u�����Z����8f�t���^4`�C�5�K�gd�wL;����A�r$?th��De}H��eݱ�[Z�y$v+'Z��W\��t�:�9�~�\��a����{{��TY��
%�l2ጎ;����?�U��-�ļ�}�����ME����@�����wz����S��J���OEt��l0��vjty�/%ɪ�á|0ݫx��"ݗVeECH��9��7���]��G7�|>p��:��q��6����x�����S��%�6�	�SOO�F����ϑ����������p}z�/�
]�!�����:럞�k�Fqڕ��
�I^3�vq%}�Z�~	/��M�D�[g��羱�G<�k��>�-�R�r�ޜ� Ť��w�ۣ���NA�WQ-�9���/^ޚqo!��/6V��#����/ǹc��@9��:&۠���y��O��S.�p\TWgn#�����oNz5��d�΄��	k��N��)G>�3�#�t�:�8�OAN�SX��ǧ�2�߅0|jgo]Ps���T�|�ֆ	QJ�q�F�S����S��Q.>������(sz�v��:��tՒ7��&7t��74���A����0��:Z3ę�Z�3��x��� ���s� Mkk�]�V��"�'O� "�z�@Hf "�j��#�?��yJ�n�w�������_�y�?;��������{���o�����jɪJ���]6�U%�m��t���j��QZ�|�j��ڵW�ڵ�j�[rֶڿ�U���[m���}j���_��Sy���V���WZ��������+V���ն�� b7FPi	�S��<`�u�#`�
�u4����he"D�!��$�$�d$� �$�A	 Ȑ& (@��%2@	$����F0�L�BCI � ��$��2@���1$��$I�$��a��$$!$��0$�J%&f�b�dI�P�&D��HD�  �$����߭~~_�켿���k�ߝ_϶�A���B���4ߘEB��-�"�/-W�W��Y����2���,J6��(�H��(ȋE�$�e��RfƤ�d�-����3FJfD�M$��4��Scc2��ME-���5%%4DX���i4fk3L�Ȓ��l�&IE&��,ő,&��dhO����r���UP������i���B>�H\��DV��iW�kU�����Z�)5�y�k��R����=�|�(��C���b�����\:���#vy��>@���@�s�� l�=��o@P����_�~�[o�TU�����Ϟ0��֩3�K�m�N�'y��,C��W��w\ �%��~$\� ���4��t�ox�{߲��չZ��6�g���Z��Z�{Mjڶ�ڵU����gt$�%���!4(xXG�w 8�]��ƦC`]�3ɹ�E��y��:(�1��e���>�$Ђ�{�G1�p>�M��j���~�H�/���/��T��/�&�a���%�	�=�n�h�y�M�**I�n/�h	 �d��vχ_B�]��Xx#d~����fқ�/'���{�#yު��n^����>�:!���0"�f����7�ݫ�mm����򿶪��G�Z��&d���đ�ƀW7�2l��C0�d�hXj��h���\.<�L��W�������V���mj����[[����o6�u_w���_௺�W���/��/�s������[���@F�^䞔����d�\LP>�U�Th�Gy�':�PU��?c�� BM���}�G�8�@��}��� ���m��~\P�'11����!<�փ��S�����UPU����}���Dy�2������ޟ�m�ƪ��M�U�X���+6ը�F�h�Z������э��-�F֪6����j�5[b��[V�kX�V+ƵTmQ�X�-��Z-m��6Ѷ����V����Z�m��m�5E��k�Ij�m�mj�j�kh��F-k&����cmm�kU��+kƭEh��ŵZѶ�m��m�����6���Z�Z�cZ�[Xڪ5���[V-Uy��}������/�o����ӘftF�#�=={x<U���:r��������y��_�{u%�����y9�/���cX	/�d�ÌG���1@�3�*���b6(���PDA2�ּ��H"�4�E�
�1C0�S��I��H7����$�2���`*)!�"v��U�`S����@�  ���(��#�qliחAC�Gh�HK�LN�ʔB�6b�(`�-�<h����m �Ni�%��5����w$S�	
���0