BZh91AY&SY��r��k_�`xg����߰����   b<|  ��me�L��մh��J!P�j���l�5R�M$$%3i5f�6���hj��-kb��cQ�[4J�ʢZ6ضDF��5l��ã�e"�[F�ֶԈ(�)�� T�&h�jJ֙�R�l�(�ڪ����YD4�m@5Z̚F-�m�mi��X�U�6����Z�5�������5�&�ce�(bV6�Y�V��ªm�Պ#L�U�6�Y�S1��F�a���YZ��ƴ�m�Z�mR�Fl�[ l�L�Y�HՏ>���M�Kg� ��}V4Wq�꯱��j-��Ѣ�wC�z�OoO;z[Sufٻ���N�3��v�m��m��r��٪�SC�w6�P2ݔ�F��W�`�#U�cD�i���  {�����
V>��R�M��{���RPgU�.����O��
������_|�B���;��Ͻ}>�R�V]��B��^����t�"��>sN�)�ܶ}��B��mm���+"�Z��.� y��ԪT�:���AU��c���*T��{�=4zwiJ�%�U)R���y��J��;�{�UD�m<;{���T�;ݫ�z%T�%��z���i�W2͢V�f�L�Z�[&�� w|TWZ�^ynzT�*�z�zJ�)J��ëA�gw�;އL�R��y�����^�B����/z��R�c�sZT�5=����T�4�jR�R�m��E,m�{� �s瑩؊��ؽ�m�����{�*�jv3qL�U*T��ާZR�Is�gm�
U=���ҠJ�s���^�T�U�Cr@��U�xw�R�R�<�Ul��
����mcH���  ����HR��Qܪ
��m���R�t�.�wc��Q���UZ=:WzM�JV�Wz��T�JW;շ�Q
����*��积zIJ�ҫ��f��LV��jM�2#5�  �|�[eJ����R�HG}�]��
R�{�k��jJT���y�mJ�Ew�;���*Q{���K�*�����^�[2�JJܓ W@3�u�h�0kmfԓ5hA
6�[�  \��E]���� �x 
c2���\���U���Ż@���`={���oz ����wmz�y^�Y�JT�3i,j�m���  [���4�]Ըh������EW�-@:Uy��Ī+��p��tP{ۇ���w�����淞UF�Z�ѩ�U����4�j��   ��B��+��
�hR�=ޕ�ֵ@ޞ�� T�a�S����a�u����U���@u1N���       4�*J�C 	�     E=��R��D0#�F� �14dh�~&BR�M&  �4ɄS��R��� ɂ`F ��&
�(��F0�M2h�#&$�JPG�	�4�$�z�Ԟ�&���S�MI�?��?��`���V_Ŏ3���[��Sso�r�φ-�f3u��~�������U_�� {����~�խ[k���[o����*�m����n�տW�ߟ_�������|�������j��ٯ����[km�m6��j������gk_�Km~�Z�t�o�J����~�mkڛU�鶯�J���[~�[^��z��ꖯ�j�R��J��5ojj�T�ީk^�U�R��Sm^��^�o�koT�^���Tկjm��mk�+kn���u-m��j�ꖪ��m�[�6�m�֭ꚭk⚵z��kz�֭�R�m�T�j���Z��km[�-���խ�֭�k^���תZַ�[V��mV��V�W�j�o�kU��Vַ�mUn���T��ީ�սSV��R��oT�m�T���RڽR־��ީT���SV�R��R��SmoTֽSkz�Z�Mj�Mo�*ީV����6�TսR�^���T�������CH�8��I���������MeK�_<�a Bܱs͓*���5S�t�j��ĳ�Ō�Yr,����"��.sqᱴ���3yXh�M��VRk�j�����vgnuCm�Q[-�Mo)\���3+�A�Ƴ��u2�Q"��T�Ьqt�(�t�E�e])L�U-ډК�sA������řO@Q�oZ��,=�F��E��Y���QV��<c�j�wr��p#!�Ȉ�ު^�k�T:�����S���#�_HIS�4;d^e�&��Ә�-k��LP�*Bwp�Z��+���]�$mU��v�0�e譹Z�e[p
�{�7�i�4C��V���b�[������,m+����,�r�B۬��T�U�]���Nʫj��s�1t���hd��00��c/ �Q�n��E�Z���q�EI04�ء�F7y_Ljj���Ӳ�J�Xl=����YZh9�����A�v��n�ڙ�,��=�s�Ԩ�ܮ,�tp5/��K-��N)�}��7�/ ӵglQ�������� rVŽ��U2/jk��sT���mc;Z�YYd4�^bun���-�@���M���]�
���" G2��6�#¡��P:2SV��R&I�F��&C]��J�;ֳbYI��b�<N�[ͫ�'�\J�X��{�:���\��̨���`�d��)��Y�@��2�L��e�["ϰ����*����kq&��ː���]��w�fS���r�fL��fn�R����h5�0c�+`�U���K:��.�2�cǆc��	V�+%��n��8�h�"�0�W��,��+b]8����M�"͉���.�+w�J�ӏt�S��F�Q�&v)�,�x1��FY��Ԥ��GN\�T_$����R
�@D�]�wҵYe<�ѵ� �kN�[Lf��������u��L��6P�ֻ)�7b�M�1�:Tb]եm�^;u��<�ö�:YЪ�ww�k���J�}.�-� zƜ� aq�̽r�䙓+2H�1�{Wv�m�iMe�KM��3���P�9s����5k8#&��t���e�{D��2�&��]�V���n�N�y�if.����[�O7	�d�F�ؗQ�3�$3 ���{�@�W��J��ڛ�T���3�)I�յ�S"f�b�R/nd�P�h�M����`R�ym�ڶ���owq˨�VNkbR	�r�$N�?%�(M>rF�ˢ�����%�6ը&B!��v�Ou�ӊ�p�P��,��&Ҙ*�ְ��n���{E��j��ܒ���X�u�tȝ��`�&n���b�P7z&!�l�]�����q��4T�-����Q����؜0�S*�k*;��q��&l��J֣۬Ű��W\j�wҲ��Թ�t�YbQ�6�L�gjV�Z�n����H9O)������iN�V7y�֝�C"ib���ȪP$�.eh�c"T�Yh�I:��w���A���ݝ]NpE����e9�q��Й���*�cn�K�1�{�1>#���r���]RU��݁�PT#/,�U��4�u���`�w�������鱩 �3[�:�8)n�>���`��d�E�_il�-���q��|�T/�i�*5t�yV�s�h!Iiӗك�X
äo��z��ޖՔ���c�X�v&�6���,��"���fvޝg5*�c���+�(�y��w� /��-��x\�+-�D���~1Ơr�W@���s����4�L�	%�r�X���x�mY�9��t���&k޺r� ͛�K�7�J���e7�E�^	Yna"���i��ո�j3m��s���>��d���N��0nSUm��]VO�VH%��6࿴��M�8tc�:�:>�$ڬv��F֫d�m���D�s[E�X�ބ�,�#��x��Z5�eGN4���2^������V��&�\폵�Nu�x��;����{#�	�GsD���
�n��f$Y��Q�~2�l��5D	�?��ݤp�S6n;��i s{�db
�2�%�>'3)`Ux�F�$Q�A��/vF�LuΔݴ#�����'O侦s&�"ȫ�1�i<ț���޽MQ���τ��[���6�O�;db�ѐSJJ��U�Ʋ�+13��:�"�b@��]Nz�;4��9��9J���b.,��V�u�B������F�� Fͳ�ML��QX��ס��Z���(v�5��-&T�uk&��V��
�F��2$d�x+K/VwmN�μ1�`�E�g+DS�b���i�7��^�vE��
�X��C��-�V��˙�Ѣ�KX��H��RGj�h*���{iR��7,�m;�st�)�X궊��ˣO���'vh�*-��j:S�o�\TZ�q�3K�I&��	��Ppͭ�|r�VO3��!K�C�Gs��r�3 פ+Ǫ�(�'~H�j��םA�KQˮw�����E�q�H��)R׵h�X.��sS[�y#h��
���P�����>qٮ�c(k~rM�K�]���:��i?KnRN�!,��13�m�k���1i���dNm�m���Y��V4�:31mb`� �B�m�b爃��uu��QBW:[si]�����f-4�(�JT#V���n��e,�X�*�|*Mw��P��V�r"���,�$�uq��#�X&]��F�����~wn
l�����H��)m���q��Z����2�҅�i�36�eV��ؽ����0�HR�m�|VJ�4�MִK�ՋFJ L�{�Y�sa��`E�s�w-�uf�[�x�<���&�� �f�B[Īa(��n�DQ�ws��OBՖ)R�(��LS�*$,wf��7�ecz�VV�h��`�1왢�j�m%�k7�v��iW��k)��L:�Gv�K�_vލD��Z֕���F�If�ui����[+DVs%]cS�� 0+ ��s/�C��0^`Ǔi�#$j��y�������� OMC��u�;����C'+LH����7M�!V`,�Tp�=�;�=�V�� z]�����f��9t!Y����и�62�ڴj�D Zɣ���4�5@wVڀ"'kG�p<-�w	X@P*Wu��!���y�����@���[R�Ha"����K��P�k�؃xsh�x˶�Mc��͵�&��Ej�ZoP�ז���SQ��3��"���Zt��ohG)��`L&� 2�TV���^95s,��6�I�8w�lfҙoPض�qM$ǉ������,�ؚ�U�S"������X��8�dt�T���*��1�yBH�p.`��,e*[Q����6�Q�C(�H`=������8+y+�.���bJs6�J�;��/%��KGa	�7�n�|� j� ��/����n�du尳�PB��h�T�Vh
��wi��p���ܼ|�GmP4T=;�( B�k���v���0R�6�I�7�]�H�W���8�{�5ћ�R^�fV�����R���xں �HSV��9!�T�);8��<�Ơ!���w;R%:�6�捨�0�gGf��&SM2�gI�hn�(tsfQ�M�N��e�A2�o`�+)��C(f���<%+���5m��ݬWq��	��.��Z*�V6����)�T*�k@��NK�S�yB�SK +4�\����>M^��
�`+3��Y���O�-�v�7����:�s���{��8���������7��Y�ƓtYͧ���!������/_^ۡ��~7�h��V�����X�Y�q33Xo2�CՒ���@Ŷcۃ(�v[֖n�*̵6�>�j�TLx����.�e+1�
�����W�Xݢ�dp�ca�Vœ�9�I�E�����D�}A��4n�Df�0������v�5{���@ �6��v��1hG �9M�9(��a'J5�73iRͽN��7�3]�3�-f���p���}B�
�̐a��O솭���:j�4��s��Q�rYE�Z��i�5`�h�)�\\]<��^PT��	⣖��h��G�/���i�ې���7'� ��ak�[[N���Y�Qܵ��7��t�3f�u��Lm��V���Ӽ�W�9�-���2��9�Gd0a��u �u2 -�� T4��@ W׻L����3%;F������o��aWE����N���h!�����m���˯��V�[H�W�*�n���a���:uiG!(�"d�LQ��dä|�Lf�}/djr��H+)�mN���E[
�
�w��包e�Xgj�%!���>�v�˾�ӱm���v�9&��Z��ۥ6�'�&�Ty�z&X�7f�ߋ�L{(��U�Yt�����`(�Բ1��uF�����*��6yQRѭd[��굖~ȵ�&KeYV�+;>�'z��j�^�2�RW���Ԙ'�[z�d��mK4P�[������x��T$��B��+R���Cl�]�*�R�6a*�V�V���Һ��.u�)�[Ok����.�yc^U�F��TJ���wn1�Y��1ԃ ̷i�jTb�=%i7��B]h4�7r��1�-�F�!X���iP�Ԯ�ǶA�/w���m�n�;�Q��v&=�S!�(Z3k_�j��nth}N����� ֲ��j�jO6\5$na�d�f�5��i�suh�vƽ�g)�����nQ�Q�#��fMcv=ԅb�V�X^����H��/�3�[��9x0^�kI2�0�с��4�[gE(�0dH=�o6�q}vl���a	����Au{Q1�)�u�d��Si��hcz/j�ֶ
��ɠ�7DXT��cq�#
�^�6Σ/[R�S)S,\�&����:�ܤ���sT��L;ˠ�b�Õ��8n�xZ�#S��.-��W֜�ћ�K[5
`o �)�[������Zs�ۦ�I\�M3 5��ys�.�%wXr�m-��t`�\h��&h n6h�5�ꃗs>`�Tج�^ ��Bɼ���N#{�p뛀��~6�n��qj �캲c(<�R��X2c�5�cUb�(�8��Yop��/p�*ٔ鐩i�v�ufl��vE�U*;p4AۭH�/r�P��[�E*E*5[�Mݼ巕��:;�+��v�OI\kM]��P݅���C��E���>[4�	4N��ܒ���o���,E����m�]eX�	);�]&���]^
q�sL�@!������
�����g>�]a�F�*�/(�:K[�ys1m�M֍M$��tf���Vwn�	*Ʃ����޹��S!c�(���ٷ6f��ѫ7�i��� PX��T�nV6�#�w�bԊ�J��U�P
f
�W{řE �lϯ]�7�l&) pVI2�B������ˋa�a�n�*n��2�3y.�LЩ�`���ת��Ǡn7��W
D�����#.�"~�)ZX�D0�t��IW�&������z;3(� *6���B՟�H�}�6��*�X�Ř~�m]Y���7]3`T��巁��9C>(�%G�V 
�틉Jj�R�!�x��)^J[��0̂��D���F��*a؂n�)�ػ�^C�|��B��d<2�̽e,Z�G3D��y��y[���φ��N�T�s�w��11�wV�,^U�N�;�U:˛�{#��U�歉`p[��yt�B�	w&� �f�e�%0��s��<����Z���xQF��4L��
U�f]<X�w#RnJ'QcɊ��6�֔��6(էDiٕ�n[M9��jHY�l�ޛ�.�"�d���sr�ُ&�b�cp��[TIbj�cj���k�Z��>��[l,�-��*ݶ�z�R�0��eMȦ�Oh�]^�`T�F+.�S���Z��ו��&�\ he�*	F��F��KZ5z��	���)�wu��h���/x��CV;:��MۭV�7YL�iM�n�jջ�/kl�'aQ`,�m��7c�U�f���TL��ff�2�E�Y��)fe�ՂQm�p�B�����P�blV��=U`�pf:4��p�(��V�L��p`�ӗ*-�.�"����-L�,�;�ؚG#"��v�.����۳��MXkr`��,�u,�+3�$�=k��"�����e��gwW�5e�ɨv�;OS��N�>����4����}h���o�,�خV�L^��n�VR��X�N����$�,�	)E��k���l��#Twf�v.JB��D�Q�V��Ї���0|��n�������"�(e	�����P�]ޑ�3�i��r�ȝ����J�KB)z�wY���iݴ&��3�z�/+l�P�k"ٽ���F�j�u���\oE�J���݁丞m�u�f�u��GNK&�,jX mH�@�07� �J�v��b���vݸkk	�;Be�@�/��8�L� V�ν51��F7�l�׮��(�_$�,���L�#Gf%ua�1��%\��)8�c3Z��)� ��`��Ү�b����s�X��U�].�*3��b����*ka�9TeZ�r��8����X˧���6��dc������U�u}��]c�7�	�9�����A��Zk2�z�V8D��e2E=���HL�˔��֏����%S�	���S�v4�:���7�G�س�نֳ�>��ޔB��v�������*�M����A�Mc<ohq\0u'���(�R̦�!�+4ֲ2��F�y@J
۠���M�/�(j��(VCG�5]
hd#A����mҐ)�n��C��U��Dkc��4h��|�\(8A��4�?3�eA�[���c5t)�)��X2���px�'V��e1���V��Ҫ�L7;�<m��nh�������yqK���E����/�W��zn�^:�Ҥ�xQ'/R{�-�e>nT[�[����Q����?����_�޿b�����I$�I*I$��9��֜�H��$�G*I$�IRI$�˒I$R	$�t�$�M�C*G�����$�I��Nezhs�	����8��b�� �emu�T)�C]]
��o��Ы��]Q�pB,ۗmT=z�(W)��Sb��=�&���MGΛ���iP��W�ci\wˡ�Ԏ��j;��C)���3����#�a~�Y	����nZ{��Ƞ�t�y�5�*P�Z5b��حP�H�c	�E�wRn�[6�ޅ��K�:��b�-%l"fa��rWIN��ы���hh{��3f>�L+n�6�|;�%�h�Sw�#p=�oo���Q�k�u�d�q#V�%Qk6�;�uk������|@6��<=d�O/~�2,���d��	B#]�ά�b��aR�J�f�B�sXϲ��^�Q��/l亅o�����%6H�6��*�_�V����2&�P�f� X�{9_K�r�k��"�9H�]v3���}.��Ã!;�bPf«�����ۙ��o$|��e�-�C/�$JWU��O� ��>�=�ײ�VŲ�!R��vL���n#�;��[��Qu`����q5!t؜���W���+��k�Q������LR������'����u��ui]2�����Φj]M:
)�U�P9�Z�6mփ�%ӑ_<�����ր��q�����_W;H�9S�f%����3��̮ȉ5��|"������<j�A��RX7tT��)�^vޞ�**t�TMή�7#��S���̢�	J�q5ow��-�"�P��[M{��*5��$�ս��Ws5�ݢ.�;-I�Ē�yT���z����0��Ս��NV驍%бK��!²�=|a��m�L�xh���Ϫl�F�U��/���y��l,Է�d�3��7R����"0�s;C)�����%8;Fn��H������i�c]sf�b��X�j�����\�-#e3�j9H�U}M-�XU������}�����qˁf
ϑZ��[ݜ�lc��ٓ�ݺ�`,0C@k5GI�C�:-����g*N��&i(�2�nʽ�� ��*V���5fTǣ1QKH>��R��MCԦ82v�S��.�T��#�n��C��0�Y�k+�*��o<X8���7q|uI�\-^�ţ\�	��뫰M6���v�Em�mYY���ѩ�t�{�U���C9�G"np
�#{Æ�=�;B�9�%th0��̎��*�h���� QV&��̽��LH�,��O%1w0�u��C�AN�)��_�ˏ0�M�-�֖c�c�)6�tNR+&S��Z�v�Rb��F�o��
�7ېy/�P��ỵ�"m��^V�YR,]E��#�)��/�L��� ���.Wa��ֹ�Kһ�J���Zh[��as;���@��R�sN��_f�O�#O��C�S�%�;ax�;�&>CI@�I<*��kK��k�r9t�Yr�������"m����y�Ƿܯ��c���n�����n�>�^�>�8ܜ�ˍyB��m�0K��Y.����,u�N+�7t�h5�����6q	�Q�����3��������j�hk��/�9��o_?P)֣��Lm��9�4�^�����al�58-�9�B���:���Im�'RY�:��<���U�"o�au�O�_Z}/�ާi�>n�f�^�ڶ�`�z�m��`#�2}ңK*�kNgWZ����9A1�j�x��V��g*n�tr�)������[�=Zuܷx�K�g0G�J��,���.������U>�^��N�V�PWWT�d�[z�ve
�y�r�r�Mf��
�ͥT�2n�y��}m�Y3�V���S���j<�u�X��aD�I���M��J�[y�pi��{h�a|V:�A����u�F�X��u�De)]:��ah�Mڗ��;j�u���Nw�of�/*Je������a�w�)R����ͷ�;D+��I��'Y�N��y���cQ�ug��9���:��њ-,��.f`bnQ#j��g+q��B>{�u�T��|�-!)��$]E����W�bo�b�ĸ������-��,�z�-��� ���q��D3&�7r]���|E�ǽ�X��_�k�T��Uuϴ�8Xʌcm�B�]j�T���m��h;E�6L@PwZ�2i�ݑ�v�hʘ���_/��im̐��`<�[qU��-DT5�D���3Z�Yot!Ckm�Y2e��x-c��k��׍�?_]-.��*v���n�:����wtM�ʲ��1������X���r辝Ę�)�X�'4�� �_lT8Ԉ\43��-`��E �5i��^m�a�6GQW��WVn��r�up7SzS�
�49��#t��JvU��u��gt����g��d�ܐd�ɽ�M���u+�9������ꗩ��`j�,�p8���i�S��Ɓ�)<圶���/�I�A-��A�}%�X��oM���@2�2�KzYW��u8��^ޜo-2�k�l�_F%d1�(�N&�J� �qu����ki^��<�K}�	3/�ͮ��I�w[��`�ND!��u�[.��uޝKn�`[�c�!*Iq��ʹ)����&����	ޔ�;�f��ds�÷�f�QJ�`�.�s�ʈ*U�̶�r�y��;��E�����W]
�"+�[��
�V����IBw�.Zzsy��޸�7XĦ�	YL˱�Ӡ��Rf;�{������I��a������Z(5C>W�S�f���f�̒�d��n���_��k�'��c���ү �,�nJ��H��Bh�V�nz�IeC�*gtޤUs�n���+���IN�S���>�]	+���#F�(��Z�}�9�y@� -���u�ϱ�d�wΦo.Bͩ���I��]J��-����bLM���|ވ��cM�[y�w�R�q�V��	�
�OX�Ui^ ���P�^>$D,H�N/��G�c�Ȫ���vȀ��I?��x��q�u��+�Ah�St�Ӈ�n�+�H�SWu��8�����%��[�-�f]l2Ha�[{���o��_v���C��5�+4��(V+��1|kvDP�Θ��8�t�n�>��Ui(&�9����
sIr��W��;��������n2���n��x�'F�NO<j /\
�0_V�i�]i��5�74�5!���9��1�t��Ū,:����,�wu�_�b�S9��ڣ�WG8��,!�+r�
�z�<e���
��ި�z��vS��wQ��4%l��t��:.�p��������Ƿ�7Jj�ք�H�$��%�H́}�ekN&�A�QlW����A�tsҲL��r�16��h)�_�[���\���)V��i���h�v�u��"�����5���+�-g;�K��x�'��򢸛�" h��kվ�u��4�Xy���	�,]��;�r�Wq�9��A�KE��(Ӹn����[;�lTdY������2FM:�l��4(�R���e>��GQ�=���Ŵ8�l\U�B�R���/,z�JyE-�Nޮ�iȥI��j����/m0�{��3�3��geL�EjӦ@I�(s�z�9�)�g�2��2��k�}Wj䘷5��:��14>��2q��9$�i���X��%m邅��{�U��B�N�T�.��!�i�N�[� #�R/����{)P�6�$Ko鄬3p_{uk��.��!���u�t�)ޱ����}�9�a�-K%���f<�%�mc��ia;�gkh�MS��[*�n��RXR6)�|}=�|�['=MǧP�O�<])W]s��s�ε�1�&�=��3h�bΧ�ر�PݴJ��@஑�X��7x ��Z��Z�t��`�Q�݄>	8pƯ�W\��P���7]�;�����J^dܙה�X⇰�i=��M���wڅ�ٴI ��e����up�1�s:@�|����6.z��7��qm�y��&6.���Kz�u���N��i��~ ��vQX�͖��g=O0\N�N襽S����o`yA
|�����v[6D��f��S��m#*�.(k��%��Y���Ƿ[7f�P�_i"����%���ø1��Q������jW���[�K)n�)S@��u7���q'#�;9ݒ�o=(7�`��J,W]8��9n%�R[w�Oj�^c/���<�:��KYJ�՞�Ԍ�,�ۖ�M����oq�{��dB�f�m�T��q>$��{�r=q�����4Rѭ�YWɛ�f%��veM�Ӌ��fB��s8�������7G�f��ϵG�°
��S�A�a8����q�E$���|����J�h��܂]6t^�JoX5Ż��[	�y>L��Z[��z�l��]rg��~ǟ�s>K4��hnn	�/),��aL%ٷ�/_u\F�v��p	�W��l�5ӭiX��U"��j�#��{�m(T̘��B��vAo UqD��0�Hv�y#�"�������Pֶ ڈ��؎��B�`M��6&�It�w1]9�oL���1�c��#��r��b�O��Tq} �Bi�,vi��ˬt�v-]w,���yic��w�]��iW)%(�in��G5�u����9���Fru���#$D�dY���t��A'��6�Uζ�ձM;�ǚ_u��E&)���eNRTFh�\nu>a�n���I�h�f�.��0h)ټ�����',�����1��N�>
lf���^�OM"�����V�v����V�����f
5�L�l��f��;u�V�K���+���WFp��H�fQ�$Xꀣ� GVn�j��薕�(V���Ͳ���`�r,؀ɼ�̇�'����4�ڋM����@�6V'�����K�S��<l�v�R�� ���u��h�t��斖F���&��Q����X�]r� ������H�C�7W�����n�d+ʆ>3��N����OP�� �m}���V�&)��.��9+o��>����x��-�:;�moS���բ里�e'�]�(5��"���qt-�J��-b��tlګre�liV�*|���'�\�`k��1b��X��#e�g�f��m�	���}�sYʕ�j�J����+8�Q��&4-�W��s:n�����e�մ�����ؕ��J��^��"
�0u�	�>;.������Y ���x��mLX�\k�:��ڱ�u�.:�N�K�xn*o-Q�e��&�"����+3�WV��?�L���&6�J��P]Z'vVe�ѫ�R�Ɛ�r�b�¦����7z�����n�z�fR�l7/[�1Ch�w@Ѻր��;�m;4��eI�3+mf:����֠B�h]i����]��	�.����U�*U��B���윥���-�Ht n�3��ر�Їf���B :b���a}���f�J՝�F�ϴV�(�.�! ���`�H�	��3kgl.��C�{n���T]�v����t��⵸�T����]�g�.Q�@�)D�
�1�
�i=Y;n�ƻ�� Ye�Cnu3��0��7&��cy|7!4�TK�v��nm�ӎ�k�ݐ��fKS�r�t픠�l����Bt�|�8&V��r dvqm�b�M�}[q�,X���Tv�=�0ؚѾ�YI��uׂA����ID7k�]XtĶ���hG`����Pt˨�u\Z/!�;��R@<wM����XЊk�Ik	b��'t#��O��n�}F��W.6��QMvX�0s�zj�&���<H��ᣂ�r4D����֨��+�,1d�ݛJe�#,�u���M�k�ջu��=�O�ep޽f�ӝ����Sn�g`�ѫ�K4xђ�ceϺ�k��ĩ�!Xy�ƛ#s8+\�A>�ϖЎ����#ִ�=���r�!([�7�m>�V�ϛ�E+у�����ɠ��@*��}�){��d�Q����	]؆en��5������Fwp0B"���V{��%�����e-=&�[OOf���n�dӪX�.��]��9
,H�z�X����?br�0<�Vv���j8��g^�z]+`�$8bcx6�hV(�M˰l�M>v7\�c;Y�y1�A�n��W�S5,\����"������f<���k1�f�4�|�;f�^8�,���N��ٮ�-�o��*��j����[�d�񷺧��J�݌oos�hj��CU��p�ڂ�Et�:��V���������4E�sl.�%���oI��:Ĳ��D�"{�X㒄�cv]���p��+��WV��>�;N�E�'%�_��6y���nm=G'��[���3t��Y�@�ਞ�};yV]L�\��Kݻ��Z��&3��4���v`�	-6��g�D��� '�=�vWm$�,ԫ��]���@�z��=�X�lT�S��VK�c�yG�l^�:�[��.�P��|�����7IV��;��;B:f�Fr�����Uo�9�R���!�L^Vզ�Ng:C���K�Ų�5j���HŁWk'w��m'�xm*FH8�[wrn��7��5�;\y���!2�̧:��MJiu�R���{�GU�d�X�`c��m^n7/*��]Y�ء�� q���L*p�;x��϶�9|�6�l�GM�G�yWwf��n��k�q��lp�"�3E��d�����Z�vUm��p�Υ�G8*2ΎM�/�4�j	]�j\-�zӮ)��a���boj�$:�#��-_WT�Cu���b�%����O�8sbY���2F���I$�I*�g@�X:�I$�I%�ԡWVX��e �~ 3c�bb�n�h!���P4i�A�@a A+u��@� 0� HA �(�� !!�   �� HA � ��,xLҐ���yJ����j���+m�V���{Z�� >��N���?������@����������������{�~_�����5���La�g]���'gl�+X�a��"r�{�f�JF�T��H6��Z�a1���o*f+4����@i=�E�N�gZ!��)%�Y:T[HȺ�\��,t@]���E��j�h��Kp�O����d��0�X+U�IE�*��c�{��1\���b��;��I�Nٶ���ft�v`Z�{
	���Y\�n�6����Z���P}{�v��w+;�2��K��D��]X*Sdy(�F��.�u9��HZ�w���t㋑�v�"��d�Q4����i���s8�������^n]�G���G�]o#���NƜ�����g�7�4;�-qH,�=���P�����l�Z �o-���GsuL]l��ڜ��V!�d��wzv��"{��ͼzkH�p�C���nA�n>Uv/&�����J-S[���J{��fNǏ+1Ls��7s�!(=��v���Ԏ�w}���vaؔ�-mrȌ|$�V� d�1L����eK}a��!��OӥƩ��X�@:��}����)��u��̂	�n)k�G@f��{X����0��T���-w,�����/�����2핉��F����Ka��v��i*�:�;Y�r�:�;��%��+j��+��\�em��l�5q[�p�2n�H:����^���.+
3:SCp��^�V�-��CY�9�:��.Gw����pI3�ܤ� _�3v���u���̇)��I�^�����vv��{'x�F�k�����@k�{Òli)-
�}
�VmK>�C�ҭ[����r���-EO0 ,���e���n�:�}U ��o�$$��|֒��Σ�N�R8T�ج}����mb0����9��<����2��7h�=}D]���J�x^2�9 �CV�cW��(���Xu�۳{��g`���!��٠؁gr[����9k;&�׈,���=:@��O9>OS{Q�a�\j1{u�a��mQ躷U�eֻz��*��Mۈ�:�k�Vk
u��6�k��[��+z%%n�J�9��`氏X;Nl)h)����Xze�&��cWC{��`v%��I@�ܨ2[�R�r+\��ⴤ�M�4�]���ZZ-��o�+(SahP�骮�Du�J��c���9qj(�y��u���-��`[[����f��#�ν�V�>u���U����)��ΎMٜ��nw|�&������i�z����r���=SV:r�Y�C�A�=���v��X�1yh��PF�8��-|hj�YMd����� ���,0���WV5�y��87/Y2Q�YHhb�o\�*�p�^��ݫe��(5d�d��V��*��x�qi�����]-��x�wp�L4����1FU�qRT�� f*��8c�v�WM܀���f>M���vi[���9j�U�����G6���e�
˜��|���V֜���Tū4/��'u�;���Đ�v0mJ\��B�S��9I�_8f�'�x�)2��s���i��3T��1�#l^ݱ`�۹���&�>U�=k2�O,�1�˨�M���8]d4vMjҵ�C�j��nݮ֮L�1��oS��&�w9q�yJ�Y�ru��V����`t&˗�i+ޏf�� ��ً��h�yI����T��sEP7QJڛ�Q��ܥp�Y�.�X�il�v�U��n��u�_Pg�$�Y����凷&v�[aHf:ͥ�Z���(�T��
Q�\ Sc(��cM�{�w��.�R�:'�Ѥ��V�w�M-��;�e��J�k$.�91KȠ�E�lwa�F&�p�#��*Wb](�"��6:��u,����,I�5n��x;2:��z�U�
ő&"������n���h�Q���h��q<0й�$j��D��0�]'���T����.F�_tӕܬ�1C,��L���ReYL7t`�]f>����e���qv$T�,AF� �CP9+63�aM���,s"{[��1N�꧴;x��ƵpںVlΧޙ���H�V�ك�^Ik58uY��F�s��.�b���9�PZ2a��f齶,�7�6�:.TͧYo Ś9\�;��S��(���htAS1H������#�B��'L�g:S��6Z�#�N��QʸH)��SH�fS��t�<�D(�������ct�I��%f&�v�k9�
�J�l#8:pu�n�aVڌ,������ҷ��3��Ā�R��#�EH�d��X�0�fF9�V��ʱD�U��s�C3���KQ�g�ףt|���Қ���[���Ng���(�9ڕw�$7º�c�c5��eZz��:u�7�}\9������<(Q�|^ b��3��ԁ/&V��[9�cyݛ�`��B3Kr��������n�-���4����O��P�`�ƞ��3r�L�p� 0�d��P�t#4�G;�~�#���t99�1�4
ݘ��8mY� &L�*��{�pY�dٛYᚫl>�jQB��8�Gpt�}˛�u�jP�Mʖ�De�gn����d��F��fꓢ5�~&�f�C"� b�-Νh���5��(0\=��f;���i�����	c[��T�Sw��'Wi1�6d�� ь��4�*��.�9�1�M�S8��e�&�s̭��H��+d[��l�BC���6Rr��wn������L�Cqo�������^wf��:GJ�}Ru�ȝF����=�M�ܘ��c��C+��$ػ~��'V��˽��,ΫJ���bQ*$�ٶk3��S]��L��s����rT�p+:�q��1���l�q�V��nj�Zg1���Ju��雑ЈM�3��^�V��. ;��G8�M[����d��d��9��&���Y��V�[D�d�ɶ��)-��N$����M�sB�tԭ�m[��ˮ�k�&l�oh��vl΂�g2�5*�5�v�j��3��9y��6��F:6��݉�_6iP���I����.�a�fW#�D=���������"���h��V\��h/�����]dc���jg`��̣CZѣyVt5���g�)v�Y[óL�}��6E�tɦWp��4���&@6���<7\n�Ǳ`�ڔX����q�V��r���NV����3h.��R�� ܕ��+�P�y6�߭,��Z����E���.-r�<�x��#2���χm�o%�N��4S��N9�M�d���v�IY��nj\hC�rQ;ʔܭπ|n��u���}3dN�0]2\���"�H�	�ҜS&�FOr3�w{�R
�C��Y�r���=��Җ)���J�!�n"'v�;�q;#C9|�ch���@���үb�9��C8�ز���G�����R��H佭1Q����:��6�{�{�W��3�{��k�P7n�Ukꗆ�o�!�^.0EL<�k�s�J�������.Qw�7 ��eE\��z�7q�O7gL�q�j�����YF�LMҒ�r�TZsF���!�D���ë�\��n��OM}�T��˓ϊ��YW.7.��)N��f�y����Ӧ�������K�Q �a�֏�Pi���v��r�iGBIJ�n��OI#1c�2�������ƾ��+��+��,o5̦�
8�>���}��^1Zv�������P
1ʵ@�N.�9-\�\���kB'��:��Հl��"p=�ܬm�ݗ4,�uڜ짱�U7t�2��4�t�Rޕ`�7�.�hW.�#n��zK�wbiY�S�;Z��L/�n���5eX�湯`�RNӉ�>��nB��c�$�"zff��hO����8���oM���IR�/F�㭾�N���թ���k�P�[���kձ��Ֆx����̖o�_c�4�	Xi���(t#!ثy^ͧW���^�����uh�"�]*4UH>V��|���jn�;�Yr�z��7$0R�ŵ��M�QϷ�%��s�ڎm�t� ޻�K��y��;V#S���k�EKE����I�Vi�ޗ�ou�<�wn4c���-T���m�V|�o@ܭ@�W�eGΠ���V����o��6�$�i31��l9Q���U;Z��B %
G��s.�k�fWbI%���\x6e�N��\��5n��/0 B�c�3=�2+jmN�oOln�\[jCwq�k�X6NgX�{�z��-Y���ˡ���/�V<�T�ςx.��cv�{�]m^!�&՘�u
��tЩWʵ|HSD�m�������ח+�_	]2 ,F���ffmͥ���v]V������U�i�c��Aɋ���LJ-��V�}t�X��|ŀ�\S6ip��[@X��T��>����dn�G=�i��'\��M#;]Ф��(f�1L��m�� �\րF�U������cA�]���1WU8��ʛY�ȩ�3��A�{@>��yd���W=���^mY b�9�җ3Q�h�u�<u&i�M��C�kEr=��>˪Y]R�.�#}5;M�e
�;Ojhјv�i�6�#�M�6���u�B��hÕ\���ՒS�Tl��̋+2k����
��z�t�ڥ�]�#��E6��X+nnq���o�;��{�**Z�Q���n*9��
�W>��Ys��e\"N���+&����F,IU�t�r�o:۰H6�ǳ5=�A�5�okW+n�0탸fYNY��۵�&�eA]X���:^ \�z{ Oy#ّΥ����[����	7m۰�z0.皱�ph���;�@V�ʣ��l�*���"���(�{�⑭����Ǘo�;�x������skg]M�o�tɷt�i}�&qފK[�ec�c����N����	k#�	����mf�)�W|�њC!�{�R�78��]I����ȳ���ZU��.`��3r;�!�Jб7s	�&�=�u�gO�f]�Yz��:��R�k�V�lu�����U���*r��,�Q��Z�;Q8)\Ŏ�pV^E+k���WUD�i��ȷs���%�0�iʨ���ɣ�KrWt�"
�U{�@��ն�7�۴��)�5W��;/�8+�ɦ`ٮ�c�i�I>�_M�0n^t�U���b;�2��6�/�l�7�����ܸGݬ�`>C���*��S�x��nP���Rx:��H�{v+�l�K���r��gh��[��� �79M�,"9��P�<�������X�e�[I]m_kDg7BS+E��eһ�3���Vxݘ��f��IC=�
E�����i�J��*l���o���8Ҏ��+���-}AA��e��3z��ڎ�Z�S<H��\�	/m�&��>}Փ�U���:(� �M�
eY��s�҃�����k+u�y����k�£9�,=��_8��Ǚ]:�V�+&YƖ:�p�``3�W�fnݵ�U�U� �{3l�,k�q+�X��Mp�����T��2�Z�ڌ&�A]��*�1���_K��'q)��!���+2�ԕ����l�I �"v:�y�X
�r��{�vV��T��%Rl��9ŷ�/�;4R�Cp��MbX۾�5D��g���nBk:�Z����p=����X��w�b�LǬ�N�W�+ "ht�̺�k5���3S�5v��)H��}Y�u���w��}&��D����M*V�kue3�@�+���3͜VTn��wX�G�*�j��$B�"h��^�J�l����Qd��c�`�����(5%ck���Aج *j=��zv:6��W]*�[\�lM�����0IV�@9,<���ь+	ܬ:Ⱥ�'����Ӓ��*�b��B�IN�V]8� 9��%4�awS&���j-��ft�Ӯ�n���[�G>5�MX�hi�[	� x�;��j����*Sh�S�����ww)ƅ�@��.?�R�l���b�7�G�=q��Pvfc��+R�`�Z�|Fβnog�­����f����6{�5{J=-ҬkV�<����2����:��*}}N�v���ј�&�rjO;��6�y�Vc�*��c�X{
��n�af��_ee�P�Z����`���+ N���V�KB��<�v3�:D���t��&���r�@Y�r�ш�n�2l�;L�Hf�)�<GU�71o���V�[��~E�Np.v���0��έۛ5��!�����[V�4���|\R]�}:�4��4�F]+Yr�7sn���c��lpN�3bDnQ�wYr�k]���$fȦ�\K�����[�}aH6�
Q<p}����):](���joU���رᕌ	Xf��@�7�3i_?�͊�L���ِ����O6�@���<�F$�ٸ��b=��p��-�1'y�'Y���V�ٹ8���wې��̈��E��S���ԫtu�G:e^S쬋*l���JD��S���Xv��Nw<mq��
�)�������c����ܹ�<x�>���R4�@�7���R��3#Ie��6Y�Ҥr�����'J���ح��%�&�i����:ѣ��L�'�j��<�U� �٭��\�ˡ��t�m��*ˍ�3wh	�X����2u�|k��#/��R�/�]n��U7��x���bu��|�+��8X�5�tάa�岩�X5�:�2�+N�-����b�Oj�4���G�SW&�r�e�]^�0c"�=T*�ܥ�����6d�՛�;͞�m�����VKhj#Cv�k+w��g'V5^�׼�a�uݒ2Yۖ��'¦���k���D��+{T�y��yR5M_G���@,��]��:4�O�ޚ�pՏ�Z�d�$&��n����[�[�:gE��Iǔ�H+�Y���,�ـ�J�E�c-3�\
�MLMn�e7���(���	u;����/�}�����i����?������+�
���+�ʿ������������_�u׽�u���	A��~�T7������n+����mÇe񇹺�i�ک��˥�E��$h��7M�4C\��l�b
��:.���]bh�S�E*���7���ǫJ����-��բ�e�˭M�֞�yH\b2���x�C��L>��U-�t4�iQW�j��W�1��ۧ#	���Y�r�M�Dh9={t��su2�4����.]v��G��p�iv�p%HЧr�Š*-�cs&H�ƵɌ�穁9:��J���G�<i�+cr�%1�&�P��eh5w91�� ˗[FL��+��I���ӫ�n�dX�f���9D�u]@ �L��Vn��]%ѢT�LP;�م�6�Z�f<cc��}��[:=� ��$;gb��d��ڮ�R�X�^=ې����:uM彿eKoF��|laA�2�H�?��e��*HQ�����.���e�S �V�5�N=�\�ā�|�\o%�kc&�|F�si�؆R૟Z�w����-=D��B��P�#��-haTDoA2�E����[ϕ�D��e���r�_<��l�&^���tVlM���kZ�N�](���r�8�\^��e�Wp[�kz���S�Ό�!{fY K#��"NR�)�xYT�h�䅸>�lP���hI7���,Z+���a��&Pm-��%]�P��{K�.�Iu�t��k���%�{��{�蘈"������p4O�n�
󸋻���:��u�t�x�i��u���qI3F��h��w"�e!Ia))&)�4�wDj(Hah�ݣ$�BE�3	��cL��*f0K��������IBC�����\eY,���P�[�#0�K�<�a*(�ٔ����I����ȏ*M0�*��RRM7wP�$�Q)��&�&	��h��0F+[�b�#&�@����I ��>����k ��ɦ��7���o�x�U��EX�h�]��B�
8�eAcN,!*��P!����T�9Z�?�{�	��T�@Ǣ�7_B3�����oo�X��*G���w5��z���'^�ҽ�o��O!=�?�eR�!���������5�����f���;dv�q��qƺ������:[�����W	�p�b��P�CŪ7��_���{,'���q%ލ�v�{��TV�?Vk�U�f���;��P�|s�g���e��s'�5�l��IQ3s��[}=��=��C�f篃�)I{{��嗌y5s�y��r����� d�^{k�M�f�6��g�<�ȝgĪ�Ӷ�g�/C��W�a���f� 2y�|$��9�m���U�Y��Ľ,��rS�"�����Ӊr�U�}V�x�c]��E��l�{ڦ��$�����&�{��yo��b�V'���_���1;*����^$U9�&d��i@#��:���.s��לm�{l�UU��KެNp��hG"����9��u{�r��f�P^`t�׉�t����unb�2@���i�aʹ��'&ΔMf�Δ8Vq��\�@��U���h�\�G}�r�Hm �WO�b��� ����_�`B�˥��YWT�g-�e�o��~��4��FQ=&�=��Ʊ �l����R�&|)W���+�W{�P+���z�xO�Om���>'�H1$t��f�܊���=�vz���k��o9+^�׹�Xͼ��<u�C'�E�h��K��rܙ|f\��_���L����Ry��k)a4����ާ	�"�?h�y������w㡷퍾�k�1�[7�݅�֩�O�5z�u%,���3�YtVw�Ϋ~�=�����q���˪2!����uW��;�ӾO<��^�vZ�\��rY�nzs�F%����ܷj�{�#~&���u�R=��o�T=;��b�V��?R`��Mݐ:	ڳ=�;''�]P�w�^�cS�Pމ��]�w7ydO?I��g�ˏm��{4��6�H7Y;�m��o�+(O�d�򧻣�L�3�"k�:���K��s+B/�{���=��dc/�.�*~(.��Y�zf��=�I�5��չD�O�/׺��lwd�c��4�swgu���b0F�H���p�����]�bv�7��e-���H�3�5tRT��6���
|ŧ�GPzz�/=y�����Κi��/&L�����3gE)�1�Ҳ���x-�Z�M�5z�����1q��V8�5ח��Z�=U�V�P���G*������[7���s��kg��x��Zlj�=��Ԅ����Q��z�-�%��[΁��� �IL��^��3_��=s|��p���S�<�J�٪�鏦�a�8V��N̿Q;^(O9�1�%��ٿw��yk�z�y��j�J�ď�ne��9�a�u#"����}Y^p�w{+�����蟱��NϽ�Ƙ�S)�X�w޾�J��t��c梨���?4�m��nv��_�&��p�nڧ�rt�M�~��;.�ʚ_˱|S�:�Q�����>�z�V����	��������w�X�a,T3;خ;���Y�����R�J����X>8�+��fD��Vb�~��L4!Y\J�<_���M�������ٵ�V�Y�]�\���P��K���Z�JRջ[�n˓����	E<�'g�Va�.Tvi�:�7Fș�&<���e����jC��̵"��n��6�7$�.��l�|����slxX�3�=�L���r�������Ƨz�99@�L���,t]߇1!�݂�NQ)E����Սo� ���]Nu�9^�'��$�Y;{f|3*��}�~��K<��`8��sד�4�)Y[(-�\�$73�^���Z��y{b�Pz�{y�A7�`\^��hH��D=^ܩ�)��Oޛs=�w�����q�eOʑz`����f��L=�kA��{o�ջu�������6p�9�
���j�&5�{��j�}�Oq�5�>�K��{��ny�u��:x.>�p��N�nf����A�D�|ڸ���eh��3}��-��@�N]��kS���Kk��{��S�^��j|�PTv��W!75�7m^�$�.C���Zsf"Ɉ�����9a��<<��/�4��d��ս8n_;��~�P�kf꺾��I`m7�ҭ}�g4Y��R��/��]_v3�[f*���͗17�˼�ǅ����H��$�-	��qW�@��2��pv*������]�<I˷8�M�cf�)��m��K�����~=���t���B��.-����~��Q�D�[±��i�?c�?\q���xⶵ���+����#�W�En�F��VxV:�,��{P��~��u��f�U��e�^]�0�.�$/�鵑ͳ6����tY��N�Uuh�k��zU�g�·_l�J��݇|�p�:�8Ƞ0��v�ʡ8N����Sz�u�b���f �a'zF�uMY�$���EO�۴�����#'e�-������O�u��u�1��A�5iٵ�ڋ��>�I婝�ބĹ�^<qo[Y�?m��x>�u���#���X�ox��rNP��qd��q7Βě��3��r��o*l��P�7�m<�j��y��:_�;g���nm ^��s������*��9��1-{��Q��ж�V~��$��۷]��r&�3۷ƲE��{S�PK6G��G'���,\-�n�.;*v!��u��7㣽^t~x+;�Đ���/��FmI���\3tk�/h��ִQ�;��]�!��pJ9�^�~٠lŲ�9�����7��f�ܗ�JY�;�
$���fWnG����(f�2Vs�����kww������}����b�戯{���k�P箁�˵�<���5m.������b�v{)��k�Ry�|$���y�g����a��Vk�z��p�.2�׾��0�fؘ�g���%��wNXs}�f>i�z+bv�D/{B��7e�� �՜U��ߟ����޿\�ǣ�"�O6�S�Wx�+oƧ�`Bܺ^���v{��^�{�bcg+aO:ѵ��F��lv�͐��O�.��������j��eZ���L�7��X�|[so�rF�� f��`�\�e\<713��5��7�;�a�Tq2,Z����w-n�x�P&K[�����W��b/kG&����[�16k{w�Z��M9g~�z�|�S+�E��r��l��i�$�<��8W��p9t#ܾ�L��d����3�S{Ғ ��u�4�����Q�c2��]ڜa�գ�6�����|��8��?t✭������{7ܶ��ݮ�/X�.�� 	z��Z*��OQ���M�#���5��f��[R�Yr�����+�\��Ӌ����F�������&)82����`w5-2�W�k��'��z��
��[a�ꌈw�����3ƻ?,g�N�����*����G_�w����NP&�Ӽ���(s���Oybۿs�-~���vWo�b;A;�d�����q���cR8ދ榝�^�������k:�u���i�CUs=�*xy�^z��/��#Շ>�o���w4�_��3��xr�UV�\��f��9� �����������q�1��H����v��(M����V��KX�\��ڞ�5৽y�}��9y���E$����D������oo$C��N@��yTl,�����^&�Z�����thFc�M?�v�o^��y�Փ�=>��}�>�S����o����zi����S�<�u�;��Kݗh�O��hz��/Q��+*���}]g'���Y��1��_���`�-٘��k��0��;�YE��+�T�m��z��D�p�� 8�s(V�M�ޙ�f_T���Y<�8N�(�&*y�l�l����G�<'���	�DU8�ۏ��P֏P�Si�=�k]���E���΁��Au�ΗC�ݘ-1\��y�J���be���u�ɨT�O�7�j���=TsU���ޝ��Շ��m @��F$�Ǡ��0h�~jL���c2��V�ʀ��Ƹ�y���ʓǫ�4���Oj��4��Lـ�I���Ucc��˧����߼����^K�7���Ȕ���=���J�p�Hٷg�]�"���m5�<�[�2Q���Ӎ��{��KSV�ܺ�Sp\�}����1�x���}����uM�M�U�Y϶o�3���]!��E⎃�-��F��;�7xNN����3϶X솒�ݎ
��͘蓼Ko����ZuM�;J�����r��������{�b�y-{r�>g��	/mY�Z.�2�Gz��wSt�	=�r�1��Y圇1a7����������_vP~�?VJ�Y�/���v�`��W�H��giɘ���zU�q.�N��tEV��;({����qz���u�CC���N������S&�����C,���u��;��k
Ym�k ��U4�h�5ա�R����.8��]�-.�P
M*�͗V��O~�q�n�̔uh,7B�݁�޸�%��;��'J|�I���7�!�ʱ=��͞��>����V����1�)?M�>�z�O|�o��B�et��ǻM��`"[8`�5����������A,N�z�19��ߋ���Wy�5^��j��4�[lϜ���nwN��g�(9׭СB���̒c>A���'��G�{��{"�/Ri�Gȋ�lǕh߳�4��kB��cr��95w��.���:3��!��~>��zfެw��-�,V�)�ïd �ӑ6�կ�\���١P$�w��2�_z�+5^�Ү���t|��3�4'�9�s��M}R�e���xܷ�-"�Æ$a$p$Y�zA���6}S��7n����x���xb���w��_=�=I}��ν��s�j��qsy��[������a��}e�� �-�~*����^˯ggy�+=�L�F�)�y��+�*b\��!I"3g]�yP���b��c��~�n�+�kw�[t{�EcF���g�>3#Hq�3v�B��Gv��7��m"W���"n��U��'�;/-�J�a�̽60��SU1�Ũ�� 7�$2>k�}B:�8ҫ�[��_tU}3��0�t`���ϯw>���oOޞ���g��=R:�}�r�>�ZS��N�W��r%~��.t%���*}]>��uN��u9�x�b���,�\i�$�����������1.����Y��fτ����=�8�����n������ƶ���{��r����HyK�Ϩ�i�(�=2x�[[=O�����k��W�s~���ۓ��ׁ�fh�^�.�I�OF�1��x�SZ#�}ᛮ@6���m�\]+σ;�����yH_Tީ����V\���%�mW�{r|suf�כU헑2H���?��c�*&�\���?W_�)W���V�6�c��\x]��^ް��"�{����YQ�U��^���⏥m��O��m��^��E\|�`�<l,^��/ё�A�w��ϗW�����U�䆯����|fr9���G���p�4 �`p��6��~,Sͫ�&�A���:�4|��[��F�X�=°^JX��#���{p����Ǚ�3�N��i�R�͒��r����g*�0:�#]@8�ira�̽Œ�m��:�V�Q���U�r� )㷲�����5�^��aT��x��# �7��:�t�Yץ�\�e�h�:˧��<��^���y]Z"�m��،�[`�L/��N���5n�6f��!L0gp��Wfb�J(�8�G�;�ŭ�E�g3�Flh>���BМ��U�x;""����1ց/]��czpdl�I��j�6M�;�6i.KZ��F�v0M�_�-�-��̤���p��v��q�B�ᆐ��F����m��H�U��˵�o\o���<�w[��Ùw� ŴV�����l*J:��'vv��Hjύo] �K*��[ՙ+��d�8����:��7^��K�Y�HㇷW5�bup�p_err��kw���Y����YW�/+y�K��5��J5jW/�۸��Qv�9ڻ0�����}�i�m �'GN�i�r���\�݉����X��6ԕLآ��%�o]����'T�=Ȳmv^���ZB��.s�;�Ԣ�2��{Hr�z2��U�̧z���Wl/��!��txr����5�V0� ���$
��V|�+�u�ELGQL��D��G-33+R�$K�BN}�v`�&sF�и�2�+T��ܭ�hWo07����*gS�Of�JgEj������ �P�Y��35[��&mdmdnȻ�����>��P�Ƽ¯�9繋�7K�ԷW+�5F�u�@�Ωn�@sp_$sP����J��S�dQ�zh�p��6�):���ޓD��\��ۏ���qեC{H�qR�b�e2�D(������S"ڵ��b�D�����wG\;��^���o6"Jۛ�l��r�ܬ���
iVqm��&\^��0�^
�-�{)r�tf�-�M4	�c����;�OF0>�J�����W�p��սV]�Wv=���3S���ȹ�Պ	�Ec��CV�N����z�E��V7se6ɼKNn��}\܋pB�e�n����b"�sɝ��\�o�m4��0Y5\2˧��j�XW��͢!!^j��AM��:��b�nU��5��1�Z�hŔ���ݱQ$�Aw�l͹hH��I������J`�jgen>!�t�u� Z��U��ׇ�������ݷ�V���d�%����m��,���5��{u�t@�xfN��M�C�Qξ��&���xU���C���=utf#h4�.��-��&�]r�miraQ޾�X7.�UcL��p�"齜�<���=�yR2\y(v�ή� X�1��
�yX�^\��l�f9Rs]e�O5Ô�z�Z0��7x���\���7QxR���x0.�Y�bl�t��r\͍�u��Ĳ��Ud-.�]�+��������F��j�V�8��$=���	�1jw�5����e]�u�f�L A�	���(N��R���܈� "S$��0�&;Rm2Jbd�E� Rl���2X,d�#L�����̢66�ѬhA�c,Q�F����Ѱ��Le���@�
H�T`�	F1�4P��%lm$lV�������)F�hъ#F@�9&58�A-���k���Q��e�ƌZKlRI���b��Ab�k���H���{���e5s[�����Jyv�`�FJ�cH�� H�������L����/�)�I/������/k
#n�j�1R��Y����w;��Wґſ*跺�ָ����=W�0c.1�]��;'2uP��s#[��F�z �CE5I�1a���@�u�l9��ɑ�N+UN�-���-�ϿcCEls}.0��ط�o憯������Qh1)���S�w��v��2�lns��^L����$�Gƙ��Z�Q��]ǹ���ڨm����J��Y����`�t��L{+a>�X�΍�-p]��EA��ΠkX�o~���W��]JT׫��K'���-�x(���\���+�ͮm��w�0�}��"$�{/P����q�L]H)�VU�1����n&j5S�:X0����7ǲ�5�q�䲋]�S�����.�w��cr�o��y�&���U^FL��q��K�&8/�P%�����5E'�["�h��{�T�>�k�)֏R��C�I�m%�]�}��w-����1�?�ߤx�/�qq�̪\�='�+�^�*�kq��u>��ݯ]�����zB�/���Q�ϳ������n�p��Q_wTxsYyr�1���.�oN��T�'�ٹ�
�b�An����Zɞ0��]�s�KEq�]!��)�NUt��MDv�z���|d��^�5^���拱�s%���#\�[�H�o-�7m��=+�=%�)���Ȁ�g��܎�7�b�Gc����nl�漠wh�ƥ���k�Ϻ���jn��y�`ipO*Q&uN���ab�vokWLM>S5���ב�����B��y}R�o��vB�>��4F_����'��r���#�Ub</�:�`��Žcnm��:�^´7q����	��/M��$*>T	��!�C��ܑ��W�Pgj/x�F���v�	�_xr��a���ӕ�>������`?������ͼ(D@yPZ��6�X�B�����zha���l_�Q�Gis'����#"ۤ
ai��!B�/�búj�v����Z�WL؝��i�|�>f!�;�_G46����P�c�z\��Lu<n;��j�������ls�t�y�7f[��7c���<����^�vv��kp���j	���s�^�J���HO+<�R�aORWro�.��?�2}W��+_�հW���(�k�k3��aι�qU�B�&�&Eܵ�l<{{F^2[Tx�<�q�Q���ޙ������xtf��{�ͪ&u�=�>��8�;f��$�>fN��;��"~����g^����eO~N�l�dKYiv�I��>T�ᾈ��;�'�Xoe�~�j[cW����c�����*m�ꅎF?��=�/�d�#[ܕ�j�#��.ߚ����ڙ��疟R�[��w���hz����^xǠeň����y�PM��,0�7��2�'�EoPy�⊗u����4�uJ8�'�`�~O/}��od��;D�[}r�p��qʃNV;7�����|�WC�7V4go>ˈ 2�����7(}��A>�߃=��=�4��E�.�[���4[��\��(��ô/m*�qfej&#oj���wS��*�0D���E��ڭ��.�8�nY��G�k��Tl��I�(���W]X��0�?�H��]���'�F�}8=��䮐f
a���(���S62��"�A����
�Ae5v輌/�;�<Sw?g^�T6�jG��:�+yOɺ0��"����Q��f\?Dc��������; �vK��>}�cOmc�7����/��IG��j~aQ�!q��	�F�@Zjzj�>��>�)/=��Uz�ч�6��YFK#�'�O���Vdj�SHQ=�7��n9���]�
�s-[J�0�ᬚ!�9��w���-b��P��u9z���_�L�q^���8n�Ѝ��i���7����Z|(�D����5z�D�<��O՛�~�I������c<��W�3����Q��]�6 LG5� ��#��g�;b3���c�?�]А��37�Y�{�'|uvŕj ��ӊg(kިh�c� l E�j�D�8�����@^x��!v�|�=��pM��`+5m��)+���Ru�@���H�$��}"R��:��=9&�ʹ����vp�ۓT?!��~�dA\9:j��(�����4ef�32�4)J�r�sՓ7+\� l�@��H��A'V��B%]z��i�<�7���otVv�J�������4����
½�I,oL��Z�L�[`7��FDO�N�K]���h�˵��w�
�7�z^�\$���na�E�X����+��2��3k*�e�C�6}�{.��H)?�W�G�����en�{�ر8�ֳ��79�z{&����f��ܜ6��ޣ���z�y�<%�2�`��-�5u��r�UM�����*�s�+(V;T�W��Nbϻ�
kɳ�{r���8�4��[Hr�ڄ8�g��P
�ٯ��UcYJY9��!�N<D�v������Ү����{��&G���ʒ�R�R&�c��vo��CG��5@f���ʸ��'��ef��.�r<���c�M��U2.qt�mye�0�@�ɘ�ꡚ�|4ܻd8L����)���#uU�9��Ҩ���%9ox��ۼ
�m�߸S����i������Z�I�*�a9��.��\.�q���6z�皸nua��xn{��a�K��Q3�f!���vroE�ǖ�[���$�Y��f�O�&���U��^t4�*�=��]��P�Y���WOӅ��
o)$��yg�����s��B9��-0gK݃w�\���uM���-s\�VM�刞eDd�P�ʲ�x���Ӆ6s3*��y���'c��k\��N�,�P�Ǩg(��ml����(�,��dW����7��ϟ��������Ѱ�Z5<Xx;	���P�+�R։�t���`X���� 6��zb�_N��:Բ�X����h�Y�Y���8�����Ѝ��?@�̀���S
1q�!A��>)梫rF�q��ѐh��坫#�W�G���4gr����A���'5� ��R!U���ּ�\M+]s��W��eh7����P|�[j�_�%N��F����KL��Z�;L����c��Î��;G�5�[ˬ����М����TI���˽�}�F���&}����!��Е������,,��di�B�\�&�g*�'�(��$��ۆ�wG�/�uG�J�ͥY9w��(]��/��+ؙ��ܪj1�XݯsH�ݻ��wv�JPm�����RM$�{_S��q"\�}{�x��DW�_m�%}��T���Y���r�
�K�ש��䲆W4�n�I�QY���+�mH���tE�?6��^ԏ��-�^��L��AO՚�^;<�h��쎙���@���Â�A��dK� ��m��Q���i��7'�F�<@���u�`v5Y��hn,��n�A��h�uq��y�v�5�3�wd��բsWc;xҩֹ�m��j��5ctb�خT�e�/a��9g�:=��r�r�AaVܨ"]Q����/3L��[���`��b�� ���D�|2-k����b�97;%ڋ�����ƵV5����1� ���m�۷v���G�����:��+�E�tR~[Z���{��e�6�c����6�w$ߏH}�];K��l�h���;�

Qp��~E�'P���l5�T�HO9���j���������H(:"/�=G���|2�YF/;�N�;y������S��JNv�����*06�D����F��=�t���:�g��F��t�}c�A�5:��R�l�&gdW�����+,Aē����e�~둾�� �f�����W��Ћ�4�����2=��/���ƞ������I#iX2���j�#}�XɆ`��~}�;�OB8���"��AR*�T�m�S���lz+k�o�����=��'���6�.{:�T���+��*�����9�:�f���-8�zE�!�������Q������(��{H諾�}g�0x$N�t�7���u-�V�fu�A�@��S�JG,7dc��
��[s�����ZT���)�	^HLMk���b� .;�PM����^lZX@vgG=ׂ�4h)��e^��c���Е�n��+��X$�W�"�A|�uٯfGO�a�_g5�\3�D`�\�����-Q��i����;��(/n5�O���O���Fʮ����MA{�\�ݴv�ܙ��^�S��1�ks�}���n�ѢuuW����%���cQ�4�QE�k!�����V���}���R��a�l���.����ų��vN�Ze��碝&���d��荙}w(��y�k1E�wGCe>��츙)�xb�mFpxL}��EGݱ�F?���kϞ̋�����p`�vc3o
��������S2�㐃z	B���k���"y2P�W4p����sP޶��n�#��{=�Ԅ�����6�.b�H��K_9�e*�ͥ�+o�ְ�����p��QٙTji�T�>�{q&�P^8�����Q��r�u��bSkY0��-�O׋h^���>�5�V�6�q2��Ρ��dU�{B��|/<b�;�	:MO�;#��f0�6{c���`>c��W�:�4:�ݡ�����(m��ke��Xb��z)���S{X%�C��Jq�#�����e�h$�~�E��Ly�� \�̋��M�,5�!7F�ئ��{��6^� ښ[9MFh��\7	k���Iiy��a1OaEOX<a��ԇ4qA[�Rtp-�u�3�&��s�Q���-k�[��<��+8�h@��M��{gOm��?s2U����!��>����e��=��V�������t�z~c��g�y��Ps&��zt�k��o0�l�f��y3�����J'Rg��;�+|�<\�+ ���0>{�0Ŏv�x��S\�ᛥ��ʹ�5����>=hT��3f%��h�u�/�-�>��>`��y�ދ�QU}*+5��Q���b��n[^���g���׿��r��o��Ʀ"�5	�ÍQ�W�peoG4*G��b�Y�{�^�t�{�*�+����㘽�B�v�$� �cy�f59�TS)��޲mP�Jz2(n1��3��]['su�S9��ke�-���@���	1����+>��'��g/���~�6���~N���L�/�P���H��Z�#f4�����ީc�q0��8qZ�<��^�ޘ�N��&5SW���*�78��1�|�\`[4�zg��~��e�-��!�������o�?G�Җ'�zi^���#Mfb�s��%�˟}��;���+����t�ԱJy��Ɖ\W��P΀n��aU�"_���nϲ�f��N�?w=�BD�Ր��q��6��v��nwDw9�Gt4o�S�.-�^0)o�#)�O�R*����P�Ҳl
�h/Y_�F��&�?��#��?��幀���ﯯ��v,�@*@���j�ޕX�<h��,(E�6�f��[Ý�Ss��4ݷ����]К�-��ʒ�SM�P�z���U@��׺zs�৽Ưɧ�J�څءn���'&�|��e�:����#�>	�*��Ҍ�V��z���N���2��w�+<&��T�ˆȩWޥw`�x�I �]}�I�,���{��&:ӳz���I�sdk�#����D��u5�����v����<<=� �< f� `�v�����=�P�R�7hT˴lx!�Q)�S)����N��	�ҫ-���)�U�1��o�#=����D��5��j/z�2��GI��~~�N�^%tX�
i�iOc���q���^��аZ;�������u�x9�G�����X��@���C��yt�:��冠wGR�v���s�gj�k�;�<1�kRS����Ƴk&���W-��r�Q*�=��_�^>�!Őp��Y����|�|��J�c��a8��(X+��	���y�7uѦM��H��y�̘�8�-Q�{m��u䊃ˡ1[!A0+�����VGɋ�0��y��J�Ѷ��o��ƻo��7�P)����h�<�ͪ�5H�U�H�v:0nb�5���q��ف��u`��s���Mot�k�i����E�x���9��!\�؟��ق����mjD�q��en��0��2�7-��^��`P����v��ī�P4y�����{�)L�)_�Dz|&�tf_��bUB������rd�6� FTq��
��9������wa�n�l�ZE� ܽJY&�GF�]��Z��%�W7d�������UԜD���Y��ë�9Y���ĿY��I;�̞��|Uxy/e�疂�_�����K'��=��VokJ�#fJ;�Ϊ�Z���a!�Y��Ќ�5��IR+�#���������W9���Z�ڊ���F�j�h�u��Q��~'� �OĐH����v߳�o����H/����Ņ�f�L�|W�35�)�u~\���d���#W�>ǿ�l�rc�R��}�1}�@���S�R���Z�1&�j��ɛ��#tP\z=fD]�ihs0�"��������K��<��w�Wݕ,��-�R��KUH�1>u���WV!����gGW�_%wo�* ɚ8�bʞ[�[T�a,�k�	�@�8K��,�Cȍ�w��]�vde6rz�P�".���t�w�Ap�u���)�#6�����*l��2�i��;�j�7�m�u[��7�s���_�-�^.��߃p��\��B.)̪)��E�'�����a�m�v��B,ۼ�*�S.�x����]�S�߃����� ��gIgj�o%E�p����p��Q�Z���wiQ���Gk�im�����頎+Č���g�_�?>��:��~�����*��ۅ7��΃�%�-��}�܏d;7#{k�|I0U�f\_��ц ��̳�����Uɩ]����0%�z��ߍBhO@���8^= {���FT��D���@`P X �.��Kg'"쩅�5u�4�)�2��ַq�7�^���7�bX��7{MZr��0$�.]�:J)^kEdw�D��+.��]�z��*ki�m�a��R̽$9���ʘĚǲJ4�[�����u�E�sD�؝�i8�i�
j�d�	lu�.5���5�Pkb&�:��:�3\��\�?���U7)��V>��`�a8&�X6��q��JJ���u0��6������K>]P�\��@D{�_f�Q�(fL.^�D�Q��0�C��P8.���ڣ��&�֬���a+�1��S�!�;���	q���ȼ4���ᧆ�����r��S���jv-���C]"7��N����R���%�wh��g�̐�Z�5g)�Z�E��{C�XN�Y��������.I�r'9�S1]%O��ub�v(ehW�䋵��QHeE�=q�"xK��E�0�s�[hi�T�R�1ӥ�h�z���;*ZX�)�[%|/�{���r�Cd=��%Ͱ�O���b��-SǗQǍ���R_�i:$�)|��Y�R�!;D�wB����]�(�ty�+n5L"Jʏ�T�V�W�:.��e���0���t�w�7�&��vH���5uu������um�3jJ�� J�HK$�38��2�>u�W��#Ė���yN�d�����nt:¬�Rf�ZSx3 Jn
� �-@оyQjng䘲��YW��}*4���@m;Ia�u�!����:�����Ν:�ڣS*�t������ݏq[�����s(8�O�u+�w�5���3���Zq-��9����NL��Ʀ�u} ��FՅ3+0�4��e;�!�6�*�V^�{ZiXYJ�k�]�SMJ8�i����"��՘����dR��<3�\�"�A������i�Rk�F��®I�F�f�d�g(AJ��t���Q����dC�x�|T�Yx�x���H]����f�$��5�Ok�[��;�3b��<��K)U�|ɓ3oOs޺%�1���=��*7�}�JML����2�90��Ε�u���yn;�`Ԩ�Ьݴ����b�z.n�]b ���M�ߤ�xԩ�\�è�R��v	�����ࡍ�[ϑxN�8i�����|��k1˥R�u�&��)�S���&��KՒ�ju���kr��'J�*>�p����-�M�ei%!v�+���w颧$lV2v�mid�0�5�c�*<�Q�=فV-	j[��$� �wV�9%J���/XB�;Ɂ�n��6�˅��Kz����O��=juǛH"f2#ṡ���Ս����#@�s*6@��I��`���\�ُnS�u�+:2<��Q��Z�sFnJ� �t:�-'N{8��G���yO�y�Ɲ����S8[���EnF��[����|1\ε�鼘S3��3���n�f
tҲ��0F�櫓�յ��p�T���[ap�A��ڡO�M���A`�t����]q��f�^:���@bdp��?A��(���w\�����lR}uW-�r�IN�͈��MO:�^4`�QFEOi�&�[t�<��E��2�lh�Vy.�o�h�r4���Q�Gwl�L��C˵�myݴD�"�RZ,m$�6�X�[�sX�<W6��#���}[nZ�w^�[|."���(Ѵ&ŋ�k�j6��뫅��j���#E�朻lQ�-_�c@V*��$6C��cTmFъ�"*5E��+�sd�+��-�|����|�
�Q���)b���R�k��TV�+�� �V�q *:7��w?�'+���>�=��M�#yZ˙#6�_�:�*sr�Ç?{�&����h6]�J臆�t����w�*�{�x�������zr�~�-Al=��|C��R��a�����7T�w���+�a408cF='��4:�.g�����o��BUW<u���ق�K����mO�4bᨃƒ%@�y"�k���ȧ�n_H��'6�{�}So9S��Su��8�/�Ew�<����aig,\�*ױ{�N��G`e����&Y�n1�.�1c�&1z�^J]�4��SPsW)�+�1�a�����s�����5��-�qy9��.�����r&Yxg=Їr�i^p~&7�(���q�o�.ԅ��Yڶ�9�A;�"��9�>K���X�v/�cXŲ:�i����2������a��r���$���-�ʔ�4���d$"(ͯb���EP���/���WSc�(ꕯgaR�(���|�c
3���ϵ�\��Qɫ���^>�~���缕z���O��|w�[�\Ck3d��%Q~������#-��q7�Э���_�A���g����ף�s~������_�G%1��1�) :��U�]^�妧V��LԐ�����%1��9��K��=s	��>�JZI�R������Y��D(�Nx�擓�H�m)���q.� 0��IvJ���`l�t�ܖkX�w]}O�p[��Ĳ��9:�|X��Ȇ�����=��xxf�ieƔ6����J|I��/^�^P��-���}w����T�B��.��uR�MdNC���赸Ѳ�3=&[�ׁ�I�g�<��*}��d]��M���E/q�X0�+�a�mo*�v�~�A����|�C�L4R������9�E��'�c���Ȯx�,!uk\�A>)UZ;K���	x�509�|h���QB���f�s(�dp�a8���Y`��Ҡ���:۱�����!�F,9�o����ۗ�?�����R���ːGs�`��Z����B�n�2*.J{C�p�.ZH9�
���F���jsb�m�?�s��i�V4]j�0�4�v�T]��{�^��o��v,��~/V�m��6�6���">-k�d�Y��$�@R����8�%���'��Te^��V���_k���ޤM�]��[/�*��7��7N���i�8hXr>���	#��ì^9�x�ޙ�:���1�V�C_��u/�������x�C訽B~5��\�h@�}JGt�^���`������:��qS��������I����
{�S�,]dՓ.���ok�Ѕ"�_i�Be��=���
�����e��Z�+֦'��}^���W���j�M3yY�mW
��5u$���9H� foW1�<��9�6;����3���V����Q�Q��]��Q����.0�-NKV�ﾯ�����&NV�o�>�5���%��	ݝn��2��y�[|�dx$��8䗻�֋�Li&C%��8t�굢3l�1��0],^�ٮ�vI�םh�����M�j3-f�<�z.'Z��}�[Z�:�R� Vl]7�w�F�Q���y8��tg� ��x���i�ڷ[);E]�dP�����쾔���^�m@����%'�3���O}MX!u�~f�=B[�0.k j��¼b��Sw9���V��ʟ:cʝt9�e��$o@<�*ǔ�R�cױ�kG�>t�Eؼ',�������=��ُh�
���2�����R�����p��-<�!3�c�ax~Ƒqf)QN��7�ͳݙ�F��y�zUUb�`k��\����E��gk}i��q,gñT7��IzJ�O��r�N�4gN���醃x�S��=���#V$��,@+�k�7�z�e�qIjn�z��;,�[�H��Dj��CU��xs���+���	����_�@Q����\~�]|I�Z�QR��W�k����&N���D�^�K��М�'�zNN�3^��1HS�I�_>W�,���-�NQ��XVFөB�/��N�4���*�ƍ-�l�F� �`.��s��4�n*�㷬IM|�m����,��|�  ���=��`<=cz��"˩�r<���d�[^���o=*g��K�b,���#����a�e��c�8��j#4����jS��]�#k1H����)���x�Վ����o}�4��΄>6�Ŗ:skӆ��*u�ȱ��x�㮈��sz�W���߷$dj�Qr�5;���
"S�WlphL��u'i���w�Dp�=�&�������0�o9��{?]�E�mJ7�i�ΫeDw�*���h����G��hv�W�K�*Y:(cqA����n�dͿ�=ݻD�v�z�f�5�����K�:�p���z	=��^���R1JW�k�Sa�'�q�#���e㮗���h����:���F���O
�f.Uĵ��a\����V�P�\����^�m�n���U!�VU�67�ֵ�� ɨ,�b�d��n�s�Kb���7(CP�y�{��]eu�O��l
��>�cK��&�ls����k�yO�l�l�T�=�}�j[�Z��Ggn݆ݚR)Kd�õ�������1�܁O�ی">�8���U|	E�%��)�uvl�\m���zp��w}E��w#\�ٖC��Z���Я^��A�����hw��j�士��bN�fiڙOQ�67{i��;}2ݍ�}]�uN��$��{Q���̥�.��+���]�W:��1wo�\�� ���n�s_]W�}�W���{����! ��$�*i��0�B3��ʶ{��*�T�)�x���6�ETa5�Y��{�]7V�0�PM��F�X3�M��v�Ek��4>�Khed���n���b�ZG����S��șˎH^���j��]�\�Z�7(�L��wo�n|��I�dY���l�y��:ɵnf�`5�)�w3��n����H�y��B��8�jBr�9�sǕ���:I�݃	ؼ}��O�=�x���K^5�yi��t�vI��[<О�l�.�MsQ�{g�k����[��n���b�>㛂Y�eG��3fƔ�#�����8�`Ki�������!Y��޽�9~��U�].�8_�Lx��]d@]Ki}[{/�A��C��M[:`Ѣ���̸Ro&�Пݱd\�ٟB�j�X�'�+^��0��)���H�&�u��gK��w�	��J��s,���S�~:�IH���ޗƖ���y�����Eő�T;��.>�j�w\3�sˆ��j�d��(os�iM�~&w��亱�W;�ԥ�]�f^�˦{�m��'B�^���t�O<\}I�2ĸ+GM���,tї1Cۖ	��*���֨�W�+HS��H�DVRv:��0�}6��F�5[��5��C�_m��<�NDY#��$�8,�pn3��˵��=���� ����}�Ή���q�i�׸v��7�T� rk	�QeB˘fk���J;c�3#�O7H�:��+�v�u�8s�_r���RRY�*��[��0:�c��A��,�/��Э�Y�5'6X���5��؋�=�`Y7/�Q�.p�/���P�����z���q����+F��ȕ�(���t�kYOh�B�ҫ�=��DSF�S����ѯ�w#�Ib��gL���!t˾=*}�9�U��Ps2���ȕ�+�\��r��z��qF3P#��J��7��K���7>6��p��z�1l�\rC4�ڤ��3):�'�c��G��Hݍ3��͔���يj������$��5c�}u�>_��|i0�jS��%�Ή���R����%���u�}���D*�NG��ݿJX�� ��r ��4���1FW(GqVmW0(�e��11cwH<�y�>��6W�\�a!D���L7k��`�3���g^�C��]N�/k�d3�T�U�ܦ���u� T�8�9?�)j�A���c+H%����1�o���:~��lum�FWL/?A|��m2Bª�{�����8��U���4�z�F��[l�{!Ė�5}�Ze�m�8�S�/�����u�i�������\)k��w�V�U]��G�C������Vhsv�K���Xoh�n
���'ݟǓ(��*�0%���/�&���3���6t׿x{����� xh�\�JW�QH�1qE���J�mjb�׋�9��6�k
M�!gٸ����Y�ʳ�,�h���::���,ljB����[7�7V�Y�8m���r!��	�V6�Hȍ�+yKE+��w�W��I���EЗnXD}�z�f��6��:ǰ��$��z�5x��C�Ϯn��RxFp姥�{PbdD��5��ح�׶������%;��tQh�`�I#�V��;."ȟ��B�ۛ�l}��]��,��إ�#]�g�/�O�n�H�2`ϱ�֧��;Z����X�w9�k7����Cz�P7}(�i�	��o/���)L`�Q�:����݆�=��DU/G0K�N��AsB*F6�K+ެu��'qeD<┨��x��Ώ���W��cz�!�t�˓U�v��nDL�J���*Mc_�	d���i��*���Y�.�-���-��s�w�yޙc���0�ٷ!fT�ݮV�ev�+dph���:�ఐ	�L�
�d\�]6�K.�����E'��2	��M�����h�Õmpŝ�?R��/�Pz�T��xNXpJ��v U[uRq���qL���F���|=�YZ�7���y����9�5� �Q���*�w���pN@8u�3ØW�ӗ��*�j�����J)�1КX�{��S}u��늲C�ѹ�����J�bĺ���#��k����K�r�!�w���{6�n��x��{����vx�m~���#�<juA(-~�#C���W�ևV�(Y��C�=��ss�	f`�J��e����12�c�b�i�KB���� ���;V^#k/�pwt������1]��,�$v�:�������tZ��7Wu��R���]�����a�Wc�R��'�&e4�����CU�MટrQ�x���Ѯ�t3�Rך��Sߟ=1�}܍`��LX-f@C�j��"���$���6=�^(+�D�e��F��g+�xW�OO���E�G4z��(�}l�}�����יUN���ŨW\|a�)�\�R�Pd2d{�a3��z����'��jYܶ��mGEvc˝��6G,���ռ"��&��4�dv�^.gX"��5;�(�Э�
j�������v��_F�Z�
"=������������=���D���w��͹G��)��Xy�苽~��1p΁kK�E���AH{2�aiY��5{1�Ő�ڑ�����˥�?9u�����չ�(�s�j���!l5ʀ�'��t����X��_F�6�|Wڽ����5:�,�Ӊ�h�O/�2�ip��{����6�&JYDW�����n��]����$�[����v�~u����3&����k%t5wZ�R[f�D\�[e�d�Lv8�[b
؍.F`M��5����k�Ŭmy����������h����%����wM�Ϗ)�P����%$y�^�ɦ�����\DH�{/^��v���uKS0������2d�f>!+�:E6e����Օt�蕯gaMK"X�Y[T�~	ek]��w���r��[��v�(���.�=�w���Ri~��ם ���hu����|\��U��Vt	5ɳ�qF*�S$ëVr����i�2��>0�/�~ȧ{j��.�^͞8��H�R��ҩs��<%K;j�0ײ��;d)��@Ȭ�+�aF�_��_G�$�{�>���xKY,���z����&�9֧h�v��cL'����y�6�]d9�5�y�)��>�"��3�X�nX9����lȍe�l����}h�6�A.�O�Qc��)�R7�	�YVE�����M�lCz�n���Jmץ矕ԉO#�Ȧ�0a��nSB{�FK-���K�W�1��=Jɗ�D����r�{"��0��j�S�f�+7��e[Ü��������V���L��]���u���>N�Q_w�ő�tKr�_BZ�Y�O%�0/F���.���t�ٵ�~=X������%h����u�7���$ӖGZR�����=��̼#�F'�kg65Vo��)$1`;T��,H`^�n�%z{�Ԟ8�2�9��4^��n��b�/6V�d�.�oB;���$m���T��jCE:.��Ó���� �v��˂r����&�y�4�A��H�e^$c�]d@]Kg�V��y�]�5:"xv�^6��g���N��z���q0m5�"÷�T$:b����s�wF����a3cZ����i���b�޸˵���SS��t�b��e��Q :�����[�u]��>��	�3k��	�]�S�n��8�4�!� ��g�f��xty�Ge(*���y{IQ�����Ⱥ���4�k�;A,�S>92�����FD�֩�w�J���J�pH�w��Fb�I�Dt�K��v�ETE���*:��m��F�X�]�G��8�=�|�b�z]8�Aލf.�"E=�o���z妲=x]��[���҉��Uzl��/n��V7�J��怒h��Kv�<�˜ݑY^*���em�je��oF�iƯK��-�6]w?6�;Y�ߺ'~Q���b����y��J.�)�&�ؽ{Ur7�NK�����H��~!/߶:l�r+u_�m7��[>�[�C5q��C�"��x��s�O�E#v6�]n�\?3����,�VUuW�r�\:@Π@_�ؕ�1m� <�:��0#�!j��M>�H6�=ooS�jӴ4��t=��
��+\3�ĖXIw�+_upCP��e�R�Ut�^�����)�M�������D��Ta�97wQOɒfZZ����av�J8!Ab�����Pʾ,����Z���L�J�ȱ�tl��{Y�xT�sӎ�u6er��Oj]խK��<m:�;6�s>�lrA�#�ϴ�J�o�1\� jLT-��9�?�a��Nd)Z���f:ҵ�r�EA��d����W�0f:n"(��s�����:(!���|���"ON	5o��ԅv<��xD��Ֆ�w�:�T�ua�UEP�5�=��㪁}�ɢ�[;�}[���x���ց��E������̙�Y̴�7[vs5�K�W���	�� �}��6\�h�C���an��[�FU��m���Ͳt�O������po)V9���)-Ef�����Z���V��.�n�}&0���+t {�hU��_L�mL�����sN2�,570ZR�ٜ͗*p�ۏ�ya�X{XE1����͘�3q�҃�O_m��B��ѭ�#S�Z�r�KE�!��L�������;��J�Q���*���ˑ[2����������SB�cn�e�v�!�O�i���w95xXɷh]�t��F���%�t�X���H�э�Fցˉp=N[���ύA�Yǳ�w�J�l"+�O�geq�&^I��8v��Qy,^�ͫ�Y��:��.Z�l �k)5
����r\v�܇�x�#�w�$q��x`N��ڕ�+iV����mo�_<��:Zv-v7�_jǭ8�wM|�n��L�'";g:�˚䝊�V��<���>�%MG\��7�`o�}��44-�dtg4,Ђ����F���g�&`�o�o���j��'���n�e�th�yDQ�N���pWN�.�m�i�;��n����Z�\o����a9<�R�]����D=�
����\�ܷ-��[S$�tJG-b���/G^T���+Iَ�R,jGu	V��XsL2���{��
��+����U�I�l��i��=�zԵm���]8�����o�uf;i�*��2KGxl���ڣ�3�*iC^Ф�5�j��l�z�U���A��KS~��z�h!Z���8_/��^�s�R�s`�L�3sW��f;YSw��N����Xl�����W���ξab��Ś\d���]0�T��g9F��E��|ph����Hr�����O&t�I.n��n����e0������wg�I+k]M7����X(R԰����*�t�Y�Sq�e���;X�A�\6ȍc�w��	�r��2̎'�b�r���Js�]c�|�H �A ��%�X�PQ��c]z]��,�	i(�9�Ƃ�XѶ+&���y-��XƮ�\�Z�]ģkӒj�dѵ�&���:�;��Ѭm�鮖H�t�s]9�/;V:r�Us�w�s�W6�u�-��-���5O��6���Hր�J��t�h��L��W(�F�\�W/)nn��Z�דnm�u6�rѢ�]%����SYw^Θ�V��(�.V�%\ӥ��Q�^M&�j�mr-���n��'�I��J��F6�F�m�����&����N���+u���R��w���|���������G|�*�Wtp�{����vY�����i��Ja�����:1٪������^s���X�{���o~����  ����^�뵿{k����<��|ZC��L,�&)��s-��<�A)X�#1C��Ӯ,峬�;��)��aIw�{������	��CNj�y�؞ESv2����Jy�]�I�"nq�;�����o��`�7I(�ԁ%}���	b���[B_��͑5����gq�"9]F��%Xzr��-]|�P��B@�1�I6�b�8A1��x�D;尠�ϲ�Ŷ��$*��j�(�~ݪ�ûeҟs½1�&̌���N�lpL`���G����]E�^���óo-�6R3M��<k����Lk[�­Li�Li�!��1�oT���>����*��&+yBjIxf���lg޽�21�VBp��$��<dk��j�Ɖ��z��ʟ�$�X�?}��?���r"�7���h:��jsr%�P�my�co���1��ob�Y��K���J�?\5k$7�.#�5[�:����wf�bé�����aw4�:��\����-!���D�j��>&2*���Fx2��K�!\��������R�_�w���ݬ�#w��������Vbjf�P��ܐw5}��4>G�׺�7���=fv&�}�B�)�Nc�ܭ��*xr�SZ��3v*]�6������x#Xg-��{x����f:D��OZ�æ������*7ӽ��"cC�O��<?0 ��ى)W.������-�[�+�6��N{Kj5JTa-�R�!oE��4q��˦�/�k`5�JL�m�53m^⥋���e��U���b��C;;�z��#���Z��^Wp�ޠ	k�B^˾P�4	��
�LIa^&e2�Uս�MgW�����3�v�Ao˅�^Uo���j�|��7=�G�x�+�d6��0X�ɟ0��ڝ��S�
J��v�۪5���ME�g1��+q�f)�b3��ѳB0>94����͔\_�R��ST�D��EBw��w��gN�����7��rXg�1+c})?�;VdF3k$
pv2���L���t^;�����p}�!�\^%��?@�S��S�L+b�؆�'�Gʹ�٭���X-�li��DֲƮޜ2xVwK3�b�1�����s��鎳0�ΰM� ��_�2��(y.9ꍫ�YQ��(��b��2�bL����[c��eU�j�3�H�v$��*���^�������~ᇂ�@Pm�&O*��N�=#Y��S�gی�z�ɚ����ٍ��8�ߛt���uCn�I�������!J��5�8ɍ��U�;x Ժ�
�#���t���KVR��"�.�U�o;��Ŏ�h@��}��N� ��m�Q� �jff�/'u�h��*Y��C��O���h-�t9ņ����x�l�۰zN>�����K������z������?{�~�y�g-혟�O�╟�pGU�͓c!����^����wyX6��.��w*r銄��z�P��;x���v�,!�U�V���m�[?&M0u�f ���"��5-ܸ)gƽ��-_:�K���Ӷ ����Y"��)���S��Vi&j
�&`缤D�;^�t�����ҵ�MH��mQ�p�3R
m�����;��H�)_OɈ�
��{�ު�[$ة�܋�]���SQ�h��0��3^�P�����n{�k��a���# ��x/�b��`�T�n�c�\��0Ǡs�KhT�O"����ޚ\��2bķ6_�m*��Ou1ym�![Ҹێ�,�k��<4k��Tj�Hoe#�
e����:����y/�Y��ݘ��=��$�]�!����;�m�r'~V��H��R���hߖc+��ϵy����WB
�%εNuz"�u�,�86���,5�q��z;����4��WC�	���O=[<���%�(�q�d�EE��/��*��Ŵ:�]m�y����]���xLWj�~\}l��h��gBU/d"-�س�"�+��,e�mz�&p�w�� 6�uk��;]�q�Tf�rM�*p��j`�+�v�70֎�a �����*gv���^�ӻPٻYW��TFD�
|�bqX�����_L�b�EY2�ɣZ���U}�|:.�W��m[��/�i��~j{KP�r��O��]7����]���;�y�XkAT�SRᛦ�#v�Kg�Fb�μ%眛�Nxtv���d�٨M	���8�b}�K�e���:tP��#g��$c�t��j��v���z���4.��Ra��y�:͏EN.�c�`ۗ��fL5�tn5��M�%뼫X��^�]���ϛ���
�����+"߆�^��]�Ctk�5�®�6�g?���q��p�MH^$b����Rۧ�w>}��FWVEٺ�4�����.�Մz���1ȇ�F�J�B`�<�1��G�3��B>S�v��5Y.6��L�Ɔ��yF;��Yw���z_O�S�Er�P�l��Z1>���1�U�ګ�fx>QdC��z�(/���3t�J;^�js��;���������j�X�Ig�W������]NIOS�z��l������P�2���k�s�=CzZ�Ƴ���7
I3�%��í/��޺d�5R�3�;�:�:���z�\JUd/y�K�(2$�_�8�'����.IuG ��.�ν�'n�؃�*X�!�&�-IR�i"��#(讫+Z�z/!}�vM����]=
�½�ή'\���θ+�	��t���֯.miV�
{ұ�;)ö�:��ձ�2�62����������E�ڽ|��OX���S�BL�T&���rTj��/��LO�
y{t�ٽ�8SQ��ZGn�zV�ȘL���I�H��Un�������v]A����6ӍR�3���:�%��o��7GS�f�V2cd���E�
�"l-��_1߻�7S��cj�`Q�5�n���	�ɬ���g��������@��6�R���Iէ�cC��>�F�n�STߓ�����!>�����E����]�oJ<{UB�s�J9G��0}���$R��O0Yq�mJ�^�A�P|���7����MYIQ��7G�Bzra�<^�<����.���f�s�J8E����= .�������9��8��jJ�:��B�`���1yo������`�9�8b�ŗm�O4�t�b�����J�Գ��Bo��b�5�c�ņVI�x���*/F��J�n
��z��E�^����A��z��3f�k�z�Q6`��B6��}��餙��_��q�G�8<z���r�	��Lc[�g��5%��	�5����\�}X/�Q?u��\�>/_*J
!m�ͮ����ԷsYE���o�G=��s�Qv�j�j��������nv 0Q�W�Z�Ti-w���K�{%���3j<i겣����yQ���Űt`[��Gw��[wͫ��>ݣ�{�����,�iu��~�"5�����dP�^?����8F�YgX�;�x~��3�w�e޷=8{�M��(,U����k 86+P��j7��B��
�o%�B��ֳ]r��!�)8��9 ��w ��IX�VL&�~�)��o11/�N�Q��2`�i�	8E��}�%Ӻ��}/�� P�6�n=�J"CF�S�P4&�x�Ξ�OІ�4�:(d�s��fum�r5M�`-Bx��@�s�R&���dWT��)��c�^(���{C��T[s��&Wl��Tψ��dO�oA�b8�d���'��[�@���&!�|w���b��V�l��ޭh�j&ݛ[mЗ�� �ɵ��Ė�&[�T
t\��Օ6�:m�K���eyF������!FLL>�W�t�U�C�O��˞E��4��G�1`9�NX_�����Y��(�����݂ZW��̌��1���<`%�/z�"04ݎgay;Ƒqcu�m��T��ʝǺ�׉Vڞ�\9��gñ���,j*�''�S�c��fqYy����\��֒�S���pT�3yt�]�.p����Nm���N`���m���F��_��,4x<�c��YY��lsPjX:w�v����򦷫)�@P|�]ܔ�v��ՠS��#M�+.c?�a���5�l��bV��y�%�V^h�Mz�.�q�ʘ�Z�U�< aǻ��rI�3?�o~rzC��O~��Wm=#-q�X�j��4�+��O��e��M&��KQ��;4�Φ�[uM��2�����CU��
~nY
3����>�r�&�@���W�|z�:1��f���?�Y�2�����w~�O�5Ig��y��q�֠H�v5��fx�D��g9�V��e�lx���W!D��]��zO��#���=L��==#a��v�8Үv��m5I���MK;�V�mtɶu�����r�WH���#'�[�jN�͐�������$��K�mȱ;:����#�m�	��y�f#�4Ȅ+yդnv�Y��(w�۫�A���2��m�p3�m��8	Dy���K}����&j�{0#^�Q�&��UJ�csyR����feT5{5*v�	J�)fک�=���'�9�;��W�v�p��=�(b������R�z�>�a����5��<�_|Vg�[=�vT0��."7h-��&��n�[�]��z9�(q�)�X�<�ʺ��J׳��&��,[,�M��z@s����W�E-��`L��q�1d�OP5m������of�4���a��Ďp}	�;Y��n��:gi���	2�x�7Kz�!�<�&�1��6�d+��e2��FF9YL��eL��/A{�� |�U��w�A�������7�3���Q=��(1Cڀa���b���R>�c���\do�'��f��؜CP��蛊1��i���P������E6�Cz��U����BRpGtr)�/1O0�l�t�fʣOt2�����vK�E.��R���ZrWH�W4��79@���
�=B��~���Yf�m�~ʤ��g7wu��P���:��Yp��Q_w�y�,�ܪ���t��1�����&��,Y�U;�89�t+�y3��1N��!����&�=�`��ZF�v�4�I�{�x�{I}����Yy{ eK��K�~7R'�zqP��0a�Q�M	�q2Yn�m_h�;�kY25F;�qy�֔wß$��`�ǄC皤B�]��篫���*S��^�n��&���)��d�׎�����例���� v�3�N2J�[]�L�]l�4����3�+�/��#C�ۜ�,�C��T1����k�V;�|�Q	$�x��]jC�sF�{��7y[eƅ�{���;�:��ӽq��hA�.(�	���	=�W�k�B�q��l��[C1#$��rm�`�we��cy�h���P%E1�o��w+�sP� �\���0L!��ihN�\|V�U��N��3S��k�w��$R�kN�֏�c8�y�N3�)Wgnс�f�܆�{����6�:s���*����k�;B���H}l��f�Xv}��3��lb�އv��T&�1l��]Ǵ�����xVX�Qۨ������;�ǵz��2��0��(H�zLk8?ߗ�Jת/�S���W�T��y|r�nR���z�r�
��]���U/G!2�� �lՋ3��6�����Df>3�.<��r�>�%�]-���Ho��+���}H�_GZ�%�t��k��g�F<�Xn�@��}�v�j3l%�KmfKG�~.�@2�/�%<��c�y7ʡ�=z1Z����)m0�͌�Bd^��)?X�X��;�*�eC	��y���7�<pʼ�.��s��w��$U��!nG3M����%��U&��y%�m
ǥ]#w����k��D��Ľ��qfB��AA�|z���=C$�/��i�R���E���b\�dJ7c+71_v4`Y57��=�7�j�^S�M�Gb�Zb�c�y�^���A5)�>x�J�VV��s�5�c*��
�c�"�h�&���!7GZr��>�f�}j1@�P&Gg���ː�[?Idⵓ����W�ԣ��������t֭���4'�蠻6Vo^S�
�k�n����wQ���f�W��0,�M�iLq<��Sd�Q+W�I��e�;�Ω,)�5���Dy�=uj�֩�z@Q���r��x+Q�Olf��N�|�e�����fm��q��؇���2Y��;�a�L���L$(�;9?Cv��C�[��'t"�n;�hZy���G��;=�:����q��.+چK�׋�n,�E �XA/���=ѕ�������e����u�
�m�2���걩A���Q��^�M��~/T� ��	�j#ry����f=�iLtVr�T�W�i���VZ��6��ק�60�V#f4ιν��D�T@�u��W�h�&qsGSW��\�:��� 	]�21Zx�ҧ��<N����ӣ1��w�ϫ40}���W��k�7����Ej"j7���fЪ\�e=�?U]�vW]��-ʡ��{A�v#����I\���rLߍ="��$h�EG�ڣ8c®��:���e_��ds��Q�Y��|#�j~�z�!"n�VC��(�;	0��n&�$3�����"�%<�o+��@�:[V�Jxݶ6��W#��r&�cȪ��NLyvҾ����_���9��e�C�b8T�u�8Ϯ�ɯ�M�*X��#�l�6u��
�b�ثne���}�|���@}-�]:��36�/��ٲѕ QL��tl��0�ԙ��_hkk��f�]4�GӧH���i�8�Y�fdjxR�$H��o�;��\j���?�Y��P�}+�}����[qq攮���7ZEhT<��w�<�����d�5���4;���QNg�r�nx�8(�7�S0V��}z����:����sv|a����j�s�c5��(�Жs�\��;��q������7��nb��ޡR7�#�6\�p���5,P4@Žs�o
,�4�6)%k͵{��6��2[��`���o�/;Bܬ��]��N�����	,��u�VU'*wuԁW+xY��J�5�44ݲ`Y5`x0��F�y&G%�;6����C�*�av�{��N�Lƈ�H����7s$���s�rf����uu���rp��s&\��Z���V?��0qm���6ٙkrڒ�V���ֹNG�<2��<��[���_S�j���q��W�N��ꘞ!-���Z��ǁ���NPD�\h+2rX�=XƬGN�w@a������B7�-a��ڲ�2�ڤR��{F\���
�g[':.���f���@��3sE��Aҭ�1�/L��69Y]��6���㪠� �+s:"�w��jj�
;�'cK�\o3���N��Z\Zr�T����)p�%t�}�^e�v�SRd�f�-����������
��@Mik7���i����i��6��֪�R��
�ԩW\:�(J�	Zjf���f�����{�a*LQ�����P^�q՜B�]���w+[y7f���o�ȧjrX]]�,gbۮ�@��7�DDw�� �ϲ���SbK��+ws�U�J������"4A������T�M��}��{�h졍mMT����k�O�n�[\�b�Yo(o)R�X�H'����?�ܣI]�ֲ��5��a3W|��S=���\n=+N�toAeA��@�׉3@9�f�p�W*��X��{��uo�Z�3��z���/Xk:p��ɞ�{����#B����p�T�Ƒ�U����%;��)MMه5�p��[W|��Z�+�8���Zc��P�E�u���=�J��ܺiu�|��P1J��Pݴ�[4�#C�pp��9n}�ff�w��wqg������XX�WN��i��[1���N�k��ٰ֌B�˹�n�o]�t^�P�ub��N�j̻�&�Ky5��u��;Mu�sf냮�Ҭ8�yt�8�NL���s�Ӵ8G���1p5�؋B�Ղ���Z�s��d�����Tb�iq�#̒�'���.��5�dWVi��5�g�>�N���xiC���]�5�"��N�	ϱ�,|���h�]�S%*�����{N�^'G��m�vE#�od;0�=[չ��h����a���(�E��^�Wt36�Ōe�K�kqո�8��������&k��U����1 �RbC0bH�|�}�t��Hlo�}yvŒ5N�{O<�Tb"ɪ�� .��F�o��)^y��V-�\�yy׋N���nj9�1���U�񍱍�����m�׈�6�.ѹ��nk���mp�+��׏���Ӻ�65Th�r�n�W9cTX4F6�ܱO�k��j�mʽ��uӕ�b����t�U܋nj)�X��X�.S�W5���c���u��6����9v��{_=^�w�wuF�V���j���ۗ65M�����B1G"�W
6�U�͹\�[�.mͮr��P[��F9��n�ە�u�y]{�Iuӟ?O��yMV�ۭ���KM��xIN�I���sxwd�޷��볎Λ	�K](��L�o8ٝ��:��z(�0�?�A��}����̦��Bx�/��P���"iU4ƃ�����4��R�US"�tSc�MҪt�I��ш��y������+4�j��_������ �硎C@�����������v3�A���S�]C;���\jۨ���7}i�h&R[ބh�`|rE@M�^��G�K��h���O�	�Oj��xn~ގ��å�EG��}�%��_!�����եP��?�o�#YsRơ�"�Q{~*y=(��Ռdu����;�$]\9Cf�Hc��K55�ϒ�犢y���y�LA2lV�K>�-s����[�����hޠMgk����ȣ�wo��ސ�'�/)�T�����U�r�O�j�ϕj��SƫX�m�Q���y�kpF6bɾ�u��d;��s	��A�U�~�<��H֠��i��[>�,է�b����Kl�:'�ݘ)q��\�7?zD}�����;c��#�C�If[fr�s��*�	���t�*��rn5pZ�
"��d�M3��f>�zY�_Tw���X�o*�~	u�nPi}yO��ӿ(.��kѮu�7�@��PI�3��Y��í�g?G�����<S� �wAwytN��n9���d}u�n�o�	Ծu}|�V�\]��ׅ4�yB_V-[X��)�����ܽլ�������W�ߚ�z�?����#�f�`�%�X��Ӈ�������d� �|��ւ:���B���K�q�u��̼�kG�2��x�1}���tG��:a�R��=�=g|�T��������*b�b�.��V�M�G�1^�)d�^%Qf絑-k��N*�uB9C�9�vR:4�Ko�JU�CUJ�@>tĝ��`o5~����=���,�dن𭤮v�z�f�oo��1�}Y�>��)&c��o��)Q��BF}�q~���k�<zd�nC[R�ݝ�M�Ψ��@���c�l��7j�u�kԑ�_٪R�{����c��m'��3sY;�+���B��T�������������79^;d��X)������R�����r~�R�{L��|K��e�ޝ'P���F*������P)�`ל�<:f�d5�����ꕥ�)x���~�m�N�tS�{9N�7(��'�r��^�;`�k��_G%�gy���V��ṅ�hg�2Х�^K�ϝ�E5|d�#����{�퍥���-���G[G�P;ˑ�sS�X-�n\�튍mC3�,�2gL�K��s�{�-aa�>�,4!�1�>��Y�:
��Q�h=��f`�5G�{l���L�Ď���I�]��Ѽ�2�Z�.��o$v9�ۨ��Wmަ�^1c�-vn�ҝN��:�*�h�������K�~����x�R'��d/��!��L�]�)N,���©0�a�e�-��.9:9��ܕME��G��3�p��mx��6�tH��IZ��K��=�I꘭]'�5�����ތvg�)�8�n�c��}�U\�S�/��������o&�齱w��'����X-��G�O�x�-nshqg�w���.C؝BF��ai^�`�����	j�x̳����Ԅ2&;��!�j�[v���)�@:������״���N����}9����א�YQ�1K�WpGF8~7��A��I��{$�	�6>�B9�	���_S�*����R��W[K'�Ƌ�+�Ξ��[V�-�po)�k�A�9�v����Z坻��膴L�k���n� ��xk�>�?J��Q�Q�VF����V[��F�]D��wKs=�������p=��F���7�f��]-�_d�{$��;���҈m�-V���6�����ÓY�Sn�r�e^�i6�d�\��(����Nc�#�+nXV�c)�������x����9��l�~�s�7+f̌kʶwA�V��!��6Q�{�Y8[���̻��/�D����6�v�1���Bқ@�{١\��̘p�-��v)h��y��	Sa{Y���^@,��9iq��RI���0�����ԷC_�W�U����%����U���6�6�k&��4Z�̤��J|�K�^�{+$mr�2짣�UP3eTf;J���{��p�yg@�y
������Ƃ댆i�R��s2���,u���sKnZ�\fc�7�����T���\!���ǧ!H*/�=��s��ۦ��q���;S"�О{��m�5{�!�6��8�r�u!�aIP
�y$��O�,>.qzǞy�byy�Ҥ���ZP����+���őûcOn��u%Q�V�i
%��IF�_���5ƕ�&V]am��^�������K����վ�����P��P�o�4�bAXA3T�(MIDKݒ9�2^���>k⨦R4m7���n2RhNL��S���k_�Ŵ#6����St�F��;���ѹa�Dkb���b�X�<��qg���*��zw؂7P0k��t��5����o��v����΀�.+T�G��UG&�,�Ch��q�iP��F��d��c��K�$�Di�,�}�8*����b��1�Z��{�ţh?��9�> V^�gZ�ӠM���Ho�{�X�Fu�%z�r�.���{޽N�!f�oZ���>0ݔ� |�Dc����Y�پ�ԣ@P��Y`7 �wǀ挡36��{&��6�Ғ��`��P`[����݀�ɕt��M���pRއ)�a�ћ� A���#rO�M��-E0a!���c���:��4

�`�Ĳ�C!�\�7�i���*}��I4���Z[�D5�bF�A���{�m�SZt�|�W!"mt�8|F��OL;�Č�}���P��%�A�����׎�g鎥�j��Um���cp:��������o��V�1]RڌR����ἓ���h9�9薶�ze%�P�ͫ�k�S�@qR���K,ኵ���,Y�<�n��҃������ͭ�,0�����&���^��k?0��=2[����дNz�*x�Plyv՜:�Q�.n%a��M9�Θ��ke�T]��q�z�CH��|.yZ�����S�e����?3����H��m�m���������<f>-��ބl�`|ri�.���0Z9�uk��à�R�ON򯹹�gݏ�>��}���EB�')�<f"�l(6����8��V\�f����14>.�������{	�D��^����2��:/�IP6Ŋ�7����#g�i�������� �n*-mxR�jN5�IQ��c�-+Z��n��?_꼔M�/N��d���m5!�Z�=;\�'�Z�!�շb �b;��u�V�mc��A��k����Eb��dW����P��Q��!��W{��fRi�pح�:�ӝ�ۓ���d ������E���E���\�]��i|�{�x���?�_:�w���w�,UkP��z%�Κ�嵧�;�m�9�+Lw��]j�N�Z`�;crQygDl�od�h�#s�2HY9�*6�T��V�M�{��߂k��z�\3�P���<Α���3^�R��gd�6��CWZ��U�4���v�:�2f����c�K�����Û�J{�E����4������XL���1��s���eMh�
�N�i�ل3nvn2:�p;P��ԃ���`���|1M�
^̮YjgŔ�y+|V�358�T���{�b]�
���US,ȫ͔b{����:	07:����$�ޤ�ڜz/�;쪬����/���Y|�@|�M".z��{�r&�r��qK'���J��$���Fɢ{��{�E՞Y��қ�EҖ�J��.�ʒ{���bOT1��sR�wL*ֳ��&�����y��jWz��]�s&�f��I����j������u�4]-�{������[aC̸Ѯ�Ql�{��F�Ŷ�U���$���K�ދ7
�#�E�q�%㼑����9ؿV?b��srF�(��c�2�p��"�7�ӑ^A��WKD7D���m�f�\�-uʗq�k�U��iDt�J��|��e�//��
B�9y�^�i_��@�ۘ(�mr(�����:7۸�h���"恝��ӻ(<ŉgAfn��k����s\����W��0��$���U|�Qi��.�z�i��������{(3��˸��=�s���^�a��:�ˉ���Q��U�0P��f�*��Ŵ:��E���P��W��1Z�6Os�C�;�.⟎���L�~���ٝ,�o��u��]�O6��wM�\;9�\�����3�q$��1��'���Q�7�MȜS�s`	͍j@��8�G�)4��ht;x�l��eK0��sx�Bt8Kر$m!�k^�f�^.�-h�=��T��`�5.*�n�E6����r8�]V�s`gD��JJ��mbTH��W�_,�����#HC)�iv|���H�Ъ�����P��Z]B���htT��z ����@�A��D�*�#^�4��������ǘ�E�6s���)�j��@99�8���c60���'T�@�"��	^������5�l9���;� ��[����Ot�W(ߖ�[�^^�%�W�(��*�5��͢�Tsبj/�Օ�LU+*V>K+�j>
�z��?��A}��UD���f�=���_
��9�:�50�naun̿A��z�=�~;�ly-�+�:w�������~͖t��wY^4�v5E��\�/�ĝ���42aI�r䫫�~�t��)T���!�U�ÑXFkI��U��[A^0 IV:E�.����q��g$��X�p�p q}5�rNV
�~۱T�h�}�	����ȅ�����Kx����4�	Y�d:���7N�0I�i��CMc��TA��w�΁����),���J��o�0w�J^�c�%�u�A�agJ8��T1wέ���u�l �^�E�+h=�~��Lg�9�4G�a`���g�NU
f���͋:�`��e�ӷX�[X�L��lR~�[B���q[�jI��ݶ�`�g؋�Y?z�eضk��?pVc��&ܳ@�U�Z�d�ks2��y)�&�ؽz�(n�Kt��b)���ת�=
�-HI5Lx=�T��Zd�����79R��f�u`'�c��ns}�d)��a���iy�w�ݛ�C��.�,9*Sta�=��1X��?f�5�.�q��H��̕;�W��su̎������	ޘE%�Ҁ���	��L�^�1���J�6���ͮ� �;#v�X_#%�/Ö��>��H�`�7kf��E,�}�y�G��Q�
�+c*e����whW�b�	��7m�A��
�е8���˩nl��a��+�p�q��u�	�s �m�ɥf�OU'&���Q��v{�t�)ʂ�h�V��.�c�c-��6���P��@P�f䕻@�<�N��j$��#H���b�ecP���3�w�Rk��ʇ����Ζ�&b��Uv��y��n��0f��7��3�]E1�:z�z�����t�{���&�j��*q���䫞˫�kH4�0|�ʟ��Q�Ǥ m��\�&8'�Kh0v����֧�5Ͱ��[7F�|�3�r�;��n9�pL�"�Ef�.+P��AȷZ�B<��㕕�fV1�VC^��l���v��yp�+�X�;�k徂�beZ������tV�15�֍�;z�u������o���`�Y���9�%�˞�r;L�� ��;��Q�CT�CȒ�����2w�gdM�=6b��K8��,7%�[�T`�.;s�n~�#ݑ悯�}(�i�	���*�f$�U{gյ֯�JO=�oM���e�s�U6��BSM�m{���;�@����0%:�[>�p{���;+�헝�H��ژ*g�0
�ɯ�i�X�T2~ -�e���$��"Y{�}S�ը�d���x����|w\��b���)���OƠh1�#!Ƒ23&y�& �$r��f���NE�io+Z��'&�w�:D���=EG+�,X�}ԉ��s�9��; P�����y�|e��A�ʮ������7��͏�S�¹< SYሙp�[�GV.�[W|s��f��mCw>ܬp�ʊ�-]m`O�\��w����j;�4����e�ɉ�D�V��*-+�p4��r�b�s�:N`�)0�7DAn�����苌w�K�1)�*�7q�m�s���|�j2�ِ#�f��!Y6FwvƱ�q��TおU�����ǆ�:�}��Р,br@)���9Q[�	"8��y߻c�_T��g��.�0ޭ$�2	U��K���u����E�Ӊ)۵�X�7�wA�Lq�8&}���X;�m�u~�r��5�J���qEܶ0

���G#����N�9ɾ���#�0O\&,�u� ���n�.o_I���?���S�_*R�S�;��wYי�j�ƠH�vE�;m�-f�P����Z����t8��3�R�F\7YZ$�e����z�[�xn���ml6m5�H��ְ�*��͇���{<�L9w�Y�psc�z��Q�r�4�׊44R��������k%2G��<��[��_]j᱘���������O��l;o����;�o��(i��00@�t{�Kb*�	YwC4xOlT@�d;��Ӱ_���х¢����w���N�A)!��K0����C���0���U*�]���!��W�9����l�O�Y�4D�r�Y}�`	)��ҋ`i�L�o)�����7Zx��`�)ʗY�x,�Jd�S�3)d2�ז��mmπ<�M:�[�+n��η9��B+yڗ���e�&2�ՙ����i���,�I�h\�,i4����&ffncv_L4*�؋vs��!�Y�,�YwI=�N]2���T�;�U�ʷ�h�,A�ݱ�����Տ
�z33);U�䘂W�in���������1����TCU4=v{z�)\�d�ɍ`��u�e1b�]����6oB� /z�mCz���Z᳠�I,��'Sc�s����޸.tá����#;�J����z�V�Zllk�U3WS�|��nJ����vS�����*X�li���V�\2 ���[u�2���K¹��t&-��ZL���[+���m0h��V��t,Gbk�����ĳn��Ռ���6����7I�F�f�OKY���:'t'eV�R�	׀�\�@�5J<����{r�Xb}/�;_;���Υ.'��N�S��������Wm�+�mЩ�=a��gp>"��̃%�)V>��I�<)��櫋Y�Vqjnskx�$�|��z��R��,��*M{Y��Z5�����H:�zt��|�m�8���3�k�(Yr�9��&�����(��Ae:E�i��N�6�{6_It~N
jn��a�+*9GQ�X>7ȉ��[l���mX��H�E/�6#���˾�rU���J�q:݊�Qy �:V�\U�w)��wN�QM��ǆU�oJ�O�n��hg9�_I���ƗSL��]=��u��>�y����E� u���j�l��V�{�R�� ̨h@w1�@+t�A�m�q�ׄj'����u���F�D��������Y�"7�,'����U6d�q<�6�콦3[j�:�t�'��@	��g{X�7wڄv�骲՚\��f�9e�[X��溺�W��ޒ�0���g�c����S�R�ZJiGC�k�����=2�,���k�S��^��v��:G5:VqU�{�������C�EWkU��^�������ۜ�j��N�t�ob�����Y��;��u"��-;��캍�8{k���C��1�*�3�j,����&S:��z&P���&ݴM*���/�!Aٓ���V��T��Q\iC.&���8��ca���j��?
��=�-�����\�t**`�5�MR�9[\PoZ�&��-T����hTv�vvKF��A�/��yo����g7��.��;,��w._D(��PcRYW�GNGc>���#Eav�u�*
ڹ(]A��GQؚ���8+f�1�'�� �muoH�5˫,]���q�t�oP�K~�:��gF<��{mɂ�l�'zQ�Vε�>9;*_^K��d�sy�3�D���p��̓�_��|}�z�v�k���ns�-��nj.t�"��5r�U�ܸT�ѹ���͹cb�m�栯��ywX����cnh����M�����j�o��r�Ӯ�c\�ۻ�6ƫ�ƫ�r(ەsU�KF�][���.r�����s�1�]�m��94o�vƱh�v����sW1nj���b+����������-��b�\����F�Ź�ni5��fguF�"�����
�k��6�r-RElcF�w���Є@@��A <E�y9��w�����i�A��op+��u=&3��N��6���r����nȘ�b�P==Iǻ�_��k4w����hm������E���j=��7+ux)�W�C����w�v	/a��t/~V�����_~�� V�6��#_��H|n��bp:�'�� �����sÞ<^>4oW<�[�������Ù����k�Ѧl>ɤ��'���x�o��o%#�C�-6��7T.�4���d>� T<zF):O�tR~�R)�{�n�W;6�z�=����/��S���"�7��s�6]�1��Wb�a~Qqo
J{ ����u��ʶ�q5넭|��pl���˓�����x�f>�L��-&��YF&��H���|b׷vbﺺ�e�nov�9-�C�N;�o���G8c�%�C]��h8`[�&�m�˴��+��P����S�T.��������?�.f:���<�QHҲ����+1GУ�o�Z�� װɇ�G�&-P_Ev�vmC�h.�q���?��%X�$n�v��j�Q��z�6���B�I�j3��n<��g�- WRa��y�:͏Eo�MsQ�{g�mY_:�K��5�Z~߆�rc��O�\��;l�o�T\zhF�j;����^��)i�|����^k���^e�G_���#��e%u=�����h�����2�S��d�d|v_Tc6f�|��P׬�&�a�L^���-��iL��Gm�ޟ��5�\|n>s'�y��C���N741���#�p��~򑨃��M{޷�'�b\����W��}���Ud@YK����;U�jrslv��z�<�k�f���"5o~�����4/{׹h#�6��`�a�@v-i�Ht�VK61ç½�v�����$>�����[3�:��m`��`��yk�V�%}!1�W@p#�ȇ�rt��}v�J�u����L�y{�FG���M.�~&7=(���q�o�.���/Ϲ`�4����r;���y��w^��foq�:rq��:a2��J�f>��$��<�;	R����ށ){e����$A�-���M�O.����{�z91���)>��'�a,}��!�{��Ph��U}�I1���S�A>��yp��ǜ������l���ǵ{�<��H� �oR�2z���Br��]�U�yWK��j�g��F�,�S�֣X��U��t�R����^��B�<_㽻]���	��rh�?|���(��|%�e�2A|`3X�Q{f{W4'�P�u��"&5�M I��>�-�loM�|���N<v��;5���[Yl��T���|ō��M�GzD��f�pJ���g	�L���=��63�u�d<
M����G�����;.�"���[�\��ZJm�f�R��ͨ�Xc�n����Ϯ�g�D�*+�7y�Kn�}�W����b�"G?5sІ���!��^��"�r��R�wD�#J'%�t�D�%�jSq|QR��7;�Ԅ���x3�ǚ��tq��*㚩M�k��<L�8s�c��a��������ˊ-W0(�nH��	a�C��mM`~Z8���Kc�c�4d��Tf^X�Ƨ6+g�s�
�ҭC���;�z�b��P��F0΢h����9�lϣ�i�Ϟ�h+%������[r�=E�C��cR3�޵�u�UM�$�Ƹ�Z^�k�{���t��n�0m��|D�d���f�;�N��7VU��T؎&{e���r�u�u4g�R�KS��N0M򆍧���踭S�!�?����v��6��K���h���tUp�p+
��<K�<d���H�[QцP�8\P��)��;�Kj��i�i*�2��I���=j�I�> |!��;���r��ծ���OH���|:z׊H���_����w#Y�8���2p���������h.لG�T�/P�>�*���{5�|-G�b�������	���B.���I�\�S�;^��C[t�N̮�7 �v�\'}jN�	�>[}�v��r�v��n�C���M�8ܦk�]\�R��,����A�;�H��ni(�r������g��������eT;,�.��>=�;7�p�ưu@���K(V=�v<�ɵ�eé�En�|~ry�ڥ*0����Z%z~��VO�e�R�b����ɦ:.KowL�{O�YA$�osF��|�}ۙ*O��x��4!������-F�W��=�X�,+B���D�'��<��0�(��3-���5����T_L
��:��|h���l�	�>�r���L�Y��ˉ��qE��Ϻ{��q�1�2�����썵{O����.~#��Z6}�m}�$��;������O!�Q�\j������ǆ��RÃ��EG��`��1���G(�ߧ�m��1l��xc����|Kȍ���A.�:�������H������Y痝x-���c��C'��\o'�5uѦM��K2��(݊&)�\�k�)n�㯕�S��a�	���Y�y�D<󦆆ֽ�궱ܧ�����4�
�U��᛫����%𾙣�%��5�p�Ŗl �I�U�~�<��j��ǹ�싫�+�;m�J�]�'Ӓ;�x���6��(<�pޓ�˾l2Mz�Vf\5�ny/u�x߄4�ʄ��Xh�P����w�a��x�&��@1��w�cX�#n_Kôsev�b��V�E�1�b�#'�� X��'v[n��f&l]�{�GU��%�پ��'U�=���[�/X�����K�F��͓lzD����E�-y_z��J��IG(;9����v�����7��޹.�{dX��&x�R
#�[h�Jdӈ=��SwR���^�f��Pk�Y�q�D!YΉ5�U!�۔pjj�L�)����O�T�2�y����Æ��p�Rx$ρ�L�-�).�׸\���2f[y)f�	J�C0��<�6���t'S����ژ$[<|6�/T��R����y��
iq��_�W�5�:�\��G�P��d�Y�X�Q�'䤴s3����a�Z�a��>3@�|Ǡ!�C�"�FM0Yu ��Y��v8K{�i�$^-���瘿E��F2Pd�^5�s-�\�Q��	A�ܟ���u�T�Y"^t���c��Vl��9[J�-��f$�߸�'%�.�OؠK^��1�ʝ�֬�vU@���HJ�|k�}Y���Ф��u˶�l��_�g��R�:T�{E�'P���l5��\>��5�^�����co}~�S�#��c�����]�K(���Z��EE��_u)��+�u�s\������.�-�����W��8h(���'r+��De��rkG��G?C�2]=Ƕk�	��Dw�*<|q� ^o2`?_#����1,ՙpZ�֛�(��%�j�άU;�d�r,���Q���mG�*�+h+���o8Mm����3�Z%�Z`��������#���!h!��a�U�Q�΋3����.�����!�slUevp�h>�0����{k��w�N$�*���f�S)�ߪD��(�4�2񝪨��dS�J�k�g�����=z��=��U8�$n�Z�@|�٩���_L����sm�T��I�v0�ðlsru���99ö�������%�o
��
�$��s���¿h�t�
B���}���&q8�	�x��S<�TX�FF�@�>G�x�����W/�/�+<�V�C����_g���)�Z늌��dR�>��ȍ��]�g'29��2}���<i�q����_�����^vϬf�K$~�����}]eǺ��]��P��|�Gߋ�9nZ{"�JN��|��9{��~����GT�K���A6�%�[8��͎�l�Uӳ�3n�G�TH��yfE����z���Y��M�N$H��,�(j��^�Y�;ρ��ƟH��IGݱ��KMmq�t�E��:�+D=Y��glئh�m���N��N��)o��5Q���1�7\)�N��]�؏'(yq�gJl
<�
�;�uոz_¯TK��qR�K�{]R��M|��';
3;U+�s'*�����hǵ�J��w�nγMG8�F�}u�B�Uɾ���U�S��+ d�S�*�m�{���`� �^�E��[B�ѬaMC�C���J����hLb^��p���}���|W�}	�2$�S����8�d^�ؤ��$VoER����>M�QB��ooDG2;u�Y&���.��Pr����ær#h��3(�`J|�lӓJi&�|��\�GyuϠgo\�R)ZBUo5J����P ��07��#�����W��uVq�[�+��g��}^*}�)���Ss�,5�!7Er'�Q�syG$Bp�'vi��y���A��s�%��Jm�_s��ۜ�M��C��xRP��)	�=B^t�3,.�S[�[��g,�v)��a��0䊮�F\P-W0�#E��xC�jJ��S�QL$(�ڲ�Cw��)�ګ���1���b���T=�l]�T�������ydw8�	N�5��z��g6c"�7��PI�$p*�%�oq6�V����\d�����^ю���TU����M)J��:n��KS.1l��b ��`�k6�m�³���]��¾~^������ǆ@GO���k��s�=y�?g����+հRFe�[�����Өէ\8���ӿ ��W,  ����ѹ|��Z
�aۣ�|�a3gÔ�͋<H�F���]f�ݕ���q�
cr��Q����=�H�����������0�U�s;�1l♲�Ӵw�o�_u�U�&e�.'��?�#Zϯ`�9�.Ɔ0M�Dڐ�`7n�P�yY*��ۺ(q�8v��y������4��
 n�����<g徂�H�Z��l2"D����2#VKE�;�0-a|u���Y��.� �1��}�j�\���`xw9 ��$�Xҵ�3B�d�>٭�"�r��2�+��k6؟�}���j��ͭ�jmb��P�*�$M���p�Ӱ"��?>�U�����0�YA�[��轵�V���uV�gܪ�X��HY ��+(V<�=�3᳚�R����Rڏ�JTc�|N��*y�W>�k�S�C��O�m�p蹒f��qv�u����|=���s,]��Cȷ�}OP��.��'k̐C@�[@�[��X��)�fp8����2�p�T˜��l��DO���z���y�Vr�Ѫ��{�BmM��v��wb�U2�Ҁ�*�yY�-	��8���7qSM��N?Y��|o
a@�v?�����+�;���ٽ\e��4z,=7"���z��S��N���T\�}l�~m���}b��?��O�]	4���af�@/=:~PoG6t���~{�(L㏶�ͤ@V�i�A��k��0��kU(�Q��\��/s���4I~�\��Z�VΒ-u3��3'���s3dJs��u��ۊ�^��ܬ�a7�:�o�x�|c?!�����}j����Ȗ3��W���"IU�����u#��a���T�;�]����x]˒Lb�;�uBxD6��Cf�\Wx�6y�UI�:�5}��â�'�'4�Q�����xz�4n�`�.����S
-q�
����5�[a#��7��U�쪷�a3�ү3T��U�@q�vF��ز�̀��o�H�qV�k���Qu3;�ٞ�O0۪h�W�=���Oc�g�l�g�lP��&���g)mۂ��f��2ޯS�u{)�X�
8�q��R1*@�������^(ȱ#�'�����"�F����Z^��������\��zY��� B��Q�_�/3jQ�c�$gtzP�Z�)���~3N-]ue�Mv�K.pT3j]� �tv����U3�6�����3^SM���>=��3�H�L�Y}y�Fo�⟆!��}?&"�*bL?<�Bj=׹l;B�5�\�Q�D�-2�n:�u���;:,�S�Q&��RȀ+��q�R��j�G˸��!�B`o/�dp�y�D(��A���L��\A�<���������IL V�ͮˌ���HQVu:n�h��0Wq��mѱY�峴�a;�>ܥ��A�rty��^�2v2�G���NeZ������й!D(B�y6@�έ��3)Dtu�P����=�F�n��W7����oowuQ�/���A�,xb���7ê(����> ��d��
�s��.����s��`Wn�hk��Z���m���\�"fӜZ�%X_1F�}�ǩ�]�5kQ����/)�G��=�~���۔�dEdr<�la>��<�U.s�-9+�V+�a��
Lc��(3R�&��oT�yiY�L{.�g�a"4����y�.���Q���;5��S��0̣ͷ����_j��(��C9HE:۴�WN��t��K����� �I�9�M��g�v�w�#��e����%�ba}I�܌_�c[(��CbH#��끲!<�?B�Y���8�199Ŀչ�O�^��/oxB��{{'��\k��=t5��{���q�H�|݂��@|�Vd^�̕��_	�
q�]S�<���]�*�[М�\|������M�K��h�ل:ǵ�7$Ϧ��}�W8��ЇW9�T]����-8�	ucx��U�S�hO��ѳ0�o/s�7�Y�x*��p�H�5ݫΌ��q�d{j��� ���/INli`�`�p�Pj���Am��=�����q�iZ.�+F1�gVc�d��;\Tū��o/��dhUx�6V"z�zV���$���l��+���P�5Lt��U��Wӛ��!�
�ʬ��S���]������qK��S	|NL��lᘳ-�-
�넮�Gጹ(��b<�&�9�Z�=A�"�_3��A����Iv��BV*�g8�U�ڙو �d��fZ��`���V�l;�Q���l'��*T��ѱ+��D��)��0/굼�㷏:�l�ǎSK��P�'L�uj�|���m@��x&�𕒨������8�F�@F��d�n�@e��H�j�S�O��ۇc�3�Y$`���)/�����XK�3�������5�9C�!��;E*j`'�.���r�oȱiv�PF���5�:�n��&������;��v�fm�K��4�SQo'��|��z��lO�2�{w����e�Gs0�õ;T�89�v���%��=��;�)mJW��D
�`h���̹��oubm.�� iU�KD���A�Û�w�kð��s�0��R$[��v��[N松��5D�yu�r2�]n��x+vv<�f:�\�xt*�j���ǈk�Ε\dEx��;�!����sDkHE3��љ�-�֟Y��Wr!��훊-�o4�3:W]b������$�ܥ�+�_+)N�2�.��$�({�f9�Te�m���e�&�Ei�����x�;p�$ξ�:j��,=,a�����WPe�&�V�k�Aۊ+X��F�K�C�n���:�\�Y��m:T��7�J�U��u��i�
(<�ugz�u�y]6mp���8Cf�w</�o��;�}��78Ŭb`]�Σ׻c��zR�Pm���=����ʣ��e�+/p�
�և�S�SX�+W�����!�6�(�}��݇����E�n̡��L��|�)�������D��&6� ��/�w�xS 5��5̪�g׏w�r_��*�XN�r�^�F�X�or������Z�!�v��뤎�D�9��v�A�B�C�hr�L\�Ei�Z�Y���L�6�N�s膦�cƃ��I�k��x<W��63������������-�N��omtUp��,�7����@ӭ�GEE
f�l冑X*9Vh��{nԀ���X�e�3/
אE���]�)J���]�u��t,�'��e,��9�u)�5�,��P�x�2n��-
&3[9U� �Ǧ�-� �����!6��M�e�l�Vud�^�(��ݛ�b)����V˚�Q�a���ê�N�k�UFV�Y��i���E��rCH�+ܨ���&�>��M՘���kH�S����g���Z��﫞�q��[t�N���C#��%���廛űr�̠�c��rݚVl$e���ThP��X�WJ ú���64�4�q���rhi�80�2��'�:Fل�ŰY��Z��M�nܗ��.rX3BL�nM�Y��ue=��K�;y{���׺�O���k�Z5�ۚ.[�m��s�E�n\�9���3.h�jRTQF�U�滺����j*)ݺ��.k�Eܮl��EHZ��F�\�mt�jB�iw%F�\�ss�h���E�6̂�w\�����77+0Dm�bmχ�"��j�gv�aM��j�뻆�6J�N���[�ڊ��.Tp�r����4�"4h�Qi�D3TFlE��p�^5�(�1�r�r��mW7"�FƠ1.nN��(�؍�p��e&9���&�%!2����Hwn�\���,�+���׫�����SG9����`_�N>v��7Xp��B55�0�+��)�z����S( �=�0>��*�+�T��ѣF��@#�#.���]}���+-*���_�CL�g<����v�[����Z�ľ�G\�/ڶ�e�t�v��\��a��R1BW�j�����!���^����k���C�ө��GH|Pˌrg���S��ޘE{���]?c��8����Ⱥ�Sı�ٍE0w;S�k�fJ|qmh��ճ���tä�2�r�-u��RJly&c%�[-�=�(�\�ؾ��M�k�"�o��̞��[��g.�u~��Be�lQ}Y,�kSW���iP姗H�ЎV窬�S�k>���{�� ��S:��Uzl�4�ё���.�)�-�{�}�MU}캸'^u��t��T2;�SG�/x/��1Fao yi,	�W�[6d�k��:�z�5���c�Iއν(^8�b�����v�^���">�a���R��-�E@�_�`ǣ�OK���Z��&��.��"��x��s�oG�=�"���Xk�~Mр��0�7s�4�Y/�4�Wɍc��ZC�ޫL,�&)�(��u��ʹ��qK�Yݚ|=o�@aQ�ev\�l8~�{�N�m��N�V�m���in�%1ߦ�̭���d�#.ڝ�θ�&,A�U�t�Bm:�7��ع-��7¼�
 }�A=�fh�Ȼ�X{\�oZ�]³]l��M(�5���������CG��w�'m%7d�ܕb�&�HԄ��/�\rr���xkݔ��p���n"KW������@X^Ev2�׺p��z{r\YK*�j�Uc�gFf��ʲ$���C��n��S����$����@��b��P�[��dw8ģ���vk�ޜ�a<���|�����bf�}�}Ne���k���I�cR���]?S�͐�Yy�r�yf�:�}BTɣ���W���&��`(���6}�sL�ק�sP6OF3�w�&������g�{g
�?F�i��D#��7��\���Xu�r�=�$Gc�]��m~6ֽ��Z��a�^�z`c4���x��o����8)�z�[ ��q�}ͮj�(Χ�%��3{���ft��k���̓^�S�~u�Pn��,%���bJ�9Z�s�묿;����齕<�p8�U��]]�>�}y0Y����)���sa�4d�Ae+�O�}]�{j�U��z�쀜�Vb�T�U}9��2��R�kj �Zid��B���<��W�����=Oí�q�V}s��N���mm/�m�q��u��VM PޕX�V���o�[����Og,��G�����jsMc�I��T�Z�Lڶ0���vk)�O�B��Ž���t�l=@�ny��}.�1y�ï���#����]�n>ѽo\�z��)�4�s�pͦ�����*uҲ��C&�z#o�̛���<���v��:���}����
�n}K���ߛT�4C���B�o�T!oRi��j�"E��TE5g׳ޱ�k�L��:����-�%T�9��m���G�ή�K��Ts'Ѝx���v+e�����b�ׯ�C!غ��q�^�o��t�Ԧ��U�퓎lLSt<jj�ܵ{M�0�JHߦ��<<�·�t�p|rE1Ō��!O�6;P��zs�����5��:��M����F�����?/p�V�brJt|۵f~�f�VD��S�%�A*y:w�}7�)ӐV��T��IZ,Ί�#�_�ؿ��B�\o+��ɹѦL����2����>�e��u�~���6к0y�����p�F��`��1`���y�~����٫�ʽȉ��L�Ÿe�y�]<��j�ϕj��\fu�.]�`�vZ̀���[W��u&j*p�}^��}�g�/J�mC��r�s�ۯ��W��
�6'��e-40#k`6M��J�7i�n�`vs=�HF3�딈�iv(�.dc.|���.����f��~��>��2�^��v�Krv�������ܫ9�������k*5�n�㆝��7�G5H�<X��-�7��԰1c��=O�|Ga�7l��c4m#�_��{o<��=�c.GY��$V��Pf��k�"ے���+gd������dQ�=b
��Y���.�ZǿP7��xE�;�h��ˑF�^���P�[�����w�L���b�N8u�UO��ta(e�<P��/~*�L���o1�%nl#��OI�}~ܸ�#�=�;���!O���]�G�f�
~م�2��}?1�Tǌ?>��}�먚#t�vFtS���<�+Welj��_(r�fׯ%�M���PDW?6��^�_5T�-��P$�Ч+n�|h�+���ܮ�o&PygH܅XL�����V��מ�[j�l����uc�dZ��W��}�r8�'�'������O2��%������̃�	��I�|tR~�b4-��Q��T[t�W֤t�o�jT��>����s:|��.����r���h���r��1�v���بo1����+Y��g0n�ju�[2ڸ�Lu���SR����D>�_�j<�%�5�s;_�����0Q˲�jv��UVNcNӈ��
1���zX��Z�����ʟ�3�E!���R!h6`y3�6���A�������k<���}P���b����;^5g����$��(�3p7㘨�5���_mH�	�kÕ�xT��(���?}��
B���]����2�]SC�*�ʘ��yI�q�f:?^��$)�����N�OՔ�P��5٫�>Ѽ��}-��;�e�a�@�h-d=ف5aY�Լe
QȞ�]M\Ύ������P]<��ڗ�ڍ���C?m��x�4�~O��Ȧ�z��٨M	�d���A�����M�`��_duPJȌ����{Q�
1��S�y�O*~�0������g���o�X��ēp'�^�{IO\�p�:�6ͮ2Fָ��y@y{#<���BFE����"UV���L�T����'ó��P.�r �a"i����[fC�sCv}��P�bN���t��K�/3�Z��d�hV�סM'�&��}T����0��� .;�PM�+.|t���T�+�����0�&1z�IJ>����o������mJ���<#����c���#0�ݻW����;�m]5�9!��(,���l*���#6ͪ'�u�=�@U�s��y���c2߶&��ʵ��\[Wb�cx�KQ��z���܌�}?_E$��<�1��-ޥ-� �շ��g�=0��K҃*�N�;��.��N������B|�VP���	n��&�Iv�ش?gGKE�}���BG�/qY���҉�����g$����8�b^�ؤ��N�qx�����>?�7�k1 镵�����*4GY�{�wF���>��w*8�U�h��+2@��Fۥk�g���O�Wl�<᾿�������}۲�I���=�4d-l.��kR��K��V^�¯�)g8j�`$�3�m@�#6_k�;
�ۍ=���dӰ�}��
�zܘz�����|�u����)�D{�����|Ͽ�s�s�Fd��
�����!s��w��
�q6ؼz�(m���z�>��hUP!�B�"�Y4Ƃs~�PVw;�ƍ��B�(\�bt��)�?���_��U7?Xk�Bn�5ǱE�'Y���/@*�f�Q���5�\�E����0�a>&�7'�b�29�<�@�X�C�;���Mv_��eG�O�UN�WBˈU�e�GsR�P8m�	�fδ6����=ծ0��jJ�z�lI���z�.�x�:w�9���!9j&S��E�}�Z��ޝ/K#��m���Ns'w���S��;8T.R5s�&,0VKu�S1��x]=2���-�qH����8�i5Y;��ц��z���^��fGk�Z�n4
�;Mf�B���9z$�%)f�]Sj�z�nm�3%��[�e�b����N��V�F�i;���z��i��ۭM��1�1�D���`�$v�g#��o�	�YY jc�T��(��URjsr��:%����`�딠�\]���Be+2����f�@�Z`���a�D�֊���f�n�Xm�
o�A�<�V���Me��_W;�m������i.�n�7O��)n������X�TAR�r�qd���gnP�/%�P"^���˳�r�ٞ˻C�"j3��A�TsS�;��P�mZE�	M�iFi�>�&{�Y+�����L�T���b����o1"%�iݪ9Wq��aH�|���g]/ńf�R�k��I8�b:���)�e���{5�>>'�;
���*��2���%4��tg]pRl��D���N�sRn�s�Տ"���>z���/Y��??��^�9��i�BG�HHK��V=4/ �󉝓�����L��{4��x��E�;�z��c�$�*y*�/U�6HS�3up�8�|$K��d�3)�aUL��yt�uydx+ߋQVLG�@`Uo��['� ^�o���<����(ݪ:}�p"���ğ��w�TΟw��u�5�& ������e�u�+m���qoL|фp׈r�>�	�����&�q`�*)�DUx�\��6MG����D��]���!�{e��%X�}��Vg��md�ĝ�]o_�#��.�O{�Uݑ[��㦱�G��k7�c�W)*֝Ig�رv!�'�G;7�n�L���tj.�j�g��ȄW�&31����� +�Jz��w� �>���=�.��`��l>f���˙��(��`�҂T$�~HL��3���ց\ b�N�̷i�d� [{j[��J9�q��$�D ��>�C�݉�8�ڻԧ>x�Ʌ	��K�2aPP�z5�N�=9ѿC|3�'��K��[�
�j�`���&,� (���S�(�ǠxŘ�ʢ39�qYf�p*jdn��1J9��쩜�%�f�Y���G_�Y�b����T��F�M���0c����G��d�������~j���o\}���mj��؝�j)�����9��)�q+A�D#��*��V��Dt��:hc"��#����i;ccv�$�6���lS��wW��*�;6�ԦM3�1�mF��+y�"kc������>U��^]�>3D��: ol{R�eb�ҳI3P
�&^��ɨ�9c'��y�wLko24[���lZ�y♹�_}}o2D��񀳦,0�qA�ς�$���S��t^�<>4��ڵ�C��d�n;oe;3�a�v'��O(���mN�D��eK">�m�)J�#T�_@��^�&�w��*�;�<��p��^���ͼ�ps�֩*=H2l�jۙn�%��w�ӎ����ESS)�e�'+g<V����l
��>���,z{h1'^����I��H��Jsګ�w�욿#��5�D��8k�h����[��*��l|ۤ�f���م�*�9��r��X!yR��.Xק�1L�x
��H�Jt`U��3v�t�h�>��:���Y�f�u>�`��_ro�]�	J�_�~�[2�v��y�����V�W}�M��&���{ݺC5��}���S���tG�z)�ڤ�v����N�0�3�R��<��Zrzl�fN9�lU�����.�ޫ`Z�J�����>@r���Bپ]�~Ժ`�h���c��Ls��
΢�]ݞ]��F��V�+��a�u�i���dJc-װ����A���/�w��.=�
7�9�l^�ZdC�'Fи��6ق�{z ��n�՗�Q����y2�H庲��Fъ��R�X�׽y2�2�w��wzMs�'�(Db���j��"�1Яu�9掳&�"8U��bؗ��º���2��Ɛ��"a���v���[��__�v`��Rѹw�f�e�a�q� oP|����;N�g��8o��bk7-u��֢F���TՒt��]�ηm�^�FAyg���q��<F�8EX�ru	�v�ڮ裳�Et�d��my�k�/�����H�m26%�X|#�X�CK넷(۵����_�m���B�Ɖc����E�V{���e�]�w��5�i�4�c���m㫾�t�2v����~��|�}��bu��4�;lv�|�ŗ���5o��(L�Y3GU��Z�0�����B�C�.g��A�+����-{G���1>�I���<�*��.��/��'qQ�2�bP�����3;z-E�ūyDo��/<H�Ҧ�[23c��.��wF��G�7�2ا}�����*���z�MMmKhAB���㵯�o2i�C^0ڎӍ�ǅe���N��e��5�2���j�����t��W�R�8y���n�v�hi�XzZr��⎓��m�[b��q��$BC&�}��᚛�-��F��\�������'la)%�[�U�\��QكT��5��L\H��)LoG]���1M ��܉��W�+v��l�7�f���Y�Gv�e�p}��;�vu^��lzTF(�vnqf��H�E�Wk���IO39�h��P�*�f˒���q����s�#Ƴg�Z��wǞ�r�g�O�#�c��(����CM�mf��[Ec7 �2�>�ޟDjOG���qI�f�� H�h����v�&�^X>Qإ�t�}��z�s��!��̱���p9w�`�[�'գ��-�Nm��6u��X��-�fP���{ID��ܭ���3��;/�&���U���]@*��ᇮ�u��_+��fT,�����3L���Vs���L�Rd��E��X��N��zq�=sC��
�IY�fEa⮲�&C�F�R�CK ��(ٿ�̶D�^�`�}L�Vcx�֫�"�:��e�yE�E�|v�G����p���|l^5�w<��� ����2�=X�.E٥�l�7j��ū��� �����G8FԳ�<2Y�]4�GHZn�S��W?�9���^-ɖ�����t<(�t4��j�,4�с��]X�
��75L�5�5(b4���/!68��!�m�!���ň�s���x���1���3wj������־R�ۺv�|̳&�@(�H���g;�.rNX`ԹsW1�:����w_L3���:n��ɐ�	��^531͇qĎ���� �eJٽ�՝]Yu�U��L�],X��v��Qc�Սe%���3	�t)�kg�Ii4^,/.�3\���e�iz�0D%� ��s{��ڀ��M㵷��N��@�B����k"�1��2��&� G�Y	�m���gBwN���6���,ʐ��mf�Y�^k�2)�-�Zy
k�%��l�|(����q�/m0(�_}+��M�A�.�h͚72��H���`67{�e�Mi�i�5�Jw���=�O\$���5�We�E>��;�:Y�t<���1�+62`���β�Yc9����,]5S�������z�%���eL�����|�D��%ʏ�a�t����Sm�AK�9v�{��wn$5S����@�z��W,�	}����k���A �]����,�ᄍ��Qt�ˑ���ې<��!�����Ѡ����ۀ���i=�5`햱��r"�r�y��T�f"cH�o4<�&lY�^�j��������8�Y z)ܨ��ӭ8�&b�/����^�c0zq�cQ]Y�j��iP��h5.���._0���v����-	����:j����!7�w����^B`_*[�nl[X�1����-��G~�ZJФ9�%�&XĻ;m2.k�*]
�sye���3��I�ӌ��(��N�˸�H��w6�t��z�V5Š+�)6�Bʢ����h�a�c��1E������z� ��&������HX�=�p��@?��s�і��O7B�;���;��֎����ܱ1��zqf	g@�vw{�"��̽[K�c��č��3Wek�ì0;��x�����M}7u'�J���*|L�<������ft��ƛ�O����t^��նwc�S�� yX�L�![��edf��k��N��6E>��<�f��9t�$�o^F�e
8��sR�:��u/,`Oiҥ�����gF.'a�ddwܩ�
X�����Å��=Wv��I⺼;���џ_��O���%�{U�{v�*('u��$ܮ�$wZ����;�).k�1o)�ur��-��2��s�#wup��wv��։��$d�*(.n\�-%��wp�ڝ��GÁa�(������.h���`�r�b(Mwq�F��ӝ����I�ɢ�r��u�*e�����b7wT�f\�h�%��c����1Q��!�jMx����˨�D1wXƉ�	���L�e���ݺcE�ݯ:�H��8��"�K����%3D�c1�WBH^7S�:��D��	��r�U�F��F�����bF�u�amˤ@|Ur�e���ڕ�q��W6k1�O0,�<Omp�
!����mY��RJl��I�s�a���n(�;yh�7R�9�ԵV��M;έ+7�cu������^G��l�s�/u��V��Bj�^�����k���;Ӑ�?h�>�Ƹn,1+����٢���j�0��N	�r�)I�-�/o��7��0g�������d\�f���܇�|�>���0b�;�8�v���;�J�!�P3[�c<��ׁ����E�D�&%�t�M�COH����1�ˆJ� �LF&Pq���;�x=��v�L�a�Hk�1�LM��ngO�l�N�1�!���[r���d���gCbcE_���e=-�|��*����M�vV��4J�sq6��Ѝ�5�m�5!�d[љ��k"�S��,w�f^�r�{�k�"���ݩ3]�Qm��yؚX[�$�U�r���fUb�xl�|�pu,X,=R!�֊^]멺���R�ɞ�8���N9Q��Pqp[[>7V��ʼ���@�"������Խ-g�7�o=
�ne�b��O�|	L�#���5�y�M�ӱLĚ��~����?y�n���t،�|�WwI�ؤ�h*��(���`�כ5G�9�b0�L���kQR9˱�z�%]&�i<ܼx�v�+"�L�|JL�L���Y�o$�F�v�T�>�k��u�inR�g%RU���S�ә^ƶZ̻��زJ8O�f��l��Dp;7� �.�'x�q�몷ŲypBA�{��g�mƌ�VHܤ�'ٞ����D���'5���Y�|�3�>��'���؋� �qۘ;���A�g�g�-.�n!oP�۹OP;/D5ȇ�\�ZK[�{�/Eh�w,�(�B�7<鷤�8s:WL�3%�z�v(��h��ى	������:�5IM+��E1�}��T>.�fY����xr�̃Ws������[�n�XOe�z�6ȡ%�[@�VK&��;Գ'8���iƌ���Q̋`_-�QM|���vj�h�J�{��h�<�OCb�C0	�B�>��V1�����Ⱦ�m���Dti��׳��.�zt��= [5Н0�0��{fG�1�=jv���+�~�T��5Eeۡm�s��!Ս��<ޤ�qy�a�R�V�	45WՅ&&�ۭK������|�ܙ�B�����pmY`�G)][ì�H4��E��xˣ�b�v��B��f�Ұ���5�˼2��仡�br�Dks��鵬�=[]aW J��틫�\�n�]��C�?^=���[�h�����3�9�]Й�.��8m�l���5�YM2�mA�$�犹�[n�b�x-f^�T(���R�ܝ���[N��V��nig:��bW�I�K'Y��MyL��n8c��f�=2i��㙍\��jM��3�铚�gx��*�Tg�0�\�n��}�y��\s"��d�i�D�"�m�9Б�0���V3�9sf53������Zx����o�N�e ���B��{��׉�Z�T�Wo?|��[R&��V��>
�m83I͆��g�0�]:�����\1gu�>��n�Xy���x�]��}q���l�Ӳ��h2z��0�]&�{&�-b3MNI�Q�|K�+ZWq��P�m��qw�H��u3�w�i��֟���$��>�ހ��j�rU��׹OX��N���9U����3�8�.�r��ݮ��Ŏ٨屯�!џk`qK��)�N���0"��!ףU�d���
�k}B��N�lC5�޽dS{X�����5E�u��nc���}�O':9Y�\�{��H"�;eW��[�d��i�����v0gx�H�\�5���Hd�zi���ܻD�SD��4��0���t�M\x���m~������?�Y>m>�)�vg�p�.��2ȍ�i7,]u��U�Hm@v�s&�瀲5��D@�&4A�+PQ��k�L�g��I��U���� ��m\�8�Ѿ�ϱ�N���.��g|��b�Z���JQ=|�3n�/8����H�rV�#�����Q=�ޕz!��ge�D6�>f���[����@��J��dݮ[�x���e�H̨urPV��|>����]ɫ�'��MR��}K1�!emR[��n��N�k�eOQεU�ӎ�U�H�c]C���!uٱ.��b�ͼ��#��wj*{j���2fͺ�x��k�6ِSd���.36�sx��W�v��A�`��qH�[Y4���T������+�R��hD��ee�v��i�J]��Y3��u�lN�e3ĩB��˳���Mi�b�M��hh����)���)��H�{��Wk���Z&V�HM���̇�ܗDue������ov�U�[{H�co0���V�A΍�2츀w�-���[�èk�o_U��z����	
��oÝqE�o�Vϩ�3v��7���C<b�μ�iؕ�'�g[��O�
�����H��y+�lnHDڈ��ݩ-��{������a�d3���x���Zy�Q<�]-E�;3��K=,-S�a�jpӨK�����a|j��!��o�dF��f�)>B�}R{���&GM?]�z�^��c��U���P��������ސQ�&VOo��dCWs�f��ӆxHw�ǵ�u�o#�}+-?�Z4�|��:t�\��
�]W��K䰪���";v@~�U�n�C�%��ɐ�!�t��7Zf���!Q��קi��ē>���Z��v|��u��ZG� �Rƃ+;�G�},燐�2�e�V�3Z[�h}o�6U{v��~Hp:9j26j��۫��[�s�4USo���j�:g۰jx�W��>�ى��f ᭢��žJ�����y�'�s ���v��N��y�t�r��)�\u����(���O��HuEH�1]��koA`v�]�&Gf��e���u�4������6k�Hsf k+&��-9��k�/��(����,P9Ѯwzk0��Q�-Vn �~��n�7���l8���=ɘ��XN����j��驹�G$�AuЕɥ��"ջ��Yk��nU>{�k��奵¶��/^/�dஆ�@K�v"�&�R�9f�iY�C;��e��l�b4L��m��;4u�����Q��!���ɞ<�o�����ժ*�-�<�ຨ��9���qe�� ��'���y�l%����T{���S^\�Ӽ�װj8�n��7tF�/��M�k���1�m��٦Gg�V�h.KD$�����q�E,�RK��m˽��[1�zn_�is��&��j9MUbȘ�J��{4��;nw$aX�y�n�e�D>��B�Ġ�<+}��w�7zv�r�d�i/B��Vxwb��ǯ�O&ސ��cp|w�W��=o8�7�z�u-�u}?Ds���ue�j��O�N��c>:���}^�j�������>�9اF�/aY�fg%��s̵u�����,�p�|d�Ԗ�\4��PGr\��8dݏ�y���S�&(P�Q;�v���xGt�~6�����DqnN��\���_h�)�*o#*�`<��iky���b�^�+`/ �]^��[�_��&�he�"�����/�+tۂ{�,_��o�_��5q�<d~�~�|����}�1�iO�r�6,���;����i�b�&+f}��Ώt]:$Ϲ�:��g3�Ļ�9
�{1�K\*j��<��B��qme�ܯ$�#�Rf2���bg�|�7��_�n���Txt�j��.C��J�D$E���k�*u7�Τd��6)�D����!��͟E%u�9��&�qQUEXmԌV�-e����-9�y�J��l��K,Rpg&��B��Ad���NP	fR��M�{���n���Vp�B���X�	:Z�%���#���+���ٹ�Fل�c*��l���.o���W��y_��8i�D�"�>��]	a0Џ6�m������=�N���v�{=�6�l(�5�`W �.N�3,ֹWm����-��g¦��2��1��K^���.�A]t��岶�3Wt�\�ni�(���*�M��i��-���e!p��z��Uڌ7@yLw�[P��ܓ[9e��w��F�� �\�b�([�u�Pv���k����sF�4; {���By;�9v�NgMCh�>mP���r��(o�|�#ܓ"�_�ϯx��R^`W���ks�|���eKܑ��Kv���!�[v��!�#{���ʪļ�4�]�t␖�7+D����E��^ų?y�;gD���hL���wȬ���B��U���q�٘L�z����[s��OF}z �y��2 ��J��;Lz�s�xn��֞���7\�QM�Q��!OIT�{Tᷚ�
�aԍL��R�P���jUc�e��sA۝������W�hj����) {�w������1�UV��W�<]�?+n���2�
~�Lz׬ց��ֺ��KZ%���0;="��-v��Sz�`���5�[�$B�L�7���'����}�{�q����6�l��v��,���ŧyDmr�q"�����3�2C��>5/���u�6n�Z/>�J�L�������;Hf��n��<�o7���UXy��%�'���w��M�y^�����/����dA��3�:���!.��kL[}F��"Cp�)GX�#S9���ը�޽�f��h���Ų7>w��ܭz3.�/��K^K���������M��^�K$���>�&����\XY4�U}䢧Eg�(i�T1[���>{�c]/*B*�3�L�b��646c�?h���P��TGrH���k+(���n��h��6�0Sf�K��u�}��˳��j�I �莜��)�o|��(H��>M��ٜ�#1�h@�ukqs�۳�ͧ�c�l��⚇$e�.63���Y+�3�f;�3���,Ԝ���l�u�m>u���7
 z��>�JA4��y+�lnr�noC]N�N���A����k�7%_@kqooX���j*��<���W&�K��U���{��R�6�:�H[�����/'�_w�x��+g��{?�HCÅ�ꞹ�{sZ:gڅ��Ëg��,��G�I��H�;�os��$to*J]��Y.Dtd�+s@i��n�
����,~Z��ty�����w�w���聳����f�ZQeun��Ծ�uvY-�Hv=�t{��.LѲ������R�\��E>��w�3ah�v̫��D-��[���$`��n��#(��X��[g����ouR|w�J��p��5ٽ$�G{�e9;?,�v|�Ն��iy�@�&|�7N��,�Yײm!O��3	Ϋ6��nτ�6-�n�n��{�'�gp�P;[+'vPm�ͨ��\^�4OCvK�hA�vU�:<31<���"2sz���k�'h�?a�pX����'#�f�t�Oz�Y��O9��vn���t�<f�1R��]��Ϋ�{���
R�ݠi�]���bG�Xy�� �殗']Y؜�ӎrݙ����p�m��mm�dڧ{��<̕ߛ��	����٪k��ك�Fn3���(.^v���Y<V+��bpg�L]�	���8��=Qoh=���wTj6C�,5����JN���5]���a��r�@�ˢ{=lB������k����֝K�9�*]���mw鸕lU4��Q����k�N.C\{�Sl��|��wh� �����UA��n��AV�?����ݬ�ʵ+�R�p5�kB����+nV�V�4�t4�7���}��q<����\)��)�nuҕ+-c.��p0{/��P���q|)��뵴l9���bT�2)�]WF��2b�u��QmfW��۠,ŉ�{���T�z�z���ވ�E7��<S')>�߇*�@����16�����yx�I�u�n�өCm�����c��BZ�ќF�͏l�v�j�LՌ��{�\�]���Y+T�o@zQʷ������y��Y�f�zV<��N�K�Ʈ��8di���¦<�*K��kvu�ڛ յ�\�\Ӣ��e�D��nel���]�p��̋���W][��o��x"h�A;�C�I7hެ�h��U��el2+rl�DI���%u�#�����v�Ǒ�b[yb�wƶo\d��֞��������J�U�T�h�����={ZM�Z5���;��T��G�X�ׅ�֍b�{`u���������qJb���J<�sk{�m��:����Ơ2��-;�xL�V%u)N5�����T�U�Q�ҷn�z9R���En�W��/�G�u���Ԝ�g-�ƨ�3x r�ә7�%5l;c/-�J��o� 8�����[F�}�]=Hɼ˭��Ƿn��׵��PE��;J�ު�i�N�/��߮�\�k�;)�ࢻQ��	XF�6��� �w\	��M.�����^qˡ).������Ǭ��2�f��9���O_M
��m��U *9u��/">���6{����;�W���+tpZTy�ͮ�&%F�Nw3�Ack����U�z�ݎ��{�03X{*m��j����UV�vPĶ��\.$���B^<�,G���.��|XD[z�<蘭�)�-Bn�W���r/U��v��棔���ʼ��.�\���XL��l�j�8�VG���aXً$ضv7����B>�J�����zFgfB�d�Z�׃��6��s�p����{8h�A��]���f9�S�Rڵ��M�1p��p޶�r���cvV�� �yxLb���{��ﶝ���/^Dqj뮷5��-��Γzk��$�}�*�����/}���&S��m@���{b/�A6$�#C��A2�Xق]>�ʕ��Rg�Ο4+�V�N�nmf���m^#F;{͙0ɮ�B�V��ff�}��ٚ�=n]*Z�H���S�`h7}���B�G����X0�����0:�(5D�N��IT�ԍa�7y�9;%u	�&V+W�z餞�9uҚ����I��v�|D�:<E�%u��\�b�z�i3������"�D�n�0jh<���������4�:�!X� 2�7��/u'��t�n��2�n�ޙ�:�N<H��:�=��Wu@�U�e�;{k2�� ��7�:'=y7T�*�}���$ �@����'|�s%��9b�ۥȓ\�����L�]�$i'�]D�2i2^u�K��L ��!�����r�A'Nk���G�ڢ��2���.��L�(a�� �ˈ�b������̉N�đ�ܛ��t�<��@뮅&.s�0��H�;�w]���E��d�;�c"��I]۳#$�۵�O;�9E��w]˩$*��q��u���]	$��}W�HH�����$K2�����&M��%���u+��dy�FQ)�׸P�Y�"�X^�f��۩��!1��g9�6d��n�Mnv��vRAL
0�As����M���I$	?x	j���}X�+K`πR��"ů3Nâ�<��,��ք�F�V=]pMj6�ewv��lt�_[�ڎ�d�#â4�]f�t�������b����_w��w>�����RK��V�=��:��z@��I������5�o[T���:]�r���۝�V>n@݇���^Ƕ��n)f�}59[�z:�����L/�y���ܲ������q������k6d4�U>7�VA��}4&p�����v9jʳ�s\�����`$[ѹ�[����Y�Fk����lֆ�fY	�6����,��j���A7O1�/�YUf��~�x�K��l����%�3���V�w�n�:����y��N�����t~��F�`�����³>��P2M�]k�j^�3�����q�,�����˯Ie�TRf2{�ٮ��?��0�y��x�9>���ɦ���`^���L��>�Ϋf�r�X�q^>�ү2Ě81�=��&m���nLM�ӳ�໔L��
;I��{u�J �=YQ�Q0Gs3LU���O�~���M}�wD����-�pm��B �2R��&���ә˺w�h��5��w`k���-}�)��B%2ws�Q+��ٙ)�/:�s�zNѩH�Z��6���Aj�0M�gr;x���7�����P���??��+q�X�W=p�V���S���Ccm���˹�|�����g4�t��y�[t4ח(���� �u�a��c�/}U�MS-f�N��v)�@�ʯY�A��e�|!!��忔��u�d�M�^_��v�~���^'����t��+ȓ�S��b��[h,��ggK�e[gn���}�b:��X�I���X��0ڶQ^��a��V�]��}���۴ձOcU9@.ռ��W�F�Omj�f\�鋗�e4�ε���.@70��x�66Ҫļ�4���_B�4�z����LJ���S��7I^D+υ�[��B����V�[�i��lѬ����ۜ����Y����{��^}�)����06�d�Dv�@Tq����Tػ�W�����;M����؋gz��Ng��c��h���w#0Z�2d�n�������ư����Ws6z��W=�pS��펬���٦\[��Xs��ӣ�3�PINE�텻��y[u����L���x�Ykk�7�uqĂ �o�Ri�[p���9�-n��7����ǹZ�Y����8�}�up��"ީ5�cv��vk߃1l��X���������~@� ��<0�p�<�������6����\���b���n�c��#��W
�6��j�J�Vu��_x�m�,y�D�*'`��V��-�9*�C��7�亽�W^�uB残gg�_'b���&�����'|�\�$fP��}fǆ=�v���&��c12��-���6#�T��ז���%�t]��a�k���<s$nn�ڪ�n���U 셐f#����a��"�/ɞ���3",��QF��*�fH*��:�/t��{ic��镼m�l�Žtn�
�Hog{������D�K�k�7�mė��t�{��*�j�c;�Y�U�G�;g���s�W�"��f���F�D�%�@���do�bḼɆT���?<��O\Y�y"eqA<��3�{��FI|w��_���rU����M����tE+�Yݜ�}�)Yq�b�>냹H��`[}8���l�/�R\�f�)^�L�_�=0��It����=o�T�-���{�| ǰ�1��o�S�[�B�e���ol�v��D���?7rx�$3�!���� m����Ljެ�3ks�z e����ѰT�n�Qt��y,��=2ӯ���n�{����WGoWX%�¿Cm$���K[����������wVZXu
n�އ����Z ��^�,�+��r7�F[����=Ȥ'z3�Ӓ}ŵ��+�큪U��6(���!���ڛ��%�iN�W��1'd6�U����n��.'Y4jq�۰�H��Ϣ���V�vvƾ/�����t��
�!��q���De-��K��,�)�az+nZ�oh�����˼5����4_��`-��:�#7�5nVAL+@�d>��l���#q�S~;����X���֍�>ԎW"6y
�ak����]������
s�w���=r�6���~̕4ț�9UZ��Q�d�Ь�П}N8n�
�WB���<H��Lѭ�e8�7�IS?k�}o64�,�ǡ�}�]��Vao;ҋ��>�%��**8QKG��_U:�/�s(�[@�	�hP�b�n`Ѽ!��?E�1u���!\�%�Q�ĕ膲�R�NQ�c�u�:@�r
$J38���ֺ�t�⽔��B�]���fz;sw�!��SxJ�&��Y^ₕq�C����υ�w���'�ɥ�Ӧ4�>��G�Xn`�M�,�Rî�w��֔��,��-��6���C�������Cz�%�D�h�j��l��o��u �{�veA��y�y�b����JQ�߅��������>��XX:�M��a���p.�{ݙ��Vf�[�����e��jY��%����Yř��v�p�ð�&���}m�;���.�V���ñ�.F�R��F�`�����'q��To����1p��7�:�����>�)�ܲ�hO}���X�_k�}���5^�y��͎��Ĭ����uWrYMgX�)��e����F�5��uZ�~��:�d�$dGY�yJ|N���Y`�C�T^�KE��չ�z�=RV�R�����������p@Xf���Z@���ZLыu*>3�w$�:��xVe�
ٱă/����ܶka|㝭�Է����&h6z��t���s�j���Jj�G��@Ǜ�|�� �
V�Έ/7��l�7R=߸�s�+qTJ���w;�R���W��&�ޮ&>��޺�j�*�I��9�#��_��s#a���d��Dr(�P����*�uѴ�z��n���܉��0�Rƙk�&{�5�t��P���9���?V3u�����/2c7�%��AV��:ቭg?�>n��-2�]�Dt]�R�x�M���b9���
h������Zm��*y	�8r���`Z?J�J.!ON�g�Lz�+�;�^Y'kGF�Ul�d�,���;y�i��v]�+uБ5C���~V�����Z*oj���i�4��dg6��^�w:V<
�:{M5�M<�S�Uy�������;�l�mC��H(K��%�
=�&�Q��9o����m�SY�Bn!Uݭ��ݕ/���f�{CrH��n�+ ]Y]4���݆$嵃!��u�{��X4u�Nq|��
˄�o�����zW�F�7$�d�t�.�ڝ^�FD�9�=ۏ���Ypɋ�����&��x��i�7�����T�*�/�����f\N ��<w(lIA�8���1�O;�d����ېX���E�dH�ё�(n'��]��g_pY�
�u��f����{m�����zy�tg�h�|��q���e������˸B� \n�S���^�-+t��;]�٣��؛�7U�?\D��|%��3�!�͑�"#�c�Mn��Ȭ6���imU-U<�n����*�z�M�8s��݋+�GL�M��+�i!/��,w� �u��:���ϡOIT�@�j��6�Cb�,	vl_���Ɵ�)�*��޼�Md��i�v�ђ�ϻ��^�32a'a�2�����N���D����[��sO9i��^F˷�Q2f3�����3F6ُ���&��̫��H������DQ��H�E�D�4�~5ӿO�Y����U�C1oV�W"�oX9�N��Vc7��!�Q�St��Me�[R�&}쩭U	C�̦=�b�vzZr��I���stv�P�n���zxE�:Z�RX ��o��!��ߵn���o�NM�#�5�K��d�5��*�$�l�'��I1O3-Ĥ�䬎	%q#N��z;#yG��諙鋦�ODy�)��91d9A�;nܣ�e֤�g&��a��R틄�g��Y����Z�ݛ۷�"��台���Cy"l���m�Z�*�n�:�^2�w+J9B�g�Ԟ�f��wc7Gft��2���j��Gt#��"V�꺹�\[TV�FvPY,��>i�]a9+W��Y��m�ӡ	��R5�0�r�ݾ⺸�-n��Y�k��
`ּ�Hj�:'j8.�nG��6ћ�PF�Pa�u�V7�]��;6�$�0��ͻS�~�;��ս^�=i�ʇ�;Q��Z�w�^.����$�'�)c�GT��/I@�}מ[	og�K�uW
F.���N�qZ�z뺐�R���s#��	a�)��<=��_8w��j�g�ww3:Ț�1�q��m"�#�-
錰;����%-O��,೷ܾ�,Z�H�o�Fk�Ǌ���ܖ�'[��N$�0_D�;��V������nq;.5۔>ِ +2,_G�Ϲ���VUg�3�_S��z;���)#S�³��o�k�]��F��ˀ��(I~�Mx����@�yC<�4�V� �5{���Q��yɘv�&d��fICp�R{�f�Y�J�:�T*Z������M%ԁ(4=8J��%����mT^95T��g��n�(xI}#�\�2��Yn�K�,2#<0�Y������FX�1��D��ѯ�Me��Z�i4�L���=�Wt�R"l�^��]-��ۃN�:�:2�P�m:rbN�f�B�xu�,�]\��:`�q��(1���-"���1ٓdBC�=�Y��M��y-�*����f<")SQKY�`�ylf���a�t^��5�Z��R���@��5��YC�
B��8����	�eT��LC���E�]΂-����]�oqg�ZP&�����0�W����j����f����zTw,��\���9u0z�z�.Kh���S%�5�������ۻE�ky!����Mª��sQ�3�y�hT|&���=Z�Q��.��p�����ךTN���Σ%�����o�Llq�8�K,7�p�� {'A6�r��Y]
���x,��U8�.Goǃ5�`����=$�et�n�4R�>q�S �M���`d!���K�V��C�g�}
��]ʹ�v���~9�Z�ߊ�}[eӲ��mn�w�ߒ�X���E�G"��jo�6}�Lt�f�/	�y�W;1��y�vQ���Ԡ�&k�Z$zycz�m����R�j�5���CU��fH�n��J��#7�G��}Z��22ڟ"7|UƟ�$��;���x=�m��ȈԨL��ߛ�,��bJ���b�EZ�n�an���u5DJ��77Zj��g�7r��N�u+x;0��e�1n���z�cbgd�{�a���@F#>����O:���בwy	�نm��H/�ґ��#�!��6t�A�WMk2.����ΰ�yGOD�ʹG̿卣��-@�[����)0ݲu@��.s��������2qF���{����y�V��DX��^A"2�TU�һ�Ŷ.�K�\�f�>}qj���$�dy�*�)���YԹI8���_�m�Q/<��3	�T�mw�b�������WJ�\�\LԲ�*���g҆�=�R8vfh�uw�@9;�*�Z����v�3��.���� ��p�9�X!�O�k�{K>�]�H%�wЧ�-��掳@�5v��9`���r���T\�e�us��J��i�Yf����,<Eue���Ж�Y�7a����M��Bk��zN�ak���:㬡{u��;E2�RQT��r��;��;��۱BC�m�{�4�n��J\,��֓��
�ќN��4���q}v/���©*�:#	�ھߦuj'�Z���2�(�ct#N�Ǘ��y�qb]O����FηNԮ��Ek�]2�u̜��L����x1S�S�Cc��2E�Y���]��HX��n����!�����t�7��8AY8��ZB���z���c4H���������l�M����Y����_Z;�L�I*r֋��[�j|q�;��S-Ew+Kn�ç��6)K�5.�5G\Gy��I�0r'fŸ��i�˱�l2I�����ξ�[q��+�2�[�s@���%f�%�r����`\|�V>��j�l�f�P�9�ވ}��V0�h�]�)���԰|5�`1t� fD���Ɋ3��|6ea��SAr�B��K#�=j<u�+��٣��p�����a�1�J=�d�1�͞wW�[X�㩎���b�f��/��OW0�j<H���N��V��#cVx\I�ɬ���l�B��sf�\�_�'�N���Q̘3x�����J�&�A�ү+*]ԭ}
�, wv "i��]v΄�I�ggXP�1�aOz�[M�e�W�D�q�� G!�cαJ�b�dUyS�4*��L��iM|j��p�'���V�u�C���%.�k:v�p{!	���,{���kR=�n��x�����ueܝ�[.�r�L
=�:�#���Nw�K\�����0��B��
ү'��9tf�Ԛ%q�˱��A S�ܚ��QcB��B��e�zcL� �5^Z�tJ)�P�n���oV�֖�|��v����Ll���㹂��fo@;I��7�f�����s&8�	ե]��G'���b��65X<rN�U�U3$*t��a�ޭn�a[�ԛ=O�	�U�)
3N���������A+=�&h۱�D���Vzn�k�9�f����#����:��tȇnn�35]��M��*�vj����U�:*���"U���9&3�9�ig��+D��ƌ�+;a���Mu�J������|���>�*�v���,�J}�L��R�盛p�6�K�V��]�`w^|�*��5]86�6��i3�J��r��l�̆ov=5j,-^�%����e�;�[T�u\���Jinn��ۯJ��-B�u��y]����FŹ�v�Yn��U�� �l��i� �<zxEyN�Y�%{w��j�O
��[(�Yv��s*���f����X(VP��ŷ;����
o�ucuc�u�z,lK��=�r�a�弙�m�I���,V]�	�:d4��oa.�b�N[3;[����4}�,t��:b��{�s��(Lú��t���.�$I�4�E5���;�D��P��HstY"#X"AM���&e �dfCu�DH�a$]��@)ewbwWbB�S(�)�����]��D���'wF�L�$���>s��˻s ��d��)&6T�c��%ˉ�����Q3�뻠ewqΐD�bf�2�;��E2`��L����b]�N�A3``daf���%��:��)���I9pƔL�����������20S1DZ4&ɤw\a���Č@��FH�cHP���`X�,lwu���ǒMdJ�\ƽ���n��z���mX��1�${s먥JȾ��U�"�r<��<�V��=��J�v���e��0�B�7�]Iu&,Z��f�I��g����z���rJ�TV=[-t�[���Q��=fmm�0��M"Ou�ȝ�#�]��r�h��V���̶b�1~���}K�#-����б��3R��$�;3��]Y]4��v�搶���3�T�[��KF%y*}}MW����x�䯣s_c@���>w7t
���Hi�O�Ɍܱ�"�\d\lm�T/�z1��4�;�5Y�g.�n��6T��u�D�v3
�9���Dk�����aC���3����Ȯ�x���ŵ+ݾ7��"�g����!��uGj,�MeR��me�zUW�{i�$T���=��ʴ��Q�7�lg��T|ok��MA�yW��DL��d��=t���h����5@[j,c���s��o�P���<��LP�oN{x�uy�k#9��WY=j<�p�r�C ٺ�cnp;0�F�$����
p�C��j4Vu
ޘ�+�T;�ܣ~u���{��������fO�d��{ވ���:���p|��*��x<y���82�F�2���DV�ê�m�ë�Y�����l��';���0ǥ�_;�8"o��y�ho��!�G�,ڦ���Zi�ZwigP&[oS7��/;k0����:���Tl���xD`������>�tm����h̇9m�>��q�ɥ;� ��j�š}7�-n[ۼZK�,t�=�ʧ�a�X��=��Uˤ,�Av�I��n�MY�E]����^�Y6�bUS~�9
��n��&�>�,�ձ��"�A��围�K{���i�ɓ̎q]����s�Qo����*���&��hM��T3s^�[6C��-��Ό�����۶�=�M^䈌�������P2PB�ꇁt�qD�Fo%���i˫����a�oIi]en�����{�����.���^O��Nzq��MaQtO��:�kG.���@�Q�wO��}����s>�n�#��	#amOҏD��IӶ�n���n�G��]�$f͂'��G��ҳy�ݫ�Zw9N��$�dAؠ�Kt^�[6x1B�][΅۹vӆ����Z1�jjs+rj�Q����7A�Y*R�K5��l)���ao��[�*o(��W�cж]�D��U�-���T��?�T^�U�'�+�28���-�����Ke�9��U�G��ī��x��d��m"�"��Ӓ;��؎բs"*{w272�͠y��|�l��9g�o��6���Vl�����*��ìoLjڋ�z�����6�B2�e³�/�n-���zy���]KW5��.}���x/����.�͸wVHeH�s԰㜖�T+Ot�_KE˵�yv��bsz�@&�HF�b7�
� �d>�Q�o1�&`-��qF⺻���K_Q�7���x�I��T}�(�{+���	�G���w�j8�f���Ƨl�0�Hۛ4yL���*�����w���@��k��a���z��f��=`������m��Q�4׸��2	� ةm�(NL\OnӼ�c4�����4-���kMtF��)s����� X������P[�5�"C�����b����!�k��τ�� n${��;S:ގk�l�{=���wĥF*93}�H3,-$�ݪ����)(V]��� �hNj�������*$I�����D=&M!5N�܈���)��0q�)�{�߽�f.V�-S���OX��kK�Y�{L��=�7A*ѥ�`��s��V�8�Hg�SC�XԊ��z�-�7�Md탽���ʐ����ǒE�x�����aF�%���+�E�k�籼��\�W���K��b��Z����QSo���ː	\&��w�w�$D}#���Q��>�;բ���6�ȭ\�\S��]�,'&�\�
�ҏUnd@�;���6$��]�.;��w�\��'t4S\Aٱ��#��kk"�M��8gEF��}V�S7����d\�}ӳ�	,��Q����"yy�U��ls@���ᅅ����f�f-��j��V�u�2p�h�9�Ɵ�RY��#�D�i���!�8d�q�=>n��^x[���.�K���Q�d�}#�#��8m�[?\I�Q�.�[�2�^�[����i\�ް�A�V��]kWn^��X����`&��<̍���$��ի[��Y�����p���% ����X(�t�h�y�N��^�%5���sg!����T�V�J�AF��TH��R��Y1��Y
uv�Ѝ*T���8����31��^�z��v�y�El<Qڿ��U��y4y-�)�����S��ݮf�o]ַ��/jU1dȉ�473�ֹQ�@�xRDl�j�]�dl2��=�WN\�;=\��N������u>�������+�	��ԯ���ˊ���`�σR�r�ⶶ¸W,��L��v�1���>\�f6�5�쌪���rg7�����#��;�䜲��x�ʠ
���Q�d�]\L覭��4�	�����ev-~'��[~(�Q��Y��9fD��#l����''�8;Op��d�#A�C�o�{5.�䒴�wl��+�(�=�׭:bbfss_�Z�>/2�3��#LT*�f�]�@���ty��9� ?<y�)��O+o��Xf��̳�C�u�=q�6ҪĹ.�B�ޅP��fm��ͩ���������{(�|�|/ -��y>{;�sU05ᔾ���N}~ߍ*��T �C��7�C��M'����pI�ag$�ZI�B�-�؆ܫ�lѢ�Xն\[���|E携iU7�q:?�/�+��:f��=A,�԰o��"��e��}s�	����VYWl�ٯvg�&[��0Y��*��b!��_�w�����71!^��坄Kny�{z_����V�[kw�z����5^K,�^+eʍ=�	�zF"�>��Nd��q�����˙���WM�ŧ�8�3K��.���H�������=����rm�'fߗ�<�E�:C�p؝ͫ�TP��W�׻���%��h�j��E�\{����?A��k��4��+3��3�vcw�qU"u8���R*����bV�����5!�7��O�6���D�UfZ�Osr�n�,�y�/_r���>�Ҥ�.�l�@��}�w������(��c��lm�zCZ�yc��R#�P0���nn�ڙԓ�6��흵��ٓ�swz��K�MP҇?+uc3ef����U�����g�Lۥ���(7s�8k�)+�k�]��'�C�mi��3��)kk9{H���J^U�-oe���rwE�P�[%	+�yIE�w��Y��̵�^'������;���j�y�zp���PJ��T9!��:W�P�D�&`��0%�<�C�Ow ɿv�:f�V֫�e��\��;�FZ�Pt}�M� �"��k��y	���!�OL��ꮯ�����N���=���j�͙ɲ`��"�8�%Ō#/q:P��я:���1����tw��#{^3v��N��-��mu�e�e�7E�nv��s��/x�.6��[{�M�̀6��,a.�wׅKÂtf>�gdy٨�w���;��J�J��]��}�4?�0C+���)
��"�qPk2�ꈗ�*���V�+�����۫-,2j5�PCr�Q1�a��+Ryy�kN�<���~�;���2/;�N����}HLj�؜�<_qټ�~�;��W�fpV�q`�B��ցQ�7e��휰�:r�^]�j��rgC�y��޾+��eԯ���}��j��&Vy��\4N�-{ �^�/��u�*��4 �k������}U����K���l-,}kw�I@29'��I��e#:Y�ជv9�~��I����O'm�2�+�X��.Zy{ś��Y�2��W6��%�9�W"�-�8��T�fIɕ���s�뼓)�E���Q�MXܪ3m����6��G8��5\J��om<3���dm_N��}�%���Dk�7;cO2bZhM;y�L*�؆�7ͩ���ץ��;eǎ�D������&'54Cg܅@i�4ө-����mY�B�9L�cR�[fð�!t���7�bZ'��J��S�<��v�EuOX��ێ業Kմ���Z)�o�t8�g�㯚u�k6;�c��;��12�x.���n�C�<�P�G�^QIy�<gsn��׷��o�y�6J}�3�@����W���S*��,�\�Ⱦ��7��ܽzV�R������~*�u�J�����ןq���p�����0�Ld�d���Bz�4ټ{X� _k�b킕��0
Cv�a�5����]�j��?�r��0)��~�{��}�r���m�wzU�u+;F��_���t�f�!����Bc`m���渧T]ֆ����B�Q����u쒞ކvE��.�a�.�<]�,��}��J�趺�l�5��&Ϙ�nbu��ׄ�Y	��󻴽+Mo�=��NG�,��D�}��%���ə�S~�u<�<m=֨*4jyJ�̮J�-�l���a����8�I��|(+����:��жԒ���urɧ'N�o�F�z��Gh-B�����V�z�a���^�����Ϲ��M��Q�fo)J~v��/�7��%��^*��ճD{X���4�{]��e�1��U��e��]�w�Gl��aS(�������ߎ'��Q���g����!�m�5�6j�����-�|7dB�U�{�wN6�=�qk�HcL��@���7��1X�U�\d,��:gԘw���y��HH��!Y���2i���E�C�1t��5��5*��2"n�e�δ�ύ�+��-�Z����۽�R�tl�:�M��KYj��L��<���Ki)�.^炙��'t�/UGô��A�	d�W���$jdEݶU�O����lSE���ݔ�B�Z�ϴ̜���7<jʬ��E[�l�X�N�j���gD�~����hC���L��0��(�c&����r݅�c_L=]������c�xb�(n�0�1��f�^z����5�٫}d	����j[����k���Ϛ���́[鲽};^�x[�ML���[��H��-�Q�5���Z68��0E�'i�t�ްִ-� im�%b&�o�WJ��`�ܜ��h�E7(|ևl����<�O��$��+2m�]�(ڞ��3������:�ͧ����g�t�c�	�y��9��3��p�{���=ܪ:���٥(9>(܃���YN���h��n66Ң]��M1���|2�sĻƺ'd��Ꮨ�5(����׉on\�Ueƾ�z�3�^gAւ+������1��2�Vt�B�{X7`����
.զ�v�nXpv��H���7J�<t�+�yg^"� B���̎��:\Ά�h�z�IdU)g��;64m1k�[(�}��13g�[����\Sԑ���4n;��Wiy��F|ᧂ���
��������l��U
�zC�_^�7����w�����ڥ��Yx�fDM�Uك�l۳�M���*m;?��n0�K�hDf��ZA0,g_զ��1Nkf���~���o��@��j��ۿ׶���6��u�[Q��[ko��n��|W��k�������[j��;m�]KU�MU�Mj����m���j�6֩MmT�j�MUR��ޯkW�-UJZ���{+V�KUR�m�R�T�UR���+UJUU+��m���e6��>[mԵU)��Skm��U)���UU)��W��U^R��)��S[m�֪�������mUJZ�e5UJj���]���UU)[m���S[m��U)��R��)mU)[m��uyUT���J�l�UR���KUR���J��+l��W������[e-e6�MYMl����)��Օ緞Sm�ՔՔڥ5e-��l����)m��]�)k�km���������o���6�mV5�j�)��Ț�����������_��������o����������������mm<��5����������_��_w�}������?������?���ߣ����[Um��������������V��������m��l�������N���}V�v��o�����k�6��[o���~�m�uߣ�W��ʻ�����|��_������ߧ~Y��_���)V֫m��Vթ�m�M��6��SYj�[MUST���UU)��ͩ��5��%UQm�ƪ��m���6��kl��b�TU��eT�j��͵j�t�ڢ�Z���g�mm{������?���kkU�*�*�*�*�*V�;�kk�m��������f���k��O�}����-~Ϧ�w��m}����m��kߵ�������[������?=�������|��W��m�����_����ﲾ���իV��|��Um���߳k�~Z��|���יV�����5��y覵j���i���~�v���^k�[��_K�]�o��n��꽵�k^ժ�[gݿ���~�j������ů���z������_~�u�Z[��ѯ���۵��[o�ʾ��?���kV-��+h��m�mF֊�*��5b�ѭQZ�lkQ�Ŷ��*���V�F�+h�ѭ�j�����kjŶ��֫�X��cm�cVՍkZ5�j�6ڶ-UcZՍ���X�Zƭk��mm�h�ֱkZ�ڵ���5�Xիb�kj�j�UjƵ���-m�*�h���Z-�Z��j����lmlj���jѪ+b����F�-X�h������~^mv��-_�_����v�m��|�迓������-��io��޵[kmﯝ�є��F��@���=��������?���[Z�~�ￖ��k�_U��m���_�ڿ��5�_�ߏ������d�MdG<�d�f�A@��̟\�o�TUT��(��D�
E}5[2[3Z�"D�
H
�!!*)E �E�
��R$Uh�R��T�"%@AU*k�p���-�[��J�mak1
�d�lY�Ě-��uڻ���v�eL�}޷�׳;gf�b��³`�Gs�Y����Xm6����k�.�k[�ӽ\4v��T�Ѯ�v�k�ݗl]e���%�r�����+X�;��Gc+3kl3�v�%�V�V��Ŭ�Z*�ɻ9�m%m���T��Ye�m��+�mJն&�   7.��C]�T�˕]knsZ�ӱ�ܰ
Ӫ�u�7s�Iv���ΪU�^����=�v�TS�kc��݄��5�m�Օ:r�]N� �����k.�t�Ms:��Abm�Z�ѩY����>   �� ��(P�@\�� (P�C�^p�B�
 ��K���CCA@��R�/v���:��\�vu��Q�f��Zi�{�n7]#��;�[�l:[P]���A����p�yU�l�m�P6�L����  �z�uס���j�n�nk�w����M�#qӞ�Щ.�x��v����n��m�ݙn�����v�.;�^�{K��]�ۺ��KW8[�7N��Cկ{�V�����:R�#�Sn�  �u�o��M��F纷mO@�u3��H����:v�6.��ێ�v�sv���	���mz[�m�(�\�9ճ�n�ۯ[ޮ�T��]3����m����m��춭���Z�g��  ��������=P]��꽢�t���v���汘z�u�wk@��7:]�-��k���%���<�tt9�v�6��iO]4�]����m���  �������ێ��T˶8�`��)@ֺwu}���mc`��s�^����j��^������{ڍj��ǡ�ηMu1��	$����fJ��   3<Q���r��eU��}ݬ6�.��;@m��zk�����<v�&�e�h����v�'���Tw-�x �^�B��ڪjڅIy�(Sm��MP>   f�  �M�  ����(Q���4
M�p  s����=�\  �P�3�ox��K�  {���7{y���D���el���   �PI�k�PP;���t���  :��� �=w�7` 5�6�  �( k�p �{�\ ��l��E��N���wgw7=�N�|   ;�@ ���  &�p  i����� ('N�  5۽�  =����]S tUک�  ����R�  E=�	)*��db41��PԪ�OD  O��E4  5OdJJ�L� �I eI!2�⟏�����U�~)~/��u����<�r����]w��]�8�w�}�N�P��	%�����	'RII	��!$����	'�H�$��w��o���0֌D��[[�r� ���n�@Z���6{��l:�j;.d�Ц�����ݬ�1�FPZs5�S���W�'�;�P�[*��Bu��SF��4��]�#��l�1fa!ա���×H�UԖ@`�t���NB���l &4��ue�XU���7����YR wH�D5i�v\��^�.��3�hO����4]����B�#Yom�X�WN0�&LY{7)���;���:�d�L�MՔ&�ai�	`.���w���X�"��P5��1���m"��z!;�����H0ݩ"jnf�i�IW��f㽴�h��y�o�)��1�1�K1Q�0��ە���䱟�:r�Qh�X�+5�:J���V�/n]+An`�����O�W��f�јh��*�ʴԣ[tm��x�r�&Wz�D]�Vu�;wt1���+L�9�PETʴ̑e;-�;{�&�
:40F<ʲ[2�K�K��f �"�����z��ww$u��C���<�)��~�YJ7��t pk��r�̒�ԛ�]6kb��)ju�n;V�z^�هM��,�O1���OLN���&��ZF�I�^;�sM�8�L@ɠ����+Zpc��Ƴd�SsLX7`s�	��֮�׷��� �uz�4ˑ��*��@����6C��;.�Q�Wm:�����f�ovq�� b+�-T��-���޺ے�sF���	BiaA�l�wVj���Z0&ّ*�/!�-�f����6v%n�ۼ'.hG)���Rm�kv�Q���� ����V/����wۘ�Gdt�Џ-٬��r
n蛬n��ѳ1-�/"�q!�昲8і�جв��,]���zwP�����i�Y#iI�bԮ���mkV�J�Ȯ��n�wZ2Qq���Ͱ(E64-��.�V�e�%�b���k���<0������
�լ�r�[{��5Z����R�jn�B^^�x]�j��n�[.�P���!����/m����YEJFc�2R�
t`͕�6 ъ�F�#PNϲ�Z5�VŜ���V>8B͹Q���
�w2AD6��q��ƥ�����BT��R�U��k^�V,��J�`����"܌�k��8���@�?�&	��-����`�)`J�W�@��Vb�˛�Aˡ���8憁�^VمQA��M߅�M��X7F�u,�PV���D��D:X���J�1Tj�h�6C,�0�Au�n2�5p��U+l!��qf�,�N�o�4�nޛVը���tk`"�M��R�8@�VF���.�u��Y*��UdCS��-���Vm晚I43/m�-�ݭxNt&M^&�kx���#�%d"#8��&Ƒ�N���Ԓ@��M �������+/`��ŝ���*wMn�ȫEe���IŖ�=j��b�̖	[V�[@c l[[o�2�ݓ���%��.4+Ў���ŦV�mUe0�y��Ѩj!�8��Chrڹ��B�M�p5ys@̉8x��,���k����mjB���2IR�e�c�.� ��!�Hf� b�;����<��懧4��c.i�Ç(�+˨)5I�Ţm�v0��m袮�q+�/2��P�`�f���)VX�O:��lYk��a�5*��Su���qXu�Lى���8����Xա1cVIcU�K$�4��f�M&�z
b����ڕ:"a�{Z�n�y��l9��.�B�R��+Zg�i���A
�Ñ+oP��iM+�l��n�#p�	�,�0hĞV�A� vbn�����S����Z��<�%jA�[:(s޻W]Zj��F	�'��k�4����oH7B�x�bU���̹��q���z�7Ҙ�Y���[�A�v�w�^H��zH�":�$��� [M�r�jt�Q	��9��%M�n�����Î�n�p�i;Tbː7IK��b�V��r�:9�az���"�-Q��Y[�P��c3j�S�JdR	e���Y�E�~ܤ�^"��J6�j���]K�N*`��̹�Q�lE,B���������'��u�y;e�nł3b�CV��z��{NJ`�+0��w�ܬ�K��#�jȺ��kf�x%�hGHv�u��l5�AdWam�L@	4+�m7aX�j]���i���v�.j8M$r��zF�P�e,�On��f��@+LV����p��Ѭk�:wIֶ�X.�:���TX�4wi���5Z�L�HY�i<�g��jڗn],��5�h�ʹ�b��'=�(]��R��h27u���T�cdd�j�Q��G��i"�t�V2�t�^�� �A��/B\��Y-f�6�
9�%CI�b���4Jv�xu"�Jr�U`�f��~����T�9X�����"m�7q��Hon��)���V�ZY�n��-���i\q�+A�-�#>���zֺRb�"�D�1eI��`X�	���
5h�&C�7%�8��"?'�.�c��1^@�:5�����l$��oǪ���{��Y,ST��h�&v��u�RU£��,��C��m��e9LJ�.S���ڐe�צ��Za\����U��5R��tN<�J�%�@2;m��
�̱*�V��G)`�ܧ��s,S©i �i;
���t�	.!����V%Y-��*�%��r!i:m6�$��sV�V͌�M�Y��Q�ptTմv",'Z3m�����p���%��N�>͇4]3���.��I4V2I�!��E[� ����U�GA�{5�+"Q��^��$��x�܋D�|��6��I\BY�[X�˩7vKW��	{�b���wO"�h��c%,��C0԰����,`4,^A��iAZVY[Ti�uf�{�g.[5L�`��J�@�n��V��V�	�{�Fe�i-��L�[���+6*u2+ʍ1^m��O'ڞ 63�PǸ��27��$Z(@ݝ�eMZTO(���+u�Z#Hi�b�}D����(�PƋسX�aV.��f#m�U1c%C
�5�(��)^H�n����$V����Q�q�"8ҕdc�#u����69Vw����6�
��Xb5a�p�E¤�,&�������J�����( 6��CA/�[��$�g�)XnͰ���z������z[�j�>�w��S�m��b�@N�yL"�V���
i%�d*;���YMcͻIn�E03bd�(���L ��q���1@���Qf�����%SXvụ�����QB�N:����dJŚ���81R�z�V+���(�oUbk�4�n�I����F�2Tz�wyf� �Ħ<"j�h�E�t���-饊T����\��:[PD��Y�r�4^�Sn:�0����7V�u��*�ݖ.���	��ãUZ5��P9��v��nK�	��J�"f����\f�k`��ɭJ7��l�Zj�S&�N�bV�](S��
`9��/�j�R���AQHm�{Yy#�mF���&u�]�Y6�y�J7	��*��^:Yl`��1!�b�^�P�(���ܽ�r�Z�C&�fԆ�W���mj�z)����k�)?�[���d�N�9u��%ݜ�n��R��5�^���O"t�*�@�Y�Zr�l ��jL�D]*�o�IG7%���U������lK����I1�����h܆B!,��f�[_7�p��R��@�D9�ee[a_׍<U/tT�"S��f�z �xHk�;�Y���/2+z�нZ��%P��5*��])�b�!
@�t.�P�f�H�m�MU�dzTW�:N�h� ���Zӆ��y1�uV`
C���\�y��,*������1`�Q�M��#lR����q*������z٥��	,;#W�Y�ң�ĵ�$
T*���,Y�)�enB@�ϖ��AN��݊�$M�ʂ�@m!����H�	R���b��;,iU�Qp�+J��MH7yG �ף-;��}-��R���M�זB��TXԘܫɗ��lDB�&��x��,���nn0�[*��
���ͻF(W�ƅ��Z�X\��D�U&;Tҗ��Фŉmág���i]�T�F֑@�#~�Įb�G^<L<��	����ۓJ�i�Ed8�f�m�n�h�}�����WOx�#�
��[. vZ;{B�X�G*�U��\"P��/��7�)�I�M'�DkB;g������%��	��[L����IԮ &�]:C5f�cm*r݋�Nl�N�K���X�;���2%�wI]�f2��n��0�4_׶�F��i����f��s*�Y�[��(�����a�#�1mve�m��n)	!��:��e�C��.��iXNۧH�c��k���j^Y���YN�!˖�IX�U]jt6m8�J4��Y�C��U)�ڌ�s
�AnZV�n#P�a<J=�p�]�g��ȧ�li�J}���%SEf�{i����,S*?��AՄƅ���8��q�٭�"҈���o�#V��"����j�+�{v-��̈��b�S{R��U�p�4�u�}����R	m�����	W�����R�MXaVM�6�S:��t�j�i�ȧV7UMr��2��&�ڵ���nY�QP�T�"��fؚf��Y�K*��c9ajʊ
�m��8Or��N�b;Y�)hU��jw������=Ҵ��p6��leЏ�HV�^�+|��uI�H��{��t`+�q��'���-�sB��N�,�ݺ�LT��DjdS��(B��7n�j0� �4XzA�PK�wM��Y��+"�f��PN�Gr�_`�ֽ+rMܠ��@Rp�pA�T��:�.�me��6�]e2� K����ݙp�p�X�庴#�F���T���.9����sR����-�3R֡,�
٤�Q�YC"�x�4��4�˻�#kK��j��`�J8���c���sLG��0"[��V��ވ���5P�@�^F�Y�q���.�[
&3`B�"Z���8�Ʋ�g#Z(� pv�ӡjR�R�J�)[x��N�!��Kz"�n��h�Y;Y{�Lt�mݻ�����8)�BĴl��oV��,��f�jX4�c��̠A�nʻ�2�B;��/L!f�D�D1Z�H(rƚ�r0(n&��U�N;w��f(��KV�^��S�V�i��h^V�2(�uL6N�j�0�ˬ��ݹ�D����Ҭ�Ͱ2?�1P�#�,���٣uTݣ@i�%��h��As)�ͬQ36��4kN4PVoQT8��Щa�mM͌�m������&��5�7dZ�-�*�-�rn'Jd���@+l9�fb��,`�iP@�����x�n����� � � �Ư���XF�{���ϊn儶B�X�bx#�khRI8���R��5`�Y0h�׶�%��Yq6��x\�i���-�8����kZ�*�wv�P�.	4H�Z��M�Hςͭ� u-Q�f�lD�zi�,��3[L$lk�j���Lԛ�Z� �a'5Ә+l�9f����4GN��[Xq`q&c����b.+8����0S�;�S��q6v�N�	���4��^���UiYI�뒷Q�b+�S��n�^�m	x�AB�����JJ���:�ˬ��É7�ֲ6^n2�-�����8�F�n���*Y�*5�މB�!B�����ƭ�����+
��k��]�"�7N���^R̍ht�r��.��fl���p��V	ܴn����V>r�$��HJzM��w
�a��oVH%��Kr���ˡR�QrK��!��m�y{t����z�qj��a��+�bt�f�8���a��8�Z�1a��H����̠�0��en�PI17��d��(�yY2���m�f���n�%�����B����j���g4�v�� Β�7U&��{�cy��!+�˅b/v�5[�dc��VfeS)�D��d@ ��&�bUuXCS�wv�CM�t�L�ё=lfn
��c�J��jMwo�l�	B7,����qn`HfJ�.�l8m�q�L�7�^6�NSI�w��"�a(4�׊�sS�Ou����V�2s5��2�vLI���*Ԕ;#j�̼�ò��Ô�ֈ���H\U�-����z�ܖ�R�P�ұ+(Ո�t�W���!�1F���
\�C5�v��S��L�x+���!�2��3�����Kr�
][�=�C�[+jn�j�٭j��-(�����M�vK-"�E�2�c׺&�p��tncjX�B��<
��e۰7sT���aJ�4���I��a��P��)�2)Vݹ��앫��H�[�4��ud3xJW�Ef�xֱNm�� u��0�R��m^T�чl^G�^�d�.�Mڽ9*�*Tԥ��^��	�a�Cj5b�2FQA��i�)ä�l�6r�fc�j@/�t��R:Pt��z�v�iawY��Fb�&��n��&�4U��_]�l���R�1h�Ghb�1A��a9d{Z�Ũa�hS�6��ȦLu�K4�?3f��y&ؤ��޷n��jܹga>UlSr2�V��m,k0+��c�h���@U*:����f������)���j���K\	!2��ֲo`e�ۻ��Ӕw.��Ԙ����2���r�`;h��0���9t�EM��oM�oF�`|�r�W�!��F��!�����*�߲i�En	c^���ql�����`�5ϲ��LH��Ɲ'OBx�b�Z�̷A̖�� ɒ[f��N�f��u����(h�ʻ�5�;����n�L��D)e��	Z�"xs�I��F|��Ƥ13���cw�^���B����A�!��Y��g7E�{j@t�<l�������W�%N)�[�Ԕ���g,�YT�ka�Yb�9F�Ӣ
��^`��,���Lf�QoQ�M��=�Z�
Ϊ{w8�KZ�x�-� �)����)��F�q�ꀃ�a�)ť3Wvs.4�Ea� ���֮](�;k�9$4l�.g{���'���D+�z����Q��R�r��<��E��0�GfM01Rzsb�L뵑�y��������ɒYI\��>{��*]�̠�i�VT:�Y���`Ό�I�]��@&�m�.��q�a��3��7f�i���"�^��E2k��]^V��ޜ�S���n��k�\���޵�(tmg1h���5��F�=�s3Ms��j�h���'5�}��E��S3]���!L�:�j=������*��*`��5�8����T�FE��[b�VJ��z�-{u���"`�����k�\��*+�[y��Z�u=�{V�Ǒ�8��5��pㇻeZN�q�h������)0��y�G֨�碈��!�z}��S	�zn��g&��fd��+�<�;t��VrPQ���{qqvI�wRS�9�ݵeAh��y0\ۓ׷���d���t��8�˄5�U��i`\�N�kIU�I�&���8�LIj7Xo@H�xFS��Y��һ�rm>�,�Vp�}�U4�/�a�N,���-�V��|%� 	��T�.������� HM�D.l�U��](���wu�m.R�*KKM�A�eX����}0�7S ��0v�2G��]��y�,U�b���ҮG���c�����6�KrQی�cj|qKp���D�/�ܷ\unP����=;Ʌi��o�d��Z&��FY�렘�+�.�R�{�_>�u�t�.�Ţ���i�����K0umA5��'�n��b6��c�u{|��e5�R�m7�^���mr�ʗ/���jf�W�M
9ue��)��z�+��EԷ]l��Jk�-�7Vu���j'�}jXRg#)^��ZqW�*pAՙ�a
�;b��V�"=a�5�d��iQnR��5�cK(����FӴ�7K�ܯ���b���j�;:�,te�Y{2�,�hȬ�O.�Tz��lj���
���*u>�-i�V��[�g�5��I�u�hI����`ۮ���{5�獨/֚:�������j�wh��f�{(n�*�*x��7KA�6:m�^�|�P��Hu��
�q�Xhdp��b�
[�g������Q�Ԏ��ZA����V��}Ed�����h&h����O0P�p5d���*ˣw(.hƈL.T���f��:�������/:�{��x9�|/E�����91˥ݗm,}����b�p��m-Dv��=���w�|��
mp�"�O]��l��e�}K�;w���Ps�}�w!{�n��u�V;I�A��ږqY57��aB�����v91�g�TX�֪2�S�*3J�)��DR���w\�<.��"Da�-�3��srJ�yv"
��8Ʈ,r!r�,)z��wv���P����]�� �k'!ϳ2���q��\��n�@r��� ��ڵ�S�NsY �@s��:S�n�����#��	��۸y�27f�܆����x:4�vt�!�7m�lJϸ+o�zU omY�̅Vم.�k��S��nCZ��qOݩ�� ̸�����h��[J�SO�+���Q���4W��E�)f�p.;�L�]�ah6�]�=.�.؝s���Њ+B�ӽ�Ұ��e\�G݄+��}�(s�yb������ߏ!�#Y6½�kG,��!T{��-.YE��5��,�lT��@���]��9e�"H�aWk��^%�Y �9�oqT�.Yz����6�a�N��]R�������\*�ˁ�q�nu��v�
Q�3�*kM3��w����y2�`���劚̛֠��6�	�)�Y�*���!�� 6y���|k4�3i6&��묤4�Z30������ċ}�IFU����w�#x�IX;�K���v��G~�e���
�qvu��׽9PDDܳ�����Zޱ,��r����������5����pd�^s�r��y�<�k ��C]���L��e�xi�|f� m�0�8�����
���'d�غ5��s�ZM=tTV�lGȜ�]X�Hu����X�ˇw%4���Z��B�Ѫ՜�i3�O*&�uBks�JIv�����;k��}Ң�����k�!%�;p�6�>כ�dXΡ*���$z�cJ��TZV=Ҙ�PȻz>�f�>�g^��@[̛ǲ�II&.<l��5�ޙ4m�����1hҋ�6��W}ۨ ��1�k(��q��xw/����P'���m� Ȯ�����YD�jn�*��s�\��]Խx�C�w�]�՛��lKE��ԫWN|�:[h��2�U�f}j��.�%�����2��E��e�DM�1V�9��|�hq�>�wp�ڪ���DH�R�ݥ��_�'��7ws��B�q���Gd!����Ym����+Y�&R�J�&��t��fp�{,O��9�9���U-]�P"/�:���U	b;-a%�	��
�Yy�"��DCk0��&N�Y0����R�f*�i�f�ԥ,��F�It{��6{��4\�K��ڲ�TZ{�y�s�Aad�G�6��{t.�>#	��"/*	�1f��E�Kt�C:��=�.�gn�}�$
���:�XkYT���ɝ�]�+��t���׊�Yi�j�6��@Es8퉼�����C(��L�S�V���nl̼�އ��ձb;M��b��`��P=[�h]�J�Y7��I���	��*��k��׈�X��Vͷ(�fsK.K�Es�'e��V&,	�Q���G<]���6�ëN]*��ٟK�{������&c[��U�$�af���n��Tu��w5�qQ�=��ђ:�v��_ii��3oXVvd�+�N��)��ѯ�EY�qȗwn����C��e�<R0��V���1�:v.\�a0���V.X+��P�˚�Ji �)M�����w;�-�+���Nf���z��Ū)X��SS\h�W�l�miՎ���96r>�,0ĬI��N&*;/�ų�K�n�g_kʷ�$2�	R�O����%7�I[k�֪c	�N�w+���SN���{l�pîL�O�\�E�Ake	7����rؽ)�LMu�5c6���;m+�:�	�r�Z��,j�κYW\�pu��^��j��G���ؓe�Uwҫ��t9IƵ^�K�VO�1�r�Z�[]|Z�Ka���PgF����7$��t'E��*��ևPn�5�o&#��K�� �{sl�.��^h&wr3�
x��oE�WV��u�M���x����mps],6�>F��uUu*E������6-'@�rҕ:`e:�04��ɰw�r�L]=�:U_B�2j�2�e+s�笻;3= 
Ԉl6�3[F}ysss7����v�#t���9v���Z���S�LҲ%��Ȕ���A��{���i��R˘"Ӿ�S��vkv͗�ʢ�(b]WG��x�f�99r�V��f1J<�sR�[{[ͬvF���u[@n�mK�o�#0rCǕy�"Ţ��tmĬE��'� Uʒl
�(�Y�CG1][{�Z.�ᒲoC^�����ak5�Ӓ�jcU��J����� 7�	+���gr�2�s]=��sX�Y�"�y��S���'dj��o~}��t�:ž�|U�M�Q�8tU����L���-�XT76�ˀ�5fB[.�%��:�S[M�ҭf�nЬ]p�U�5�5���jt��Zs�I�C�n�f/�Gil'`ǧ�#�)��R�Z��SsI���E��wW��(Vf2]Z��[�Um]�$�K�W�r���+�/VVlE��!�+{��{w1Z�����}^��[�cE	1�Q��v�F�)tޕ{ ����}����*�(`���7hi�QV8���nAi}NS�2�9�RGp�9�ta�ŏ�;�!}2��!RI�&���we<#-�
�j�Go�</h�gm���e�kq��d�j��%;��B�Z�5.�bNݞ�����3)m^t�Xr$�l�:��+�p��K*d8��θ��¥oc��V�Wvb���N!��uQX5�*˾�cY9SM{��w��A�	��yNk4�G)s¶wXR_\�tc׵��>+HQ��Ya��|s�9�T����Z�}4�ƶ��G"��U5B���]��]o#wXc�\Xj�?h�1YPq��6�uSɿz��5=���(�Fh�{���f��/�]`��u���L��C�Q=��4�Y]�wҁw",�*�Gok��l�Ơ�����V�=�������o�n����t�絯�ݬ#�W\O,�=�{9�ʗme���x=f�L�$B��(���4��������,]��Rh�(��5�:#TH��g� ��򜷥��I
�������S����+y��Y���!8��z:�{��V��)O���UY�i���� r��R_s]��wڂ��9}�J.q��>�	X"��W�W�s�#/IFh �4p�~V8�ol�Uq����J�j�����I��)m��_t���nj�������v,�x{M[7g�>�ZZI��:v����-EUq��8��-0-gD����S�����5��5�UG�
��T�.f�B���dڜZ��@1Y�X��z�͛b*��)n��cW�#���A36v�^�.�k��Mk�nc*��Vr$�m�XG������ �r�9�b���uJ����V�]�-!�Ē���t]r�{��u�.�v!}��d�ˌ��T�G���/��gGet/e
�s��/DMl;塋�h�wت�:ю�VVS2��q�c:� ��9������5�5�c8̞9٪F���OS�EN��P�=T
O�)�8��@Dx��Z��9����.��!��4[Yr��sy�#c��8���ԠQ�,Vd�{No^���Y:��B�a8�n����\�$��1��M����$b���Kz�|��9�ڎ�렯i�̔3�)s� ��,G�����vo9ĩZ�U�эJ*�4Y}%_��z�F�4z���j-UR,�8�#Z��ʱ����b]Yن�l{hR�y�M�-�PQ�ݠ���[}[�1;�r,��Q��0��5l=u7ifWs��� 9f��:�X�7�Д��X���S��`��)J/�0�Y�]�Q0&�y�����L])0�)��M;n���/VlYCK���4eu���jS�»��m�xvl7ǟ<����R��iW��<y2�Ӕ�sB=t�фS�R �����vץ�j����2�9pM�k��t�-7����d�ǿv��8��r�A�k[]w�㯬(4���l�BI�ެ��pO�S�:I�p)�7����J޸k�!�Л5;��D7�H�kf�N�]��c�!�)Ssmn�Ǖ��Ѷ,=���U����%�;���{��N��m�ym�����F��m�p�{�6c��J^��������t�JDɚM���O�o��Y��G�ɋr��|��7��݁���6cVxL�p-T�k�˙�@f<Rt�H�A�`�<�w9w1�����UN�S|[Yyv���Y|e���W�W+ᒶ�����4����M4�,8�y�6�Ac��I����]��G\��,����_l{��q\�%$��`��@液	�-��4��w�l�C_@��[MvtdZOq�k���([�h3�^p �ŕyN�A3�4�u��ݽ���敬�FB뜼
�9J�u��U�j��1�W\�>���lr����Xu}�Ҽ�*%�[�lٮ.痸�G�����W�s�:~۴���!}}L>)��2�MS,<#�j���h��=v��ze�b�ov��6���+�J��$��fLM�rf;�w9Ju)���52�>�i��֪�UȺ��XF���)�*��o,u�ꜛL�4� ���}S�w��.Q#)�K��"�=���ћ�m��s�z��� �����QǼ�uC��ٹv"&"��!�hOoo�d�9�q�K�l]��6Rb%�](�P���uF�N�\�k�ܔ�LA�+�L[���vʷ�G/�c�P�ʶgM��m���X�[��4܎mW$����W3̺K���
�c��]�����Vܚ4F��/�#K����m�<�|O��MFkw+���|����%������.4�i�;����W	)'�0�.�V��Y�Ψ�Q�x��O6��I1��v�]���iǠ�ي&KJ%�����Zz��}�\��&oP,���ơ��z�X��zR>�U�/�Ԙ��%��K��p�}�����"�mb
Q�L�2�G�>Yݳ��ȫۅ1E̹��
�Ʀ�{/���}�$֩��V�¦��y��N�����:�uzz�mv�X WLvf��"�2m"�0q�ؐ���Ϲ������ڽ%���Z�-^;_0�K���Zj}���0�֜{�ou��}�1�Ք�'{�6ͩZ�=
оnWT�1�ڷ*��0N3��(��}��Iq
��B�.�g&�B��S	��7�^�W������K�ܝ�iW˂���')ոΥ�u��{��D��f�8�::�^+��9��M����u�	�8�n��X�uw��mֲ�Ŧ��|��J�,s`-BE�J�*��}j���f�����o��fgl�{NvG�1�6�Ns�c�MS�&qy���\��䓪��]:��.�D���V\��-�s\�dz��}]��z Q>��j���V��{��t�å"�Vb�$���ױ[5
�4]�.��=��I$	$$?$�m��~xw�?����Ci�P$�En���`#��7j�;���_�'�Dv�M-TI�7��\�����ۧC
��0%A*�K;�a�wn�1m��3
f��h�Eǧkc3VZ+5u;��qq֍B�s�\�I�\���gi,��b/*��U�:o�z�K���NL�Lw�z��[t9͢瘄���;r�-��-�ӫ�L�._g$	�����ٶC̊?�&�j�c�on�]C�*��7��F77F��RK������DTx��q�8�_M�6?��&N�ѥ�4���gy#t��UMβҽ�n҅	��G��2��v�\/núԞ����2N�醙q��P7�yE갸�6������6[�<��q}���yC�jx7�d�pE������e�B�f�ʶxʰ��[}4u$6,��BK��[��-֮��?�*�T-��N��B�Jo���uv�p�]YrnM�H)��ۖ�˰
X{x��y���7��; O~�#n��immdb`�#!ڽ�^���{K+��WQRUAՐ�i5@wvw�|�5j웭Ju�<e�5��4��1J'!�5��(c�a��9����]@��K�bGVբc7�K	�qX�'G��{�-*bS�o@��[��#�����2�kV��c��Fg���5CZ�����S+������p����fk@���w��b���g۸GZ`k:�X-�p֥y]�`����dꑴ����u���io������I2lv`L�4��튻<�U�w۽��F���Z(�aob`�òb�+�/�YF�5L��}�un�.�N:īP�+Q�_�d�N�i�d�;;*�r6����t;p��;V
Ќ��`ϭM]-�VV�u�]��od�ʎ�7�9�őC��p�#suL��ȩ�� �-�8k�U5h��σw#�Ì�D�%˺�ը�]+ܨ�p�vZx~$tW��@^
��d�!Ql�_jC4ġ�V�,u=��ɛ�����L��)A.�u<t�we]�Vf`�*DS˽�/m�G�L���;mp)�i�ʢ�75��HUM��U��t�b�vo�8\kt-�^󖷎X�M���
�B���/c�1�7Y��u�o��������,Ww�tx��|�Ř��D�n��3�<�h��B+4ؖ�cL|��1��:�Z�څ��|˭�ɦa��7#��Ai�go�V��v���G.�f[���˘6126��E�'<�96>(�@]�9�u���,c�\ź�f�Z���amtnevS�*�g�m]��DrvP.e��)��o�뢁���IS0�t����ƩgpՂ���
퇜�	yAKh�U��
ʶ�F�h��n]��M�R���$y4���s��L���Ю|B9�Y9e�s
�{_k�tw�w��dg�Jv��y�n˄T;�k-���o@���.��0���%*)��Z��9�ei酊��u�y���Gk{r@�b��#io����aP�pÖ�\u��hY�έ3����8�gb�:��%��;0�����S�Hl����>ky�w	��F�o\u�ZZ ��b�76��)rTm3{�{{.TĹ�h���*J�v���#���mA��u |-�t��{G)ܔ��Aۍ�\$���0b��ͥ���ս΋�2.�٫F[�zut
»<�IK^J�J<���i�L��Vt�$�B�1:�ٌQVv<Z��5�)m������r�&[QR�Q�+��Y����l�M4qgќ���ܭb=MrJ��6f;�����o��!H�ے�L�����8��^0���':m�
ˇmnRj[�>'r�z���]�*��-J��e��y��j�j(VǬ�7Rs�T�D;2'��)���$<�H,�+8��Ig��� ���y��*;����l��wʔ��=	lF\�u��::���<�[�+V��2�����&�ѩ�Ap��h���ִ��S�M97\r2���"��t�XRͺ�U��Z��sWJ�E=��[��+��E��뛕����w�ȩ4
����2]YO���B1|g�z�����j��F�w<�tP���X�Y����8Wjs�E�\�yj�ha���Z���[.��9E<�r: .Y�W]�a![�p�qC��-OE�P�g9��S�b�1C��V;���&ӣP���^�.Y;l�M7N���a�9��[�o(cX��\&H��N��X���ִ:����]M=�����Խ&u�}��=BYK+2��*��ו,-"�Gsm"/���GtlD{�-_&�޻1�^5Z��;��m9S��G�����<e�ކ�28��m�Fu�%�Ֆ������ ���!��Վ�CH�Tmo:j��gc�4�2�f�%#ˉ����aT0�*�4F��/���v��%�]�,�]���n⇥�%�$7�V\�������Lo�*	-}e�5��EѮ̴�[o��\�VQ�[0,����ӏ#N�N���Nz)����/PCD����f��PG�]]7��F�q��h��)�V�D��c�ÜJ�®��g��uטӫ1�s�&�F�̻�e��8ڬn`� �T�T�g*z�lq�ܛ���H]{���=j��ň�GZ펺��P�]�v�[sOk�*�r�΅��	�nZ-:�<f��!2�AM�ְ�Έ�5�z�ӵͅӅ]�QwZ�J*�!�Y��U�cGE͠����S�3��1�,�Θ��V����k�Z�r��*0>�ۡ;��Z/��ı�Z�$Ž�ф6�	��4�x�1��ݷOut�NXb�;BoFj󘎺��w��kՖ�nv��x�>B��
�7:�E7����"'��XJҫo������VcP���k/��/_��F�ؕ%����y�ΖJ��h��R��wƓ����sn���ys'i	cln���9je�M��=�-U�LX�NM�p���oH��3l�ʩW}6 ��=VoUs����wdY�_�����8�&��e��)�ge��.���aWe�Y�X����iC�h����^��	+^;&V�՘�
�`�����M���#��:�Q�z��R��Dtq�X�x��f[A*��:Ӗ�=zm��*V;&v,SMҐ�n��K�
<��${+J��p�$ec7$�v>&��V\E��˪r[j����G�4�'7fh�9�:���t�cjrjو�|wu6�j&���U��>��H�!|�@�\lm�;���آ)D�H�Y�mo`���c�-
���~X�Y���{��U��1m�N�	�R�����:��1+#�X�hp� �]��ڑ4����W�;q�|�Sw��"�P�'VMh�(짹�r^3_±�Pq�q�X^=�B[�]����mk�8p�&�}��wma��#�6�źH9o��>���Z�j=z0[bX$Õ��4\],47bS|6���*��ẚ!��]�'J9����pK{n�ԩ��$چ���냈��sK�s-�A���@h,�n�І��ٷ\fnm_Zᬼ�O�z	׮R�a\��j�0�w����C�G^Ԃ�G8�q�l�;��[�7�M}՚���B��G������Y�QGޙ^�!�]�!`�+f6�uJ]Nǵ�7wlM7s^u�Q�J�d��s�h�-�K2򢍾�����̾*�߃��w�q���V[w�"��톷���/\����ìlRw�ݎ�sN���r�d3���{b�^��a��:[�<+b��4*�R�47�%D�ַz�n��v������ɖ��\e�y]hU�E]���t�wk];lY�kn.�_U=��k"�%��ڝ�m(�t��N	�¤�B��[����gsFH^���tS����ȱ l���n�g�z)���ܳB_f}��r�i�3�����332�:Yqg-����uh�j�:V��[Z�O+}YY�S-�z�� �{�-thl'.�j�3d�6���,��p�h�D�ힱ\�~pY�I��������F����m�[�O����lK
]ؖ ��(��%u����d�����"���+iH9���F��pL钬�!u�1��Z��㲄���d�e�|��H�Y��f�4�Wu���} �1%t`����+f�3�Ț�������x�s��*d�Ss�<
�*l��#]9�%D�F���t&�+��ʷP�k0r��a�`��z���ޓK�m�ҍ�d�0؅n�T#��-%|��V��My�0�M��}�f�!w[34̒�Q<Cz��xW(��ɑ^��/W[5�w]�e�"%�7��N
�i%7wX����;��{Ce+[�,:;����'X�n�&�P�����m�wļ�!�3�>��Y�/~�{xN�5��{�8��C��oOUMM��D�d���"r��,�������XV��V��Y�<�����k��}y��Ļ+�m��d� jܭ�pD�YՃ3 �}����%;k5Lm���#jJ����
t�aRǣU��mFv���Q��j���s��,��1��`��jО����RM��M����dNd���v���á�e�wZ+GI$�sN3xSM[��1�mV��.����R�|K�UќպlP����˚BO�p�w���2� �}�U2.��+[vN���1Nƨ4&�����u�E��rxE[���ޮ}u��J�C��3��aS���Wv)#���@��לJ�c�}��Z��{'^���W�����h��r`'"�:�MIc���慅%K�)��p�*5H�j�o;+�@�*�Ѭ�y�������+��v�qc�������Üwz+V#ئr��� z�sޱӧ�����Z)
�����.��-��t�Ew�.$�n`�M�7��������"f��u��٤�o�˖����Z렭��E�pW������1���U�q9�W\C# �^ѡn�Q�u3H ��5���t����i�8u�,�[�	��ғ7�ٜ�\pD__���G�/��<l�L�r�=Un�nG���j��l��6�©N؞҅��͋��o���O��u��T�)�'�7`���J�J�[K������خq�`�D���N`=���ڕ�]����2*ug�4��l	Zt��F^�vYWGS�nv<����KF�<��fH�,��s�lP�7���<��gw����jj[��L`��3�n�pwQ��\�.zwt-���
iU�Ku��j�t�Y�vݦ-J�E�]��I��_2�����<�,K�d�y��<����!�|V#�b�f���^r�E��S$+2�gY�V�XǨ���m1;6KƩN��E��Rܳ-���nҥԘ/�6&+�^��a���*�:]�����l,|��n��V�-ҋz�釤�֘0,J�ͤ6�v�rX��bU�����ox�K`ѬWk��	N1(��x�r�^�xv���y)W��
�h�Wm���S�v�eacAK'�;�:u���"�	#�u��'��s;���O4G�;�3d^�t�D��%���:P�6�f��k-r��8�Ƨt�mE��3��������v��u�ݮ*h��|7t�|I��%k�Ů�&�l���֊'�l���n̍��ukK*a�.��k0��f;��&���r�-X�q�w΅%�;~UD�TZ�);m��������r8���_@{x�5/C8;e�H���(����}��T��,	�݌Yq`�7!�v�����
���Y��vq�b��s��S;�
�+�1���LB�L@�5u�:��z<ȷ�-4�B���^C�Iܰ�XE�m-��E\���V"�e��f@�t{���"
���I�2^�r�}��v��vb�Y�0r���kHg8bY.�'�l-�B�$�y)g,�޵�o$��mq�g+�ņҾd�;@��<#��F+m��gT
���
*��\3��X���K�"e�7K)�J^_V�tk(����T���b�@�KY�nДW��Gt��A�3�[�AùH�3�Q}X4����
� Yf,��nfVWm�:�R�
���}	;_=�5 +U�Z%��_@���#M�4����5�w6-�.P}�x���11C�<���{Y|�U�:��]�m�/i$�;|vJ ��]�8?�_n�����r�ŎO�-��S/#i�,��>u4td*g:�ض}�rVPň8/0T�*�P|l�-�Oq�*l�+��)�G�X�9�%����en�<��
u��_0kl�B2��&���)�������u���m�Ϲ&�܅s�,���������ԤA�СY��r���sQ�!y ��r�3��j7�ve�k�@[�����/9�n��C�������o����B�8�jQ�K�VV��\�)Xj�5�ݐ�fad�P��k.�Uvɚ�vc�8���p.ep�� �} ��M��1mL"���ަ${�-�O��Lĳ���j��[��V�\�.�X��o���1:Z���{(��xCܴJZ�l,+9�t���逃W/���A�_u�i��P�ն��5L����:,���?X����n�`�Y�R���-�k���~y��]��{nw&��ޥЊD�����T����v����OVo!�1rCN���r�������G�mZ@��Fm�ma�Ms�mLZ��|�66�W�|$y��t[2mb���]m!A�\�s��;�V)��j����5#toW�K���~��pᎸ٠;͵9���:�U���}WC���'���]h��p��t��I@!�IQ��:���N�����P(���F9��N��8�i컡�,�:�Z5��>5l�xW��z��.��oo��K�[��:M���
X����ц����^�ּ�o�HB@��$�=��W�U��u�O�W��kHoEE5��7 $S�om�� 9��6�/�V�V��5�V�Tv�=ܶ�y0�gCS��>�<�t���)\�
I���'���81Y:�՛rs|���Ҙ������tG{0�Z�.���v,ճ��լ*%���{v�@�ǵbWB���]��b��Ф�	�#�zY�+	�S�ͮ�q�V����GyR�rYF�!cV�Zx3�����^��[ݍڤ��ʡ�c��j�ua���Y���k��hjMW�Hz�	�f7�O0vv�l+�h��u&�Qێ��YW�%��ou>b]2Pt�wlMy�+�B����*'�Z�����Y7E������=D����y�^:�e�[*.�o�n[���pҒ��-n��V�:f!W��NKG`&���]w�l�㼙}�f>�E'DT��#Yd�?2��WXJ�Bv��vXs'e��u!�7�p:�{3�Z�X��n,�A��}��wz�Bu>9fnt��S�$�D*��Ys��v����1��tuǅ�k�n��r�# ��U����ҵn�j]:��܅���N��P��-�����V!�03�%W�}�sU����UU��6�K�(ޅB�*��K�a�V,nwt͎�8A�	�7�ƪ9�&X��r���5�w�{������+��D���n�j��I��\۰�vv��}����s����ITP��Le����}DETb#*��**��B�PAV�`[�H��֪O�fZ��̥�
��f6㬕X*�rŪ�X*2)q�F�TH��R�4�ED
ʨ(*�U����D�5j�8����L�V"8�KK��+mU�ZEUmcaV�#�5%X���Uj�X��EH��*��T��q����E�+"�kQX��D�Ab�$T`�P���a�aJ�IrX"
�����%j���(�mT
�W(V(̭+-(���(��E����#�Rڱ�W2�b�ETT��X��8ɨ�"�Q$Z�Ҩ��阈�(
,PEi��",QH�+b.YTX�("2 ��dU)Q2�EQQ)�����bfQ`���AIU���A���(���"(�UL���4�Uf%�XŊ��iW)D��[E��,-�ЬV"�*��VՈ�h�X6�� hQ$
��7�<ᙲ�˧Ϧ����\�CqЎ
�.A�(=�/-.�8<�L]��Q�a%�5�H�dL
�Vkpo^ѱ9ڧ�~�Gӎt����+��8hi�����+���Ժ��T,(oL�f�'�r7iWx�B�z�g`�fe�_BrD	�o�W$v��8�>��H�U�!��^�K�I�"��ys�C^���e��E�U}��$�i�v�\+��8l��g�_�tlp\�� E���<;�\c�����M��5�"r��\`�B�rPvc0���DI7l�-�9=���Bͦ�J�C�j8E��F�w4'�T��'��D:ލ���@P�>θ�yŚ{qB��7�@�Q{L
<)�"���Bw�\s>V뚽Wܷ���]�&Vn����`��v|��ο��Pخ�X� ����1:d�b��Ư�i��50u-�ޞY��r�~r^�����CǢX����˞ڡ#b#P���q�%��O�\<�Q�=��]8=��W�!	����*���aB�[0����c���%6�Yj}������s����2� �����?�U&o�^t� ���#J��� ����̨�`�%�5ٛ#��{�� p����|�H^N�ŧ�X}�V�Vt1&Xv1���e�� z�0�^u�u�%�F�5v�
�F��j>� pI���1���V�oq:�/]�@�R��
5P5.�3w��7r�jʠE�q��7nWP�IWk�>���x�/�Og���貺����l]�u9�i3^>Nt�RY0�V_9�]DB�:(o�5\>�w>s d�v��k�
�Nx�)�#���2���
C���b�_,��#U:H�<q$_�c���Ǌ{��n[����2��Ip�w �"3�F�V��G1	���WNUy��6���o1�����O�~�n��}| ��fT��L��72��������l +��V7�H?n�l��vծkwl/��c�[U��;�Rn��@i_]�g�>�y��٪�%������GWz��' �aU�>��%��<��9/n�ұ"ta/N ����؍�Zf��f,z3�����:2K�҃�N��/��)�MQ_v���@��EF�=��Âi��NK:�b�!<�pB{��8��5K+�j~�cۄ �����'�����P#d���TUY��=�};��/�|�㘓g������Ɍ�)��޶ �4�%�]lWc�=���������I�8!��:I�_=��p)1�T���Q���4��s��l=����fkn�;�w5Ԩ�@GJ?gƧݯ�N�k�@7%��`����Eb�Rj�	��֥�ơ��sr5��z�W41v��asT�p�v�#�Π�\��P��K�V^��j(պ��8Pޕ�f�h��g�	<�� Au�4�	��knկtQb��]�`aX�O�<_T�+s=�7/0��Z=�
�Bc]����gވ��+4tzg��K<�$���9y�-.�j{'�3�_e�v���������.?�z �n�;�n�Rq�\�a�t׷+���pu+���moZu0'b���?O@��>�݄̈́{̏�]K����۞��??K�s�œ���J�ɿ��
�]�aKE�zX�p�J���7��!�!��1�
�qa)k��2aq2Ɉ�S e*�n0�+J��
�����8#�X̫���l���i|��w�;]�S�Xq�u,�.�.�B2\�!#��\�/qu�F��?&�
�v2�4fQ\�,���t����8*Z�	�ą�	l�'������(�u�
�8���>����j%8wü�*�u���3#�BuS�c�5H\�L'>DJ���-�g���C�G�fjk�+��
�(?���/�1���;>uJ��@8S���SԞ\�JY<I��D�&h�7xƬ�Ux�R�����M��g/�*���Lc�Qo�w�u���2b��#,�Z���Yhp��j�*i�t����޵��Uk��*�zW4�qU�y�Fܻk����sɤ�>�vfu�� U�v7�f�b'��r���$z㰪�ؽ]��������x���Е7���3}�Md�k���ΒO���� |'���tX���;'�b[/�V)�FD!I��S�{�V�pH�_W��̗�P6h܌w�ʡ��M�qO}��j]���o2�\cwZ	̌Ϋ��[s�,�s$�ި����-�g}�2�e�����C��R�p��<��h7S�V�����Ӗ�j��۶��Z���w��L��~�/���o�-n-�G�u�<�s5��O>�6Ul��eu�o�s�V>�;>sDӛ��N���SՑ8pf��5[���{�ึzA��O�?#iћ6d�p��2%��oDj� 
����ŵ�=����xa
����L�#g��o��T���#�f9�E���E��|�#"-B:�qߡ��2����ܮ�=��uv�g:},�k��r�ѩN._�w���2���<uOL�w���i�뱑܌	��ԙx���	�mp�K��.�cB�W ����O�xT�8��f
��#~W:���[�4��κU�<�>�3�E�\܌y�B�z�*���(N�G�Y��z���U�I�{�W3$��*�C"U����|8g-��;,�KV��(�MXv�|XE2z�>}�x���G�G����n�	���l��/%���c�ʺ!�漣�ʍcz�0���F�"`�팎���ρ����N�P�c�3�Т�p�}9��8q�=#�q�v<�u+�OZF
y���B�yN�
G�!�Y�CԠ��۩����_a�'�9za�,$�_�Ncx�Ok��8�n`\P�Uf�$��}E���Y�g�q�L=����H_Y�p�ԯ{��i�����@Ju9��|��Dr��?y�̆݅^�BP@����UN7lLM.��q�ݿ��!Ɋ��M2:v�t�'�صoo	h
~�U`{�a	� a�7��3�QyDu[��_iZ]]�N���
|�)<�}Д���f�)�n���	9�{,��HC����ʘǩ=����_�ۣ�o.ryL�ܞ
��ϯ��0�zꎛOn᱓8y�T��1�`��|��S�.����Æӫ��5�EZڕK�����^�������my�b�O^F)zl���ub�z��tX�9Pō�à`�5���q�L
��7$\7����`�y_�`�޼6�-�k0s�&���&�yzM���Q�bd��˿8:��^V��\��V��^o��j�����^(sܯ!�W͌�ɳ-�܀#���m��!e�^<`�
��E;.n����f����b�\�2��P>�}y9M��x��&°�ܦ�d�|�kڈ���%��6+���g�� 3�_��w���{�䙮���n�ت�m-7bّ�p�оz�ip��S:<���>p�����8t#,���oa�eS{\���q�E�o,ʚ��Ja��f��5��ӷX�AQ<4�� �g�t�¼��uB2�����'��m�Ubۖ�e2�徨�l�1���*�@�5�:��W�ڲ��Rg=����8$���|�8Cə~i���KG2�7	��q+}�c;BP�)gP����)�<���U���n*����ɱȬ�Y0�֊�7�d��w�)廆"��L�@]�����'�Զ������2��e۲)�L=�$:�l�M��*�ɲ纐"�68r�!�86n&�Ԭz���E����]���g��_���M
+i���w	}y��+ސ��,7�ݔl�K"�s�q���K�tg�mU=�"�=&�e @A�lD��93�S�<=��� A��Ҋ���6����:d0ɾ.ONH��d1 q����F�O��	�ո�]�nk�ֹ���1�x&�Q`�0R�Nt�m��9�N��bz>S,���U��.(Y2��{۽dsv��s-�N�mk�m�Ms�z���mv,[3�$p8/�x����"�S��-��1�f[�݅�\W�`���e;�+���k�;1��6vt�7hC�ƥ���,�aT)��{6�޽�&���*\>�������T*2�*f�/�����^� d�5À��S�;Y�8ҡ��'m�>�r3^�`us�d��X�EDwJ9�X�TB���h[����M|�u3�;�8�ڞ����52D�~�c��+�]-W���u���T %,1�d��q��Ď�U��-����W$eٟ�кN�%���v�a���Y��3����+2�F�Y�9N���YoR�1�KݨX�ă� ,=�٦O	�)Z�r�J���tR�b��R{��ϝL~Jw{F?7�U~s����[�����x�#��"�������N�_c�vM�v[�ᖥL<s�*��:`���eqس�{ˏ����tn�Y�l<[�ҟ '�B�E�b�~��z����Ŭ�Q=QA\��֚����r���1��}e��
��!�ɣj��4�%81��Uh:�&��	b����X��D�1q	�&6%�r2�Z�bOw��i)����i�y4蚬�U���zM��V�p�V������(���(������YR�g3o��y��*"�V�w� ����a��^iA��3{k��۶ٍ���V�1l�D/M!�Ŭw,%��ъ�,�a���Vt
����֞�0,��O�Xo`�ˉ�5˽ON̔S��*)��v����t���vk����U�=W�(Ԋ�u(X^@H]��lx=�����H�C3ҷǹh�z���S,�N
���B۪�
�-��|E#��U�򴩢��c\{����;i"���Ft�Y1�8&N~��Y��_ȇ\A�N�+�ݨ��g�>�gl���_�u�����V�7�vD9�Nb��s3p�GL'w "�D��½��/^l��Ѻr���X�ą����Q�X���Hm���
��[,��@���庡�C}��;F�et��<���e(��-��O,E�.�5�X�V)��SB�u�Y]I� ��u�m�g�
��ܻ,h�G9<b�Cr���{\i=��ʗCK���)����O���!�<�aj�U&��૪#D�wp�ඎ��˙aa���Q��r�s�=�Յr��Ҕ����6�N��?�Ӷ9�(��sMkο�Na�,��A�rP����F��]X�r�u�!��b��-��QcV��"�ͣ�����^�]�+= ]�4,�v6�ٺ�5����+��6�m?;="�3'��גgd�b�uɆ�SE�YB�.9e,�죍�:cY\�Ƿ��������b�\U޵�M�rw�3,�>�p��>�8EǜлI�p�p�8�.�o}��C�~Y1�1�--wCW�U1 _��4bE�rmK��u�z�Hɍ�4�\����ݤ�
E�I���gQB�gy�+:˅��nc�F+ Zd3}_j����t�]Ϭf�Z3r�����R��޹U���`�<qO<��崟�,L�ϫ�"��F;>}L!s�H_�VT��*��⺫��Y���=C)��X���	Xy6{�W&�n�E}�=�mOSg�c���B�L^�UU�!0r@ޗRZT���8�;�3q#�W������+��ѵ	;H�4&q���K���� .*��k�Fv
	�쫝ԁ1�k��F�����s^)a/���x�eӞ�f-�E�a� yVM���odQ��H9"r��wǳ���\$!gC�pJ�q����ʚ_3��Գ����ݑ��V���q۹* :�W��J�q�Q
5�XG���(\�^�\���Ԏ�j�a��d�EǗt�� 5�xl��9"�a��3�y$v���.��24eиK���l6bk]�t+(΃���"a�0�]'�'���1�'n'������/^�֗r^�ҭ�sf�\S%Г�u^$�8�4��X��S4�9\9���Ul��CϠ;u/[g�tQ��n�+�]����s�0vݤ�rK����;��of�&p�r��:�U��D��y�TȠ��ꢃ��2�RÇ!��N��G	!V�'n¼)u-���=͂Pj�-���MS}ۣ��8��],;�<K���U�_�C�ɯ/������:
\���1�r���Y�k�
hM8��U��D�@JV��{Q�.'�7خ��<\G߲��y�佝���-�9P�DYZP��	��U�X	nH�Ki���q�Á5�F�n��yM���9��7��Q^6!ݙ��!Un���@W����JW�Gy���򼱵'rw���*#���ѯ���'���Y�:<���_���7���S�����P�Ŷ�m��Zb�.V��Ѧyq,C�MJ/��+�g� H��C����/�]7w۬�4;�Kq���r��[���n[�aa����Gb��

�cpG`��j�L��T<͎I�/J�|)<��P�Y�q ��Od�a��YU!�5�>yKgC8�qȆ^���[��4���~���9Д���Z�z�˷��_A0�Vy���ȅntP֚����{�]yP>����[��GBC� Ě�\vNZ� �F�ۤ>��}��31ݎ&CӕkO/X䫲d:$l��u����}{��S��s̽�dg�����YEX�h�%�.���f7'"�x]���m����K��V�d��Q0�
r�۳2l@���(�ɹք<��R�0���'__swq:��'�����f�[*�hy{H[�2k�͋qk�@�� �)��aog%�:��n�!tBѨ�wYsl��'l�Ŋ҇�L��ݩ�R�*\;Ee5vU�&�)jY(���1�Ί^o��sy�ڤz�1'^�D��3YL���K9+J���b�)owh�{\���,ؽ{�>�����4�q�����e;��IQ��1Q
���z�My�+bP��H�0����.���i�z��*�Oq���o�h�^��s��,�)Xhu�*��b�Z��f�E]6��}��9ݜR�oe$ڻ���b��n��R�]M�&70Q�R

��7/"�:�؃{�ЙA�;2��M�6���Mn���_D��/.����FI*X��u�A��ټ������s����L�\�]]���ݼN1[M�ݚ���8s�q�rL�H��8�-�E���W�w1�uC"ٕn��F3��Mu����Ҏe�����f�w:��]%�qH�Z��<"�X����m�Z��G.�ܥ�#���R����x��&B�S����+���\�6#iܳ������,�NA�Tc�f���Ù�%�͵��56�iu�U��c�PZ�Y�����S�Ӂ����U�&�6�\��	��7��K-"*64���P�V4�D ��rۻ`<l@�� �7Ol�A"�Ƀ�s��"zA�A��{7v8��Z9AH�7N͍�Fmj
�����fwi�J���W�g^ �fa�lKJ��1V�i`א��g2ƈmeLN�
�93�[�uξOC��˶��W�B%��j��������!�WRÑ�!���&��@�3yq`E�K!7T�r�O��b��:,-	s�\�$�d�eu���VM"��Ǖ����Tl��YcN�iuB�ukk(��|���72Q�g��m#�{jV���3YEdsz�rk|mfn
�:����f �W���rh�2� �Y�%j�=,��RӺ0�.��v wɊǔ�.���f�T�z��HX������h���]���h]Ņ�����!m�씊���;ɥ���vW`𶀮�0vw:�'��Э"n���.����g� ���R�8U��9��7��j��吱v�;���6��\e]`�WP��v�k�[+'Y3*�D���ܥ���Iu�Q�mb�d��^P�̹u��;/!����M@�(u���x��n�:�"[�y�
��<�UaJ�r�1���J��=ɩ�����(4�?>Ck\�d�]�6�g`��r�\�d�ӕ_|�y!Vq5Fw�K����G�-�t����po*n�Nk�����>��k��<EQ��cH��drت+����Db�b�+EH �*�d]RR*���� ��
,����
6ؕ�QTm�Q�UAUAb���,X�ĶTB�QAQ� b)kEX�X�V�4�Q�PTը%)R�eaQU�@De�`����ŕ*���
"1T�*U�I.��k%�)�F*�&�m*�b��Ȳ����EPDQTbH����V���TD�+*UF�A]S���(�XAE*�֬��1TQE:h�EV�����QQH���WIc��"�*�b�H,&��X�)��*(�**h�U�t�H����Y�Q�UD`��U���b��]%VT��*�WZ�"�i*���X ���"�AJ-n�ckEC��B��lE�)7+��b��v�.��@�k�r�e0�Ɏ�q_!��Bˊ2�Å������˲�K:j�:��Qރ�TAj�����ٞ���y�^���6�Y��?F��8�:H*�["$�c<gST4�P�m4�g�4��Z�3�i6�hb��	�C�8��{��A���:7�v��%@�T�{�Gv�6Ɉ^9�����E�\���޽߿=���LT�/�*NЬ��{ֶ��d��|�P㧴�ͧ��q�Rz�EX
M��C�0�����hz�0�<LI�P�m��=g��� �N2����y׋����Q@�E��TM������R����9�Xt�ͻI����x�$�
���|�$�
��U��y�:I�+�;Փ���f��ҿ2Tm�%I�/,��|«a������1�=�};�&$Y>��5�"0}H��F��Z�Y�����}��C���:9OSI8�`oz�w@�b:a���2O��J�ͽ��'O�1d�r�VT�t��t�]����;5{d�iQfv����^{ǳy_���">��?�'�+טO���!����d�Ci+��o'V��Y����I�l�A{�5�����w��ԝ5�P�n���i�&0<��6�C�<C��wr�%/�0x�<�X�lz"#��S���:C����~Yҳĕi�P�J��d���06�Cԗ-C��I�+�N�|ѝ�`bI{��L+Ǵ���o$�OYU'S{�j�D}bP�nũS��?A�].{��W��������
�a�x��z��q3�;׸$I�뻤<OĂ��Ag<�b�=��t��*c�;<�"�hV����<@�8�N��}c�,��B"Fz��Հ����S�u��g�ok�>r�|d��}hY�%I�/^��Rc:V΃�6����1�z��6��z��4�Y�����>��AVu���I=B��
��<t������Y+*v}��ӽ>u���<�o�>�7��c�C����t��%��&�����|ɝ����S{֤�g���G״4����єěB��q1�^d!���;�ïi�Abh����P�"b%w�UP�����W����<V$����ߵ��*��4q�����gL��!�=7�� �0����A��Hvg<�1Y�J����4�$���&w5��Cė-Ld�>B��`O��ߴyֳ:�'-S��JWM.�22�.wlP�%I�Ȯ^=���i��t�REu��Xn䏺��WbU���B��*�l��[���5��:T��t���)U��8M�
Fq���w���8Ȳ����)&lI齮�M�{�"7ZWQ�3���]���}�ڷ���|�=@�]���$��ѶN�tʬ��C
N���q;a����gHm&&�|���5�=C�b�h��N��&���`*� ��䘌	�xw���~u��f�=3d�W���0�$�C�I��M��י�I�>C�� �	�t^��'�'_o!�d��3b���1�!��71���(���/W	�wϫ����Y��H/>�)�>B��i��&3��tugHJ�Y��d��&<a�bx�P�K���v�i�q���ގ�C�1��a��k<d#��O�DP�>�	�zln��a����]�0*�kR;����0}�����|c�i%^왺i ����SI6��Iє1 �=x���%k�f���3���g��ϙ�3t��� ����Xq� �{�>y�}�����޺���=���jϒV߹*i�����N�b]��M�Y���Iַ�1��ea�n�>2�ϙ*M��֬8��

m6����"$|�ЄH�<>��^����9�7{������wx�Y�v�N���4�P���jq�������1��Ag��g=�*bNЩ��;��;I��7�& T�E+
»���i٫���!����P�>���Gׁ�->�7]�{���߲�3vO���=B�d�����@�0�w�p�q;H,�����|���k4��T�!S��`q���6��|�;@�VN��Z�3n�m�I~���DB������܍g�+<�k�w�^E
�]���n�$�n��&���+X|�'����fH����N'N�����:v��)���>�h��7I�L�MRb�O�oξ��� ��+�<���ww�}[�3؆&!��LN�c6�!��;5{C�������n�ă��h|åf�Vuߙ�Hq%~O��a��B��oX=R&ЯF��:���,G�>#��b�}�9���m��j{����T�g>�iI�T��nÉSL=a\gA�M!��0�w��t�Y�>g~u��z�$�3Hz�Cx»aP^3Hzo�;@�T��{>�ұ|n��uB�Ȣ���va����e����0crʳ3v�գ���[%܈��Ҵm���*��=~sS��dyY8՜�#��]ڰ��Jp/^f.�M�`Ν�1�ڙ�뀘���>4;�֯J��e��9Ʈ���Z�rr������w#36?'�%|Ue ��v0�+Ϭ�ּшt��q+{�b,�����Y>f+��$��'�\z`T>a������Af�����'>����~ɥd�*LC��=��ֳ�]�s.���� �0�O~�ol:@�V�4�3�i1�O'�`�g�.���'hv�^'�ߺ�N��%I؜LE�泶j�I�*|��sY��B������Ciu��ߣ¨�WW���%o�}a�xb����4>L���t�'�� Ұ��3�q��'9f��6�3����4CL��N�s��bAT:9�5��@�>�r��Cė��Ĩ|��>g��n^+�s�|����#�D!���V��g]�3�K��g���N�玐�{�&��J��s�:T�B�9q'I����?r��=Ci�:=皟'i�C�u�C�1 �U���j	�}۲Ѝ�6��r�^����gY3�J����X(%I�h�N�1'�~P�+�
Υ�&���|݇{���%@���y��J�+%z;�Chu�'��g�[�������{ >��c}���������|�=�*0�}��bm1 ��i+�7���VNҤ��bA���4>za�J�<��i�v�!���:H*͡ў�wI��_;7��~�|~c�|{}{��=�={���Ë1#<��"öVx������S�N�:V��+��<ԕ:}`T>��&�ɯ��N�f3l�t�t����U����z�3l��w2�C��Ͱ�߽�0G��}�>�@y�?A���6�_n�ߧ}}޸m� �p���N!��~���6����SHJ��+�o�2v�hT<3~�1:V����i������e����=x�;:�c6�R�I�iRq
�5�}�g��~��|��}ɉ>OSxÿ�gL
���18s��g��Ag�i�i����y�'P�=C<9��XTh��;@�T����1'��Y*� WFXm0�+��|g�s��-��tU�uس�5�U�"�E������1���ʓ�z�����&��4��P�z��+���u��Ǵ�M�$9�J�oI7��_p
��%a����� �d���!Ǧ�����W"+۟~QU�)���j���/lY0	�r:�^�k�B��i�\)0c=�f'��d�[��=*��Jf����������.~@�o��=��s(�id���\1��6%-j�Դh�kkD�aW�t��5ͪ�)V*��Z�,�o%�-��ݿ�}U���Ie���{��>goI1�1��U�'�ꆽ��@�)�ӌ��cY6��'Ο����B��s�sS�`):g2���&?0*p�8�O̙�i�|��B��㦾��ߢ��L�R<v{3:�G��|��R
�(��Z&�Ι�J�Y*��c<Oub�H,��N���mCա�
�C�1�d�h|��'f�6�0��3�i�LI�����Gׄ�� �1��@b�k#����W������'=�'hz�����7�� �L�:�08�V|�U��m=La�w�4�Chz��y2��5��>gHz�!�;=��I�T=ODg�f,G�A ?+u��=b<%o�o_oߺᶤ�iY�sShv�<dĞ�sAXV_�:��M�R�W��:��1%C���i�J�*2�'��>N��X
M�}�S�x���(��,�~W�)�C�G���XlU�W?o��w��|��g�>q'�P�<���%g>�E$��'l�� w7��钲���c�:�P��
����D�I�bMP�i���w�HJ�}���">b �B-,ꄱ�ɪW��:rgx�û��s��}��Հ���<t����?=׮�i+�&j�N��g�%����3��x�U����В�f?0/g�s������s�C�� �L�sx&!������V>C�1��N���}��z�R�{�"(} �ى�J�әA|O1'���$�Z�S�(q3��5��p���ɭ�;x��Y�K������I�_��i%O�ty�5���a����W~��>ןs߽�6i4��ă��N!Y�8���Ĕ���<��S��nއ�;�=�@G��2ܐ�O\�{�7+!m��v��T�Q9�d��){�]�����3��< ��~g��}Es�)x����y-d}n���]l��n������Ip��3�Ϊ�O�5~>
쳶=�{TEP��ޅ�gWE*x�/H0Z�2s#ŵ�4�.��s�$N�7��ݐ�.VJȟt�f�t�U�'1�x��mK�9�%[�NP��w���G#:�����%��\�����I���<W��
�r�r�s�U���$���_�|>����5�~o��d�����������CR�	��t��� ���{�+·i,�W�;+c�����j^!�NBx��A���q�r�H��nc�}1������K�P;^� q�|=��H�*y/ �V�7����YU!��;������Q�W������7�t�8�\�eZ���!8Q;F�쁪�]
&�j#2y���W�n�P�i���	�;�ۜ�+�c�F�h��]��2k���$v�j[>��Q=�bԣ��Ȟ���R3*{#!L���Yo�����}���Q,J8*�7 �h�H�WM
���%#�&U�wp�|ʵx��u[���C�HTm���C���� EC̩���]%�E
=gG�%�!����^�1n�Eo_-3���\I�����.�"�⭠:�OnIb�L���-�<�c�8�K�l�p�Hu;Ӌ)���(m�t�6�S70�͞�W@;��T�|d��횎�Q��o� ��z��n�e[����]U�{���w�'�!ʻ܁4��B�AY���Z!J-��=kc�z�p�`��k�&�#��p�v�N�y����t^ד~E�9�����зpb�|n�e-R��l�4�
��8)��Iu��+��l�v�/\t��C� }�����y����ځ��t���ݻ�p;�VQ��$8�� $�E{�<󯾱؍}G��G�䥏�Cp�b�^�3�AN:�������p:Ɔ18_�k�����O���*B���y�pȗi���]fU�_�,W�w���En�:�����2v�9����ww�C`�vW\��[W��q�b6h���k��y+s���WS�q��Sk9���I̘��@����)xH���/{��Ӽ�������y׮��ϥ�|'��I�´��u�F���䝰q�g����i���_ϲO�ۮ�*o
�Zɺ����K#�>X�=��W�J����z:���*��g�jZ9�,.53ݷ�!��	�^֣�}c�\|���iP��\�ͭ��N�d�a�ʨO�*�,dA�cz�ؽcr�N�g���[�lW��l���`8Ƣ��a �\M���Zt}��o�*����'�
_Z��zR�`nK��0O��\ ,�/�	M�F?_�#�݅��>�]��۞Kw\+��'�x������6_���p���w�tbw��:v(���x�f۫�"�(�!�&��%�];Z�b�w<�G�֝��F�1���1��t:��_8�ܻ��N���prN][��#l��,���K�����;��,��P��)�Bη�	$"�-�Y�
��[�q�4��X� ����q�v$ţf���|�}����N�����k�.w�^��s#e�P�+����l�s��~!Ҽt^on����M��D��i\����#��ī���'�`dM6��OG��y��y,ր~�)���g�l�4m��E^Ԁ��	�j$�f��a�#n;
�l^��f�t!Pʔ�[5�Q�i�:/y�)>B�E\����i����r��>-WnU[�??��"����������_y�^��-�MF���L�b�*�D)۰�@8`	�rx�|G[G��k+��1�Y�wz����9��5�����G#k^�0�,�_mD �7^��͙^5�:K�ٔ�p�)�	�i<�p��V���V�͔���1��!��Q8��5oO��Q�q��R���Y���Û����mK6��C/&�m�&�Gk��u���1���Y�=�+�wu+0e��Ș���n��n̕�6fX��.��"��*��1H�1-l.yc�U1 U�O��,�}ϝ�{}fo���{��6�[-���iHp"2����;2�b[<�Z�?�Tf��;�~"���ߙ<l�y,fh7ec=r��
��'<�44f��u!�+;wsq��"񤧱�(OE�:6E�q����/�YĿWe��=����&-��)�П7}m��\�W���C��r�[8%$��Uݭ�.���i���4^��e�������y�y�K�y�^Z>��B��������	ὲW�2�X���)U����^w貶퍧j3�5w��l�n�����/O3Y�S���)u��/�̊� �����9�oj��)1���JiGx_�1@񨄟\8N[1��.!��y#��) :(��f;ٵ�����v?��
����W(4b��P�!®"S��g�:[7��_L<xj��lΝ=��z��_����!n���!��/�3�3��9�N{����b�_m��w^��6z)��=�� +����+��1�n�1CC���1��Pv�Z%d��HpJĔ��㜹V�Ї��U�@'�q#>�b(���i�c++zk�X�[b�Yy��7*2|����=Ŗe�Uƈ}�+G.�eAn���1`�BȺ�"(#^����c�l�`���1�)ў����y�z�2��6�p!/���:<��{�im��>D���-n)B��յ�����Ԟ��F>����s��A���5�(4����0�q������p��"�-�<bU]gc~����d�Bn�K��zV�nP>��������
�{������v-�co�[���s����v�Lg<n*�زK���#����N/�G	�U2��!+7F�����	]k���o�7�+9��ϔi���Y�h�?����꯳�Rg�s��P	���f׆�6,s��1O�|�3q��K��0�L!�7�}ϣ/�O�:Y�����}���G�y5�8e}9P�E���l�)Φ)�g1��I��JY��;i�����3�>#��`7g>�zϺ��-W9�o�(�� Y"'=�7��)*���ɸ�8�v����7A�t�6JrTQ��1]�:N��N����&�%�l��P������ITc-'o�k�bv��Cxߢ�ՃϬ��r�B�t{�vE��8���Gt� u�p�v��!�a3Q:�����\貑h��1}�\�wyz��<%=ot^���|�Z�,5��e�)��m������jh�ϙ��N_���j�irh��i��֊�u.e�@f�o̺&�i.��Ȅ�H��:4_�5I9}jx-�mը+�!���05��Ϗ3_T�*�d%u]F* �>&8;�W��k��+�i�Y��b���V�g!>��{$h�i�9�P1�b3�tТ�����Ң�d��".��eX��k	��X[����I�Gz�]��f�Cf,���'K2�%Թ/�*�eܪ�2����S���m��'��}ɷJ�s����g,��O/g�R�h�aꣻ*8���j}׻��e��^�ݪ�T����� ���{��]���n�O�?D$�ȼ�f,��{�;�Uz����s�h�h�����j���ƺoq*��r��@=�t�����I����b���.J��;�ےk�`37��XFAu�S�W�֟w��_�t�T^���a�q�3�
��@�-T��s?>5�@:k���I�X�t�����rԹ�DO��}�>��+�m��,�W#\0�n.���>���X�mZ�0_	Ww���I�3��+��DQ�OY��iȱ��Q]��j����AQW 7R�R��,�I.y��f�ME�yR*����<�).ӑc��~���+�n>^7����%L�q�l�K�� ��L�n�c�:��~�dW$E��4�'��+\/�ڕ�9=�1x���[[Q�>���ǒ1@�j���{���^[N����N�o7��Ɣ�k9�8�aY�.�Θ��A��w��t�q<��B;���s���.�fM��kVq��X��}=6��H	��B��q9ϫn�,�z���-���}���{o�4"7�	������6�X;c��_A{�f�)�%�X��ͳw��$["ڧ�U�tK0�Y\��E��E��Q�lfS�5[���L-Ȣ�
(�	d��$�t����3�Vh�wL�VS���6km��ې��k2WE/S���۾,V޷���n3t�&"&����P�aܬ�,���*����Ӹ��h�6��t��N�<��З2���͹o�=���`1`p�YS�B��Xݮ�qIe �+2�[x�MĻtI��94��:Q�h"��k�vtH�i�r�ј�2���B�.�h� �br��G���46���gw3�[��R]��З'��7���e���������k�&�읥'yxQ0�ٓw�!�ǜG37��v�.l���^I��[{���UfN���:Ό�U�1�.�|zNЍb��-b=3Ze����;�\9�vc@�ٮ�kQ����ۭ�����ݙ6H�]�F�n��ڝt)$�M�n�6��w@6��;ӝ�d,n�ݚ9�Oc�������Cua��]��U�#;&�ee`�X"N�m�ȨoL���i����S�]#ќ�?*���r�U�TJ����En]SI0���n���2䅌߄[Rn�.��lи��U�q�c�h2fN�v��p��UwP�F�w���9��1��U3�mrU+�=J��_�_n7�H��rζDZ�"j�79���bA}}�uѷR�S��ML�)ĳ42�fRN��nZ��-�F�U�<����	��v3e�&�=ݵ��ikQ��~�ȨVՃGc��B�K�W�n���hݩ��B֪��=,[�[7A|
�e1[�*
�mV�k.���kWB|��7���X[�+n�VK�awǯ���4�w�=V�F���5n9�
�8�4��wQ[Ą�
CC֨�ݜ%�d�y4K��B%�K��$R'� ^yE�����]�nb���U��\P6ڳy2[X�Z#�����Z���i�±`������;����4\{,��1y�O]so\�A�.nEĚ�V
W��ņ2�N�V���Ά���h��SVtMA�tr�qv��UB�^�8��(�b����]}L��V`����o�kY�R��+býՊ^jMv�4JF�`��(&�I��6�wf������ZK��������R�Y�+ڰ��&`[��W��`g-�U�rgv����聻NtR>+P�罟j���u��h���ߊjKm������@��N���I��Nekz1��s1\()��`�Wt�-�r=ݏ��\�wa�&ᩢ��$l:;����S8��j�,lWIEd<��m���.�:�F��45��b�]����y��Ƴ���UJ8�H�j�ּ��M#?b�2�ဲZ|e1iT*A�ʊ�8*�6�J[���w��˖w��w�B7�R:��_q��g_&x��L��b��w_'�/m��k`X,QUE�b���*�
��Q��T���M2-Db�UX�Y4�(���CV�a�X�V1���+4�*Z(��K2�i
��`*�Q�b�U��X�]Z.�,b�"¹�Z"i�P�q�U Pb�KaP�U4�ADuk* �V��b((V�")PFQDE]5�,�PP-�d�:�(�PR)4��X�ME�H
EX����"��%a1���W)QPX�t�DՋR��¡\LV9h�(&R�G)���i�X��c`�AX�ZV����̰�e��(��EXڲTJ+
ʂ�2�@EUT��Z�E
�`�1����F����!P��Zʆ!��}���q�#�c�M��F=.�e㌋�:�YG�N+3���GׯA��f�|�����x�y̳UL���A���� D?�c~nuh�(�yFoh���QҾ��ZJU#���4���b{A��}L�ӑ߆wy$�
=�"�M�����R�Xª�p�pt�ڐ�j	��S e*���O^�U*_��lY�s������V��`n���;q����N���z�3 �R+����Z������]��_yN#��YI�����E�Ds>7n��U�7Hl�@�ŷ�4.�jk��I^��kɉN���;�m&n�qWt�n�h��rt�{�!Éބ;��B�[�3{�t�&ڈ��j���F��=�.8�Cn;#�k�꘼�������
9��Y��ǯ�ݸ�qwVGJ%�C�Oٷ,��;
�b��R�B�m^�^_�r�_*{�uqV�*Ν��\	���k��.�`%8� Yb<}���.FƘ!�V�g�7�*6�:���>��hd3"�j@m�bF�0@�<b���0��4������,�|(�=Nl���}԰�0���Cf�̶2�,�b,bn�@[G���e��
B�E�v��I��*͠�k����R2 k}~U���`�@S-vl,|��sP�D 9���dʲ;&�9�:�"��I�wn��s�^��,wnT��(E���/�:iX�O���h�r��`Y2�	�G;X�_l�om�)�u�^s���9�ne�d�| �6={�i�����_��p��^;����ʣ3��o�A _3�v��e/E_ػ�>���)��5b��X'����^��s��+�L��p�[4����=BWc��tt���/��.pZr�!�Va�G�<��%b'g��J��s����^ �[2�9�=y�t.(�^�^��k���z��,�/%)"2�XHO�fU�[�"���Q@�3��q�P�k��T����ϵ��7"�1�+/���l���ݎ�~�X��w�'�����a�C!-ZK#x�̻���|��/��F;"�1�R�ζ/�1Y9 ��Xy_��ܢ��5��J���e�`��=�\)��$���r�cD1�m�Ӧ7�)�AZ�sU�Y�������ytux@��F:�P����Ԟ6c~\�3��+���PX3�e��G�.F�]8ɤKGL����O3�s���L+z�鯜���н���"��5�U��w�S�k���ᄺ�����BF�������eJ���<eݮn�\��6̹�W֛��"5��{��6�Og��5���y�E�.gH�����)��E`�"�[�s��=C�,z�#֗�=A�l�Zl����5m;�솠��G1ײ�(�}}�]CR��a��f����.o	A�K^4i���xZ���o� W��|NwNٷ��켳�ʕX��'Zx�$o��)��vR@v��T�kCԬ���0�E�gu����I�C-�&��6)����e� F� Ԟ!2D0���ﾠێ<{�tE5J^�E4^ p�x���^rB�{X��I� ~ä�[�м�����,v�la�$!�/+�W8��i���L��/�F/�V7GM�{w%űN����Vƺ�֮T�8 ��1G%�#,���"�0d�@lGq�Z��j]O-�C��ܩ.�[�<��{��#ϖ����~�x�~���Ŵ�����p�v��S�$O��nu���-���w�g2Hk���}6F<��}����:o7�
��\�y�9�1�$��qe4YC��.���}Q̱��7L��1l��CW�9�����W�v�:L�<�:�
�c��=I��ϭK��˷>��60�~8*"6������g�R�{p��2����GOg� H��ܖ��)�1�U͹�\�pH8⩁1k��1�f7<���XXS)�
�ƈ�ً�2_aȎ��U��N�J��F��=���^��� =U��n����f�m��)����ph貟���Է�V6�ބ��}[�ac&Jc�Z�g0�^�}��[�ȋ���|�I��nSU*_��Fam�B�N[ `��C�Y��{���R�g�ǖ��|�U��z����">��7Fo4��8W� K5����N�y<��-���:��zh?���r->̻�o��Q�[��͛3;�eY��1�F����U���S�D�M�~����Й��t���'�ٖ(	k�]sU}��v�q�� Ʉ��0;��䌓�+�����K��>��r�7f�Us]��ꀜE�d1B�:H�r�`"�B����n �^���t܃t@�{kf�v���u�خp&ئwNcF�b�J�>uP�f�A�N�.Uh�D�&S�Ǝ�g������6E�:>?J��2 gt�I����p�|�q������v�3:z�+��A� r:��DW֤�F;ӊq��P΂����nbӟ�<�|6r]o,�&��;'���#�XWb<�R�1�kJLV�r�%�Z�U����T��~M�!�kyD��_.٣Hw�=8��.��`b�"`�=�{��J�v�2k!B��a4��TH�O/�Q]' l�Q@�������d�9�;P���;��M���>��0#�nS��b�%��׻O[x]��R���PQ�ݭ4�=y��Wp����o��&���XB���/ы"�k>X���*k�^wͫ�QWkBc7ֲ1���ji��b%[RM2�e�ɥ:5p�'�ڗT����W�]�n�y����}��͹Hg���[�c𘃇���燁�nc�7���>Ϊ���N�%dt�F*����y��<�|�����	�d�sN�F3p�X��S�N�s��?���R���xSoҙ�W==�s�zC����'g�NyV��8��/����r�V���b:$�d�V5�)<R��������|~��
,��w*�؇�Q+�%�h��B׸�b�ͤ{1,�\�Ľ��OU�����K�Z<~h!�<�V.�R��3�s�J���!�@l�����8�ݼ[>�uzrA7!<}��J�;Q�KVH�����<V����ԵM��7N'�����Ȁ�B�=�k�#u0��/mC4Q��K��`7"����O8�v�}�&���E�/��z�:#�#���֌�86����4j�{���nXϒ� LԘ2��|b�!�n�{�3���WBe�#��'J���Vڋ��E:ZҾ�h�܀�)ɸ�!��A�L����k>>OH����J{���ybJ=�����-���d �;��:���׷�xj֫W����UnQ�]q�צ����4�������z����u˦���=����A@�9�5[��B�i���:��6�:�t���Q�ai3$���}�u�Ÿ��V�9����&pP5Ҫ�Z��%��|>}��yw�y��v҈�?9���K&�F33��X��B��*���ݬ�[�Ql��1��F��=<��n��_��]�70E �����r���2���v�U���X��\��~��K��F%��p���e��q��0�����b��d� ��'�Q(nY���ʨ{w;ʈ���r��g8��C�g�ʄͤ�q��3�I�1'����P��+���=?+�ק�n�㖤�KP~�VXν����o^iA� ��~���j(���q��ޟ��l$&~�;7馣��	���MAX0C�
����7Ӫ�9A�����c<p:�uu�kܹ5�y��^��>~����:c�d�{�\��/&a����;���˜�s�����](�ڱ 8���1(�����#7iHM�ڐ�!�+q-�볳֍M�<����'�G�x/L7O>|���a�T���[l�y::�D���)ٯ�[���裣g�=���m��5�U�Bx�2�]�����;��_�8C^^������֨vET���h޷݌F�f��)��O0l�v*��X�j�$�i�|ޥ�d�;�7�tm�{mH�B��V���@>�y۸�,E�̼������oU���X0k2�yH�]�ݺ�Y]9����y��2,H��O't"�%ڜ����8���Lt't�2�T?� >�탻1�,�5O��&����<��1@�I�CPJr�óv��e�����&�]����^\�4���WJ�T(@��F;�G#�D�$�#I����#���������"��r�+��S��A����S�@�z���P�ia/�u�";��Tü�w��L��]H���������tQBC!���e�B���8L��x'��xߤ:��9��>>���V"����� \�r$
,G��Zz�J�q���گ��Sm��>Y;�2�Qxa��P�rbt7�L�)tu�*� t��C�"(
��\��8�A�m��zH�}u����1�#c���8$C�ܐ#+S�f�TG!���p�H;\s92�Z:�*D��tF���T^W��3;p!�f�;�p�����bm�<8
�/W/vk������6k4}m�+����j����j��1N_?7�0����o	��r�8�uJ�%�^�rb�u�.^Zow��*z�@]`�*����
���x �ꈑ��~]:8��r����L�q���9̐�y�:��Pw����]eK��1�a��]��`ވOi�9�IG�1�=�/3[,���"�۾;��f0���EI���΢5.�R�/�Z"p.n�pH0���o��Ο�J��Yu4��Gef�tZ��ys���L��A�\}}�G��t�[�oNh8+\�~�y����6����_3xmTW��X9u�M��lWu�r"_���2=�V%��j�E�wZ���:d�b���j�S���/ۡ�:!<!�o���^�3����:�/��Q�]���N�`ӷ�Y�;*b7��ȡ��I��F
�s�p8)m��M��@ ��~�W�ea.�,�sA�,,7�r�H�0�N{F5v��at�^3�[�wa}�������yr��R�}k����Psn�6�|��h�;�S}Y:���@��\�֝���l�Qo���7�R�q���~�T%2ta~3�G��Lz�evދ�w{�ͮ���Ï����g/�00�;W_�s�}����|޳N��Y��/���Z1AY����nT<��"�S��� C�F�i	˚���ch�$^G-��Fݻ�z��oHp[�ÐKgw>F�b��.+\�e9��S� ���Z���MD|�ѨxO��p��k ����GҎ�	�����&'����b��"��*���ڂ��`��YGa�'Z75�N�S���f�f��S�C�ou��C/�B9T��V���Q�L��)�F��IT��5�x5�a�{/0����k%�X�C.Սq���}���4벗.d�vAG��6��
a������6����ƭ�5�H���;j>��Ds5�~R������s�ޞ6�]6c��־j~B�W����:�|��5u��+�<Nٟ#X<�:��Q�TE�&�`"c�P}����^>g�cɊIo2v�H~��_��vY5��{�H�!�G���c�Ϊ+�]���������
�U�+w�$��Y�8 ���[�x���0;��5��w�Q���&�B��.��=��'ޙ�ؙī�����-��NDo[ W�i�M�sI��t0���$7�k&��5[&�}D��s�ެ��V������eqc0'H��[=�~C����ٙ:B=�����Zق���G�Ŋ��PU5�\dι���A���I��1�eq0����ekwT�Zk���*������~n��@r|�xp���y^5��-t�PʻJeߜ���{�]i�y˱e��ظ�Gt�ѯ���.>o����A��-mܪB�3�sH�';�Ւ��:����Oj��v���c+�FqO/Wg�n:�A���P�;־�]Et��:�e��Jv�ޗ���heZ��J����K7XRk���8��� {��A�q�9B�ǯ3�:�o1��\)V.�C ��+��"�6��f�wZ⹒�rʻ�?G�N��* ���]�w;��mY����}��^���糋=P��ݎNӇ9��_���J�&��H��'j2��?:��uø��G��9�Ց���C����$L!)����R���ܾ�mUi��+����Q�v����"��vy�����ye��Pub��,W��خJC=@���hxvTT�<���
�f�S:��\�&n�h�R��̇�QHΣQ-���}9z{w�p�ZuS���ib�g��@��W�;C��0�X��S�oX�-�빇�8u��ʐ���
�^%�j38,���x�q��czwc��nA�<��+d�M��\˺�G�3;��pT���H@:f�����zV��kc禞w�q8:�nX�oVv�.Έ٥ֆ��b��FD ��<�c&�k�U�O`������1ħ���J��s�6�t{^?'��әR�iu	�o2���(�����T;h��T�h��\��Ư0�g=���(g�g�DxV[��N��C�e��N�g�V��ϡ9{`L�SX��v�9�zVa���3gF�P`��o�o�ϭ1Z������1ʍR���p�\D`�%����ۃG^��t�\��%3a�"�Ϥt���u�f+�HHk�cO[ZH�%8\�\�eS����)#��8�NO-�A�q�}�4��p請X��.�� �#2��S��/a�$vUjQ"bV�BD�/	�hm�б��ܶގ���a.�v"�e� Ia�{5p��x��9.[K.��]�L�\ĹrX�W%�g��C��#"���;j���w,��Z$�V�wWX	�ޡh/NXQbuȐ��`	��G����e���9[j>F��C1�#F`�{h	(���+�W�ڋR�IY�1"��]��G�٦�-�V�$aŐU�b��;�S�E��q:���ͭo
t�n���4���K�w-��ˤ���֣ZV69�b���j���y�$��;�V���9Ѣ��Ū���W�!��@�5�6�.Ƴ���2��v!��]\b�q�R�ԅ[d;��7
��&\$>�f�9+��#Z�Ф�x�o���w�M*��noxD�7:��[ }�\�a�N��㵹1�x���	�g^�zXf���jhޮ;��T�z��V�Y0sf������$��q��^jJ���sts���Z���?�'���Q�wo^%d��N�[�|��xƭ�Xs���.�V�܎*͙M5��2P�F��~��ԯ9)b��N��N����"��pۉ��-��a�/-����鄍���}ef��su݁.N�[<L�ƍ�c��6��C�i�n���;׵��9e�e˩8�ƴصu�����4`g4�M�M4�)���鋵��,�7���J�@�{.ȊZ��co8jʵ�k ���-�ه��Ek���P�Y�ڕ���43�l^2��Fͻ�J��ݡk����N��C^�j^m.��qL7X*$�8=��QNԳ:��3�j��n�ۃ5���Ll-�;��rRWB�wu��<�� ��H������Tj{��>��펋^���:�j�yˣ����r��&:��宥Mog��M �u�,83����z/t28��=��#�tB�7Y[���p�G�JR[	��VI+vdT��aϢ�&-��B��u2�}
���D7kA��Q�2vqe ^�ʥ�_Ik�3��u�o�J���AJ�*��G�^=��v�4��i�Q#����GY[��\)�ߡ��"��e��_ �Z5�ɠ�sw�iV%[���H���cޢ�-� i"�<�R���xV�ҟE�'b�x���Mn�;`a�u�D-N�jd�ղ�᧩Q�F��b�li�ngS�;]y��3?k�`�}�i�qޣ�����^W.-�U�J�Y�g�������f�M�ov^��ayF�#+��U���-�pnƾ��!����gO���~���3 R墂��ɲ؄���A�$�\s�>��͉^ُ\��x��@t*+A$S���,բ��&%E����J�-YP�D�\eTU��V�Y*V�E�T��D@B��ň�TQ���7)R���t�Z؊��!R��f7*��D�m�bŃ��k5J(DH��*�(eH��VE"�Tb��i�GM�(�b�B��H���%�J���#"��q
�i(��Ĭ4�J�E\E�QE+��(eAI-(�Į5�ˤ�![�D1�iFQk%eh����e�E� �Z4�b*-m��U�Ac��1\�X���X���GX��l+"ȡR�Q���Ƶ1�,R+[
0�+L�E-�ֵm�F�e��U�RU�1��%V��" �-�(��U[hT�X)e��(��k�R���)B�
����u��i��qﱲ�芺�BAhY����h�/Uw8I����[�Ա|���%'ݡR�77�e�g��������Ho&�A�3���g5�:�Y�xi֐.�G�{gʸE��Ɇ4b b�����psJ��u:�K�>t�Q}-���<6�Oo�dC]e��R��ĉ�2�{�F��U!�V�]��9�c)����Pk��kunDS�:�V_��<7 �=PJC�T��ɔ�s���=�;�Q�9Qn�3�����<�ӏ�3�(1R�o�K�T9ֽ����7���=���(��#@qJ����ȫ�1@�I�C_�!������6����r���r�2��64��@��6?F��2�h�i���&�'��]Xk�]�u�8�m��x�7��d�`���3u�eo����Yh�/��G��/�ղ��o�c��������nO���VC��=��Z<�g��a���c=�(�Qt�����й`���s��.�u��'�4��ԉ��ȍJp0Su�5�q��a��V���i�l�k����+V���Ҫ�H�"���q�8n�b918٤[�@GZ��'f���b�W��R_z�9���Us�E���P�=�n�`�*��k�5��ˤ�f_�nJ;��mhu��]z_:���~Շ���,޳�VD�"26v��B�}ԟu����3K�q��vٕ�ʱTնi�L��.u�׸Y[�^޾�+pD�V9Q�Jb�{(_+�U�Z&�XG��J������1�_KX���~������.$�M��ї��ï$��[��Z^�F���]����N͛����3Ys��6;WњI��M߷9�֤��^���1�\��:��S�c���������TKQ%a�MOf3~l�V��
��F3�#�i�\=]�(�AS�R���*
�LT�3+jyw��o�^7�Ӻ�{�po˳m��8������mW��xU�
bu(`����B���Y� E>��*ܑ7���V2}����(.���1��K��Q\/٩��w}�-ۥgd�u:?U�H�[�܋j�E�'������I�M�����}S^4�=^^��H���x���1��ܱȐ���$���s-,E�֥5��4�O�D�N�sП5��O� H�'��(�w	F�	��Rw�����I�e"g�/PJp�F]8�m�7b�eڨ�1���d�<k��(���ro'�P��C����q���~��[����2.�~�|#��X
o��YBP�Fʫ�^GI�D���
�E������Q$�y�m�/)l
��!�[��NVM-�B�����G�E�q�g�˼�L���1��J�˥��0��sx[����]��Y�`��!S�]k����7Q��޸ o�aN��wS�f�~}��|*^�V��G���y-
ͻ��v�q�`؄��;9��5��U	d�}w֡��S6��z_7]���x|	�`ق����T^M�'��C�F%	:sp��n˃P*Wʺ�����!�_��������F�b�m+��uP��j���|�0�T���	+3ep��d�=��=K+���"�0PTx|b%N��$&wN��LW��T1qgrr���b|OY���X{Ϥo%Vzwb&�ES+⇸�.P��F�����طǵ�+�ˢ7c6ϼ���]眫��f��ϗ�f;[^u��V�'l�X=����Ug�xb/���o�K�˄�%��N��<ʜ�5'����st	��y_;��Tk�n$��=��GҺ�"S�׏=��^X�]�
ʽ���� '䥆.9��r gyROu�����ᒒ�9�G��8��63�u�����~�+)\c�G-�3�2��Na�n:���dW)#�V�۽�7975����^� �@ 쵬�Cݹ1�R�=3��>���(�m=�:��o���r f�뱕;�kR��R��/Ku�o-��Zʉ���nWipXfɂ�]��h,�1S�k�bU���n͖x�k���I��X)!�ש]����XjU�"��c�sh�fI����ͦb�8[���!iv��2��1˂g�'NG�}�}�T�=ְ,����vk�2E�t�X!�#�΢vzf6��ꐌQ�_e��x�f�m�] UE30]���o���zb�t�
u�$���9T*
�-r����E^J����z8��B%PB�{/�y���-���5M�tѿ���ol��@���R<ω��=�,.7�+��{|6��y��̬-J���208�/�;;]Xv��c	R �6g����9�n�"f�A�Ӡ*��D�������ςu\=�}�E�߻�k�j�-8�s��� 8��qq���.	���\�!3�����\k�*�����4i��+���_R�pRd-�p�����Q[B� �ɂ����0T�1p!�w�I���R3�2��坢e�R�-�"Íh��U�. �7ˑ�h�J�o����W�Y��}/��[<�hгzy����~q���?Et�!��~Ig� 4'���� /����(��_E�iS�t�V��]Ky���x1��1!��pۈS#$��eH}(H�C5}<��5����&�9�&�L����*t��*��Zp� 4h�)��)z �γ�:U\u.�q����;*Ҧ/�y���}-�[ܕ^һ�N���Ǯjl���~g������(0��ZE4�i$�-��;�q�	]�b9y��a���uv0$�1V�e`�y50+s����5�����+]Cfg��}��UYm��k�!���vMF�o����1��cb�VA�P���'�(ڶk��7��5N[�Ue�a�p)��O<�b�П<���-�TYG>�НUC[���;��ѵ��}ږJ����ˉ��1�u���<;9;�(yL�N���.��7[�P���}���q���h�!�Vb��E�UJ��,�Ži���P?G.����z��a:��2N٠�m{�'nf`�|�����,�}�h�+He�½�W����dׁ�x�����_5]�
�ݖ;#K� ��S~�����#2�g�"2�_�	�W�Ii{��/��ჯ�s$k'�AШ�_е�㑭�!���e��<)�?�Rh.�~N��e׶��z����V��M}%mC����p�Ȕ��e��E�r�
���h��a������lo����q �g@�2J�����VA��'�@N�9�iɼ�M�L�T'6;+׹����A�x=��g�X W��l������A���jWb#_ܴ`T2��,�'D�^ݭ����1�	;	���h�ũ�X�o���9�n0geՈ�w�[E��xy�h1	c��;\�ڬL���w�P�;Z^�љ�f':�uQ���j�}YC���P�=�je�Ն\R8���ҝu�q��Խ�B�:����)I+&1V�ﾏ��î�KV]�.
�.���P�<]�ZA���E�f���<C՜�F�A��:�9���pVI]����"�]`��f-h���?!��Q��~�	�v���O����dd��u+(u�;�3�a�7I���\'z���"�f8@OV}���E� <�O{[�3B��}{h�L1�qơ����MMQPԁ�bxl���,\�����]�W`$@pk���r��#�����U��[����ٴ� Ѳ�Ma�VNLj��w��vu�|��$�,�����D
uE�|��&�%35�wJ7��)��;��>tv�bXK`���Q
�{�Cٕ��HOTL�)|�"S�L`��Y71pc���2�]RG�w������C�m;�=��-7���1G�����-�C,�(X�S�t`�/3�ͼ�
��g�� ����u� ����_�3A��D��J������b��t�z��]y�0���W]�����v�������N�6�wq���+��}¾��z�����Kȭb��Jm��>{f���]�,�}��^ō��?eO^��6�.�|���ెJ.�@�P.ƃ	>���0�eM]����0���sӮƜ�}Fc�\�=BBsqT�N�gFNnGi;��G�|���-�j�8��%bΨΎ�o놯���uj�k.�S��#L0�0���Y�d��gw+W>I�|4z�_��"|4��
g�t�&Q�-l�f�Xy�,,=�2�9l�/�/K�uL����7��Lhlhy�T���x�SY�FU�+�$=��C��釉�
�j9�ֳ�p3k�Ѭ�+�C/MJ�y�@�#iĪ5H�N��
�?g��Z}��E�{�8��	.�h�p�W���w�0���0������D	ri��Ƞ/���.��Yz�hS�|����j^^���r}L�0h�t�E}�t��i�����8����B1l�>5�E�^�ÐJGw!���Ҹ���Bf��h=�'| ���eG؝��c�t��2䪬�b>�. @A�lJ�Ù �wNGM�b~��چ,r�&J�}R���B��ܗ���x� q90���7HEE�!�?gز��'��=�=IvV=K�.���|q/��K[^ʛd��^��4�vڨ;>������@o�S����`�J���;6��S�<�W��i��t-L��Y㘣�C
;}���k��En�Ʊ&B]���T�t�pu�l�m��ʻ9>�&jOMgnZ�����{r�R]#]�#���ݺ}��M�#c���
��6K�*�MP&*#�W��g���������wX����7���ȷ��'ޒ>B��e=5�����C $Xc~�TWI�,��Fؽ�+ߟ�cJ�4����R�}��</�u�i�4�o�նO3�_�%��:x�c�1o��ѥkJ�e�v�iM�M�yG��+����f�E�\�������2��es�Gz�FM��nK4�g ��+����O���uN!�V�o9z�4�噫����%�~���>s��ל��Mɿ|8���k�i�?6^��͹�����Js��G\KO�Z�w�~���}�ڃ1����lʰ�Mv̦�uNr�[�N�)�n��]���'.�s=]��ťZ����z[\��nY��/���R����P��T<�S��xB�*1��v��#�����B�u���MLm_�y���>�T��<4-t��7/Q�x�oл�j�tnE�_;p[��.*蓠���|C�6���Z�b7QQO1����M���yp�a`wW4t���-��w^U�����V�mwì2p���quʳk\b�=2�;�����4I8�yk���c�C�#O�ﾈ�I�;ukE���r���ה�BN�D��}S�y|�:y�Lb(1����ŷST�09���۹W��o�{0�m3+>1�����N�5~�X�;���k����QNf�:����n9;<ƆV�l<������+[������� �z�}"��r�m��N�������h�+[��OHҭ�U����^�.�K��F1��{7��r��#��P���
r�C;a�s|F�yפD��x=��x���o�.�+�i5��rt��_h_ڜwlV�A�SM��,��5K����������||��;���@�������=�����v���s%�N��)�������ˋ�3֌��v��mbڏ���n����p��*�OV�-��|sXN��|�9��+�`T�~�vqKע@�/�UX�V��ڞk�Jpm�+��V�l(��l�����}�]H7Y�0.�0�tgT�s������a�#Ηx*Ӯb����-��y��=���Ъh�k]��Q�¹�U����k31�Z��]������6�oÃ!gm�|�$�`n��|O`����n�m7hQ���7d����DVU0J������
�Z:]�l���Jf�T�}��~u���z^���Fsn>hw^Bxw����Z��E%�9/���O�g�.����	�=�y�Ʒ�yv������'0U`5OR��Jo�߁�}~�����*OU�rXv����Y��W�V����C�bq��j"շ	W�!t�oa.�[Z:�t�֯�^�bZ�Sd{ڼ9�tܸz2a�$Ų�BZ!)㣟Z��E��kK�WJ��I�n��M�I��cۅ	�'�YèrE��_�=/wNޭ��V�-vXK2���Z��l����#���RˉYc|�!j�s���g?��Jܜ��n8��Lm>j�|>�R�N>��N��$��o'6=#�SG��/6�t��8��r͎T2�S�g��ͫ1�ۊ��B�&�t�o#9���t7����Es��w������w���;���u�%}6�u	�9��N��v��}I��bU	��Z��S��)vզ��d*��szjf��]�{,��
6fP����r�֍�R�\Qvu z�i%yܴfM��G++�+��l�����V�=C�$*�ۭ�C3�ʹI��e�I[�*�V`*VD
��lC�E�7�X].ۋ��;Ō�On�m.���b�O�5��>�������8���%���zpY2��[�|K�͛�ēsN_>�y���)��{Cޤ�U��ҭ�=b��hdl=>�ÝZ3eӍK�xw�(��o�0���{o�C��/)�W^�s��l��i9�����R�v��M���OU��u��jFY���n�-��A[��찣n��J�@�}��V
��JG���:��[�(v��Ę�W�O	�.�8�oKw�fc������L�!颒�l1u�*=���RL87�=(x�=l��J�v=jàz��f�q_H��e���ADG��e��m��)u��vx�~:�^��Jpȩ[��\�୾���3���;�����Z���
�������˶���b��\�9�n���nI|*j��e��͗}v��(U%�N1-*��w��xp��<ka�X�I4s�Գ�����V��Ǧ��X�V�D�0̴���d�M��3k������UY�2�r���H��t���E���H6ې�jc}b����޼Y��N� ��E�Y-�-���:�@O�G(�� ;H	��9�L��)����<���4�����Y�����v�>[ge�dvK��emLɡ�`��/���&�C:Ҭ.��`ݿ���^A�k���8�KO���`�d;덺kC�2�EV& 2���l�O�9u�]��o�>\�� ����0S��;[�X��|�7yo$x��G/�Þ�]�p���0f��5:��l`�J�~��S2��]ށFh�L;�B�v"g�u~��6�6���eIjᓸE�ȳ�2��]��d��O�W��]X�pxݙ�sSpm÷ �\��*��z�|��VjQ�2�c�tG����(�����U-�n�W62�ŉ��Yr�fjL��N�;S��v����Պ����5�/�IH���J����,B�A�ng��)Cܮ��;���e�^Z�bɜP静t����զ�P�qAk1%.�rx^�/�uJ3Dl��z���bm�חy��
��{��nSj�p��|L����9�1ҏ����d{���k:�r�b뉇��S;F7��bR:PΙY{�I,�lN�8�nJ�a�;� �n�2{-���e]u�&h�L茏4��z)��;N�0��X��R4:�V�x����z��P�{cuM��.hC*ߛ��Ug��puf�C(�Y���˔�U��X�r�@��+*>��� ��C������7E���^����a��QSQ��#�k�7i7��U�#ÌM,��;+��}�u�;ff9 �%{�,r�)JZ�D
ʫl�Z�m�j,+�LqD����+�kA�YJ�TR�e�U*[b�
��ŵ�tɋ���-E��lX�2c���j�T�TZ�ZʑV�+�r*���F(�(]fH�[R��++�`Ҷ��*)R�PQ���cP�*�Dm�j�T������E+X�+R�Q--B��j5�֖��B�V�c6Ő�EK�����dQ��r�
ֲ�ڍh�+Y*V�e� �������A����Ab:jb4�QQ�"���P��ֹ���*��j"ĥ
�FF�R�Y+�F��%X�eb��R����J���J[QE
�
��hb\�T*�Kb�J�AV%�Am�k
Z[TV�D
£[m�5AhIRQ$�vs�[;\�c;ך�[�,��Kn��oL�9v\�������/���]�������x.-���ﾨ��t�Ӟz����R[���s�W�ο\7Р��R�Yf+��v���]ܶr����z:#�S)x��� ���:-�j����a崶��u��m���q��b�6.��jy=~�0�rKjKO-��{4l/�T��Q�6���|�q�<Z�����^��)�ŹO��I�G�b�cM��Շ�hnD�1}J�=�o���X���<��Qްݭ��G�Ѓ{�s���������c�������`�s�_��y}�5��_��zQ�oɊ;䧋h�nN�ꋦ��ǟ�xw�?U���\�T#&�����Q���j�5��лn{E[u}0��B��doT��40� �N���z<Ư���5M̮>y_9M&��Q�u����}�-�0�Ƹ����( ׳ٕm����+�q��/��=�!����)� �²	��ʺ���MG�{;�q�3Ms��U;A�֧�h�0�+grށ��	�Ŗ�f`��(�c=Hl�Av��^n\�pSM��f��xL�'rv�r�=pv}g�J�u��I4|򻻦
z��'k�T!�4�>���G�⬑�J�u8�[Srŵ�|>k�v�q�zq���C��Et�Z��.��)�|��=N���9Y�ݳ;$�� �T�|���sk}VI�4�EoW�����[�q<�ⲾI����ʿ���m�.��O�k6�#��2!1�I�\+{g���*Ǟ�t�@PKη[�w�co�ت}�u���s����}�f4�=sY75v3�#ʘ��Q��ZԪ#�\�*M@ڎyN��'�c��
܎}B�A��Y��o&�N�w=Q�m��������:�|�sF����j�n������U�Tțpo��8�֪������s���6/��p���	t{4D믷��9�ZVaq��*#�fQv�+��s����Q���hC�}��ѳN��\���%w5�v�v��Έ�������]�D/h]S�Y^���#�[�^���S�o1Q���Y��͏Gsh��hq�:��w�δ`�cv��5Kz��ņ�+vW_��1�}�n[�F�KE����2�*���ʷ�q��aZ��LJ�2س�\mV�V՘r��n��9���
V�V���UG/l�(ӼLcw`�t
R�}�:��}�v����e�j;rnq����9��o)>X�^��W����1�M5���М���~��B_�5\o������XI_)�w�_'P����;�\=�����3�@�����xg1J�o�ũ�zG dh��ˈN:�~��u4>���}So7_m�-�0�q����L�����e�C��BEZ$>"GO#���M	��y�"ι�Z�����κ�o�}Z�E���e	:�/��<�j=��h�<���5�z�c�}�R�u+��߽�,{p����1������N��������f�_:�f�=<T?{����C8��9P�������� ��/;�'�������{�5Hفer��9}�}iVøbb9
��Σ�l¶��(��4�}y��-�ǎj�>JK�o�9�}p�)��B"Y��N��[��:�WH����ܣMU�*�ǵ����N����2����tpSj�Y�n�5Q@+�V�vK�sV&'\!Jz�f��z���X{a��4�1=�MX�L�=�V�>�6�hѣ�>
u�z�x�o
�6�H�"t�Q\ɼ��ճ�v���;�vE���r:,�9��;�yj;u7��=��+��_iq���XU xz>��F�8��C"}�t�[Vw��w#��+^�/m�J��)��q4�>����w�>��n�����{�]�ō�y�=mmE�qӊ�ν�{���tط]�5����m���y٪�'�?(5rm��C�q�xM1�5ki"�;s��ުk�������bvxOGc��������=�-1�'��a�=��N��<uz�~���-w�ֶ�kr)�
���[ӑn�,�[G���襙�S��@@]�c�;>��Ʒ��&ҩ�Fb�rD��K��.�v
�{c��������Q}'���Ք;T����k:�� �mj���+�	O�cx�q.i�4F����|V�7�w�n(�K�\��ӂ�W�i�7�'�`yz��sl"��{�T�(K�h����]Lwu�bj�%5w�<��`�z�U�r���@h�=lZ-^�2xQ��.��K*P�L��l�{b���q��P@l�:d�ME���K��ғK�M���QpU�WbU��_�.g)E;� l��{m6ݻץ�FB1��!yFNr�۶�
�N1�]m�ӏ�.&d����#Z*To�>�n���Zю�}�K�y�e��6��s��8¸nû1q�͵�Hu�m��DH�'�Ш�9�K�٨Vrc7������}S���s&U�Gf����i=N���\��{~Ҿ����@9u��$��P�~��]پ���͏M]j�uG�)�N�)�7e��+���T�l��f��k֜�Cz��&2��=-N9�⳿>�v�t[At��	.��(H(�<u�_22q.�T�P/�TWʛ��9�ds����Y���e}�nTِ�S��u]�tu�V�M�q{�Qy9_v�ל�Sa�Z5�/��[�5:����{�]���^�٣�Bk�����PqF%�s��)�:{�b����iZ��9�p??��]��/�;�
cO<��Vqѷ�Ϊ˄�#�������(�\�u�i��i�N\��jܡ���k�,�v���۷�1���ځ��X\�pa9���l�̓zz��{�V�����s���Ԧ �,���Ń�E�{��<��u�X�Ju�ˢ�E�w�\5��a�]�C�Z�m�Jp R�`�\�F;7a�U��]���`���9���]q���$7��j��T��疹��>o� ��]�vU�T�3�V9�7��]��c;���ó���9ԛ�p9�z�Boh�n��[�A�W}k��9�I=���-��ĝ��D������t�{4�J���ָ�-8�T�(�Yb�։��oy�l��.��ل���wڡV��O���
���rS����=�SZ��*Z��L<�]K%<w�ٜ݅�JiΧvwr�ر$%�*WUߗ!��=v{0ʹS��+qѮ�����.����OX��m�]vo�y��m5r'����57���xp{-���v���r���^"y����iܮt2�&*�P��S�w[:9��߰�#zxg�xroϚ��^�8��N�+.��8��j!)hQ�+�|Y�d�z�+ɘJn�:�7Qy���-BJ��B���f�';ڔ���ӊxeq���p,T��G�f��"����zRn�q΢3�u��ƏXÙp�Qh�ɯB�="f�_+��&�%�� �s�8�łb�"�S[R�.t#��y�I�f�8%�LZ�<�c��P4���6X���T"�dk8b��ε���o�Z�d�>�6�=º�ݕ��ד�u><�Sbӝ�J'+S��nbf��ce�v^���l�r������.$(Ϧ��>��Ⱥ8��w�ʟ�|��֗�9�����X̨*��O;8�"�6�J�������sQ�,�J�#i��^�lV��/t?{3��7%��U�X�V�
��&�+����g\�[gS�����Ls�Ӷ�૯>oC�ƫ�tNT^V%����	P�V�__%P���)����|����,��\J�����y����3�JY�j*�R�Q|�\-?+z���V�>�O�g�!���f+Q��{�w��
��N�#��v?v�����~�+
Ҕ���;�"���;E׳�w��e:ȑ[K�y��3�D|e�z*7��R�ڮw;�7��B�N���	�^�#@�)�G�~V�k7��#^�M�̫~�5�JWQ��^uKC�OԖp�$.�.W�Ӻ:׳#-�v֛˪5�g1��q�8@O��o�1`֒��ϻÎ�����l���}ǉ�5e�٥�o
_oX��ĤN䧧��upf�^9��2�U��\�V`�v��-�sٷ��KҜ��r�����_ѥ=�Mc;/al�9	ݨLp{:�YY���-�����庣��|����VW*���ʇ��P͐���'sז��j��m, �u�A�����;��.{Qج;d$�6�N���!�[����,�vE��ã��=��h�4�X�E���x�x�'|o�q{�\ҤCx]��tl���������-eA�u��@�+�A}�W��nگcY.ˌK�6�Il��o.��L�0��AmO[[C�m�h�=j<~m����Lyy;s��-�ꍯ���`��j5��Xv��`T�^�%,i���&N��t�?[�0�W�b\�:16*-�۝ky�^���9p��%�ޞ2�z�7�_gL�7�B�zS#]e��=3��r��SA��u��6��Fs��>�;@�f��������a>j��J�1�nX��*Ap0e/L���/m����Y�nZ��ZM%�J#5�������L�J	���C��N��'�P�{v�EK#�CbWO��oX�w�/��⥋,/��4����;O3s�L2�'����
b.�+茾N_��\���9�1�����op�jw�Vڃ�c^}*JL_$�N����$�fSܷ�:�^b�pw����v�I�q���J67�%�%�ҭfLQk_��=m��}�Q}�|�HҸ�ù\=.�+��e\Kj%�gx��ގIYac���U9	�|��zÄ�ݙ랕N�v�s���
.��+:��ݜ%���.8��[�9�lZ�GK�
J5cL�穳i��H���~�;���T���j南NK;��'��ȚgnGp'��	[V:]��X棹mD�Z��	�̍<�5�IR	��U�>�9N��d-��{<��K�u/��#�����]��Np/7y5T�����>�w��[vW���pdF�z��zz�k�ʩ�9Qy�F≄��f֎�8�Bxr���E
�_R����M�b���U��W
S�%i�3R�;���%R�tczr����̬�՜̞�
v�֗��2�M���tt�r�0�p�|:�ˑiy�g%�e8U����k��*����E�3.]��*ھ=�=J�Źg������?W�U�s�J?y�C.�z/w��s��;���m�OKq��A��kN.�]>���	�TAW�r�b�����1\.u��
ݽ�jL��Kx���{������H�i7����}+>̒�-򣪰9��R3���,��%��\����r����5nB/�u�ޗ��R�lt�J����6oLj�m3��1+��]��T}�k��� ��ג�3�[�ӭ]�/��s6���s�v��ڗП:�.��ɜ赍�)B��"J�f�UQ���4�7����F���Yp�t·�M4��x-'M���Y="�v*�{�:��w�N�S�O�0T~��`k�6K�6��Sk^֕8��t{l��gH]^Z����CӬ���N�eG���X��]dAannn�ؕb��-��9�ߡީ�{��n�1D�����-�S�D�g�j���8^������GulԎ&�{ϳ6�NdveInn�4x-���k�� y�;���[,�Ы�Mq=Ӵ�[e�b��篳��l0U]+e=9��/6&,j[Ѝ�ThPP�RYwy�>���C�Ql�D:n��=�1a��ڹFؗٮ�ͭzU�آs�m�'�����EvN�P���w2�+�Uܞ��ns�$��>�s9��L��&;����L��u-ޞt`x%nM�H�X�wx,p:7J���b��rǜ���90k�st��PY��+���Wo!3�v�)M��*��d�a�v&�_R���4�ˎ��U�ٗ
�ιX:ޒ��蛱���jH��պ ��O���^c��%Z�\䷨7dv��oq��D*�����3K�&z�1��W���	�#���~ή�UaY������|�r�����%:{��7Ɛף�k�"P�얚�÷��3N��M�ڸɺ�H%�QJ�/�E:�lI=88���1��b.��[V�gE��,ɷ�1i䑽J6�Y��t�8����'�P�9vIF��Kгz�۳��C5m��!X�.4)�q�Z�@�s��e�1ѼV��|�XlqX9U�Vv�5b9���S�x�t蜬�N����G첃��Ͷ���J��rΥm>QϏ 00&pl�t�ǖ ��J)��]��
�@� �<<2����ڭ8yT"M�+��;s���;k�-��O�a.5�5�G@�`V�P倃��8��N_RZX��,e����V��\�)v�b�g6�de��J�]f����}W,ӌf�E˶@�vL�fq���1��-W��ܖ����f�:l���om7�a��FK����U��ܗM�Y/�Xœ�h"/�u�fn
���mE�%0:!:�1��#��hm ��p�h�0D��w��DR��2���a�kPT���doZ�b/z��m�f�L[��VA�oS2:�L%�������ѥڍ�����p��������J�Z��(,,=�����X��j�+�H�W�TlXx�X��.���E�f] ����Ujx-�T��9swsy �Gt��Ч��kL4��vNqL'�퇓��x�9n�-S�Jq54�Wxq����r�Aͤ�7z���z�����]���:hk�<s�u����0Xh۩+�{��z�e*����s޾�FD�s/r����a*x2]C��X����-#_O������{il�A)�N�u�)��5��.G˄2i�����8kYɍz�xd��;D���F&SNq�����ӤģF�2���E���D����#��ciWc���5�r�c#���&v�������_ٙ)9>=E�4,�	� Ge����*�9�s��J��2��e�fD�wB�K~�u��c/fR}F�`M7ic�2�c��`x�e��[Mݚ/vd
�U������¾%l�"��b��� uC��q�V�p�z�	]�V�Դg|�+�:M���ֽ���v%)%[`6Ķ(�aG�T0@����V)[lR���V*��cb�ҕ�Ue-��eT-mb�.3(b[U���*�KiX"�h�[E�F[p���P[i��l���Ս�kQD*�e�Z�Ƃ�*���K
²��*E�5�m+-�Z6�P��[TKdF�(d�+(ƴ��Q��������E�b������-�AjA�,�h�T�����X#-�i+DYZµXTR�R�Q��"�J���Fe�֠,YUXV�R�3�l�"
mAE�ڍj�R�Z��Q*�UE��TR�������a����U�-�aD�ȶ�U�%eFՋ����V��5+R�T��
DT�F4�E�l�(6թJ5�J��E+_����$>R[����:]b��(qC[O�,e��P�/�[b���3|��o~���h��[�kt�aʼjjg�y�{#�=w�bwg��_Mz�Nh�n���]]a�3�'�@�{M)�t����s��a1�q E�.�C2�j�E֭�EeG*��&��6�+b9����8��=^�.D5o�"x�I��]��ϱ�=��r����5�K�G��xZ���8��1�Oi��Pُ�R�^Fט=��)Sz�z;\hO��]N���,�F�۝|:OL�Qj���w�趂�ώ�OJ��j��K�Y���U�:��}�6�/R�S�[P�[C����qG���F�����&��` �u9�;1�=�L�R�׿9�M�P/��2�{����ړ��a�p����u>����~#UbM���ϩf�x��}���wCN�⻦��7s�*��S����}�j�kr5��S�U���S�u{�6]vM�m,T� S�-'b��LT_%K);��;�kyoB����fn�{su%ɣ���%��z'O�R�Z3k��i���Ը*א��)L��NL�orh��\]���ƒ��������9����K��3�(�[ӁТW��%���7���(���e¯�.o��`��q�q/���["I-Bt����|��{[��b����L=��9��F��"R�_fs[����iC�Gv:�Y6��=���i�n�Dt�_q���Z6,�K���\�r����~�T���1�
w��Ss�Y�Q@'���BN�D�[J��K�u��jqj��'8ڤ�sw��W�S��4,���:WÊf�ֲw*̾��{�Sz�V�-vF���9�$ֳ�������x�޹i�2�s����O�n�o��K΢��cg�����nev9�U�P�.�B���c싳r�����h�,�pB`��^��m�3��.{_r��9�Z�U�UO�oT�ܠ���C:&�v-f�������R�W�},j�
��h��Yʕ�w����n�ӻA�Ȅ��R� +_��,��q�_�����g��k<�ˬ�99͚<ܬ��}�����C-��xr��ܨ/��+3�!%.�	�*�u)R
��V���owZ�Ñ�u��旨�4���ܥf�)\$+]ѧ�A��.�<O��EO`���Y�沓��*ƺj�Y�#�wbgu�X�uΔ�
��ހ���k6P[1���^�*���F�L��C%Ge�
9�w�f��z#r���X[�Y�P�Js�P�.��}UK3����O=���.�)y��Q�z�������L���)o*���p�����ZW���ywq������q�+\�ob��}��i<��*�6��u"�'�M.�0[�V��6���Yg��+���W��e[��\�3R�-W���I�֡�ļ�}���%EεQ|�B�N�|�*%�l���ǎJh����3�-�܏��K��!��	��z���X�#����~E���2N�Ks�]���m\�yn>�z���n��J�%027�\�M��.��#4�{����N.��֎�}�I4���OE�J��U�KEE]�F�5�΁Y���Y|�f;s���w����MC��O���m����4ҷ~㘻I���I�������a]��9����K�q�m�畝�R�x�1�j�����<(���9~��j����so�=[}�͢�e��`���D8��SUL4|�ޜ#�O�憝�xnF�P[{���7��.���N݃�u�K��
��bk�њvS�0LM��W���aHM/�
��6�n�Չ*5�M�Mo+p-���ཤ��ԥ�;j�/;J{�'�����mlm���}�a���a\;���^�A���^���c9��8����I���k�T���������ة�8G!�>���ŵ��/�mot� ^]=�Ϝw"��0W6�R|�*�K�}\oU?\::#j�]9��7;���k�aX�s��E�`�n(�k��ڱԛOF]���2��v���Wu�]D������-j����Q���q1��ݭ�4�b�U��V�~����ԫ�e��X��Tm(��j�F*�ζ�;�W&X�gq=�Hj�wr�s��m=���n�A�o�M|����o���p)��Jp��ՉJ�p�=�ƚܧ�Mg3^��*������>��"�Z�<��n���o)>X�.ͩO����Z֛N�;��u:�@;�-�ox������6���q�_'K(���8毞��i�����8��2h��>�g���m�K-�@0f�׌b����޷��nR��EXL����(��f�w�\�7W����#�� ��F����`v`�(�˔Y{6��ڮ�Ia�$k���B�,d�	�E�����H:h5�m<"wWd:v��ͷ���g�|�YkmrQ��c8��U�YkGJ���
}���o�^��<����s��vI�^!����ɩ�O�0T~����ڮ�It,��m˸u{���N��קW<Qo���`���$�-�*w�>�)��u�d	�;UՊo��ʗ��jY�9�\7
a���<P��ޣ	������s]��e�}�Z�zVRlmC}N��������LpxJ��8�&�i�o��������iY���
���RO	��8s�ap�Cn�>0AWs{����bY�7Y���[Ӌ��N�Pu�B����yO)����"k�����IM����+�U�*���f���E+o��!0�o)ňWD��v-�����y������߂�|�H2>���E�%�<�=�����9��E�r��^,l��6����������.<�Ќu��0ܭ���f����
���3IF�ܩu"��ː���{2Å��g��͝�:��;����X�H}��J�d��m�b�w6�Yorŕ]��ެ���i����ƽ�.-��b�M\��5V�;jte_
׉G� �vA:��y,�!t�ԕ�	�^�]�U�����f'���Ǉj:�eP�ok'�M�{�T�4���/���#��s���u��b�{��jŷ�u}v;�h++*q�l`�t�r��=Ug���puR�j�2�}0Wve}׮pA�0n��#���x"�6�
�걺�̔�z����л`�	��f�����ĵ#�lݾ�af�S#c]D���¯�#\�eq�����{���z̯+��c���4�r+V�U�
���̹�9����_1��sA�Gȉ�>�p9���wL��Z��\B�e�m�$B�)��vv�3S�ā�WS�w�ku�u>�sGZcUC�3�)G�]�Ri��`������in������.̿�,�ɾ�*��&Y��O	y�b�wa�:��E��ڬ�d৵�j�?J���m������z��0y�ʽ[d���;�@������[��հ��A��wgtn�\f�h�^P���Q��hD�����^�=�V�y.��#�>��i�H�7���ՀM��t���i +��ǋ�޽��[+ kg,bTޠ^-�H1k�h��淃��ԁ�p\�cWX��d@P��U��v�w#}�eO|����P���JSh����ٿt�ڝ�{��nh�{�"����n��5�z�J]`O1�En	�Wkb��R},eL�t�����4��D�ɓ���k�더��䯾-ewQ~��T��n�>�%���N�|s��M�����q؅��̢�;TLVK����k��v�M�<�U}9��Gk���د��w�)�(5rPMj||+�b~^w���{4zc+������ֱ�1�x�\ب�o.�][�_k*�պ���ƶl8�@K��ۊ~�����/��aW?st��|f^ٙ��r��[ֻ���3���ފu;�
zX�%��񓷭]Bi.ǩd�t�H�o'�����e'&��`��J��eEĤ��*��<��!'+35]rJ�q��G�7��sI�{��մ]�q�V!)���&�T�$o��t���j�v_eB��]�!+!�f�R�����#���
d3%��X9�*�u�E^2���չHM@*�~<w1�muq�����ȝ�u�ɵ�;��n����L�&�d�̴�z�UC"T��K�)��ҫ6�tG-�]��n�;Gs��pI�m�����)1L򝽍�1�fn�Gy���W�'���s힖=�+������=��k�m�H"����^��V��d>�M��C��t�{4T{��O`��_9�{�C�g35S�G]ue�$���6=�wP���ρ��!N�l�v�&'��u�jާ�kZ��	�,�W�*=��WZ��B��Ъ��Y}�X�O�\j^WLS��+I�!���7{L�jF�djK�ѥƤ�h8�W��E�~��,�D_i��ZGw�_'vQ�N���`��:�*t/�l�]��oZ9G�������xn�0z�D�M�skG8�mQ�۹���gt��}���ʴ�6�p�<אq�G��TGf��}z�b����rhl*1�:�Sk��5n7-��խ�KG���_]�|�B�\z{[`n�(�Mc.�5<�� ��=s1��]�5؇#����bGΐ��I1���ZJ6�os��)�ب���V��\j�VP e6��77= ]*�]��혒(�{Ӯ���M��j�<�[��ot����V;��+��A��p
x��j'#�~���l��1j�~&��j�'������kQ�{���%m�]���1l������j���~�; ��o��1�XP5
TӵN�\�Y}�i;��p1���Qo�4N\�F��	�d��4{��}�[���q<���eQ�5W�ˇ�5��8
a�Za�tŹ盄l�������%L�K�_5�GO���4�|;qk9�P{����h�*�R�%ۯL���L�"���M!O�3�ٟl}3xH��K��v�#M�����%~uQO��N�$V�;ٕ��7���D�;��z�O��SJu;��q	�*�y�&)!�	�Wp�"0��Z��;��*�ݘùI�_4�ͽ����!T> �cD���::�ھ��3U�%&�l�v���Ǽ�G*_$�T&��W�:4ޖ�_x�l��MR�vF���C���@f�ٗzބ�����l[�n�Y��[���z��+'\��Dۜ���p|Տw:�ҽc /��J&��wvF�'G��m�3dН��j�X��oʧ�HK��]/�sGQ��AS�b鼲<C�)�1|�/�>�w.;�%i{��f�r�7.���1�s*��Ǽ�7y���q[6��;J��F�4���
�N�]Ʊ��N��צ��jթ�R���=��,<Q����@�^�\�n��uy���JyS�F׹Z~����h\O�O�ű���tĞt�3�����GN��W���~����|��Gim>߂�G:�ï��U������9��O���׳ޫ g�6��l�iy6�T8�'>gWik͸���uQ�fI���문�͊��\k����[��7�鐷�wq�'���'`֧Vq;���puR��e��ܦ���1O_I��Β��G��Me�"w��I%�]�'Ά��G~[��t�~����)����ɮ��B��N��ώ���{<;�')g��[�e�s=6�75�����p�d�t���_%�6��s0��g^f��7@�EA�7W*ޣ���pp�^^�����L��֭a%��8XJ������?lt�7ҽ[��AY�vE��ԭ�[�U��N�g=���F��u�������bQߙ�3][d���NQ%�l���υ���0��ϝ�̡W��a��ݛr\�5l�ګ���j���r��7*iP�T�Gz^�� ��^h`�#R+igg7f���(qK��K�
��7etw ��+VNsSt���H*a(~�?hW�R}bfIwS�!�Zu�A��b�Xf`t$0n�D��j[\so��g�n��J�0�E�\����b)Ҿ��R�V͂V\�:��H*���]�kA��Aͽ}w]#�[FS*�nM��nz|�C�����\+i�i�@�zc��-��*z�]n!�B�f8�Q03��rnGK%�2fN�`���tS�mw�&�>S��*hL�6�5G�n�rS8���[�ץ�ps����[0����+�e�ü[�
?I�QS,�7��c�零�5P�2x77a]�n�[�h���Ũ3b�!P,�}ko���c�s���s-�剶TcᱮW��K�������]]��om5�]����/�]��sV��9"�1�Ш���Ĝ�R�v�қ̻0Dc�m�}11�o���h��*��p;���+f��#
��}V�/��L�6���Б��$gJ̽�&��A�;f͚�Jޅ�Mۨ�� �((u �##|�*�W�N-��[d��u�
���9���'	��_Jv(T�X��I�	��X'�֬
�7m�r 뫥�u'F6�V� ۬��t�$���9�a���@�&%t�W�n��u�%��2�ܩ6Ƃ;.p�(�������WM���pዟ�~��yƎ<C�Rph��;�d�l�<pM@^*�ؖ�-OC�F��h�]��Z��]w�����n�ȓ��^#� ��]e�h��y�,4#��7C�y˯����+�7��􇑜���K�L���l�4�7;�=���67a}�8��Bn#Q���7���h��ۄ-���֝�EXD����y�$��f>�F`.��&��Pa�9�ANwѡ�2򢃛G5K�|;d�V�gm����<�ѵ��1o}`v	7R"�C��8�/�2s�Z�T��[���˛��s��Q�oF�H��d^.����b�VSɝ	�Мs"�+E< �\�p \�z�a�|^�����C3(�Ù�m+�7�F�]R�@���0�qv�N�)���vu^�/�06h��Ϛ��s&�E�E��Er_�1vm$K3JN���{Z���v]�DRl�ʹ��^N�j��O+%E���Wo�m)4�,�n=���:����"�Ԥ_q����ݜ*����ZI���zA��o���+�Fp�͸�=Ab5�A���B:�I7i颲�"	=��Z8���U��yoԹ�X�&��{b�:Ա����ȫ����b9ôo>�/w��f�Ƣ��lJҴb���Ҫ2�Z�
�Q�X��jR��Um
¤Kd1*,�9�-����)j±�EY*X#�%e�m�FV���e��A�lrјтʪ������FVZ6��h-Ub�TUkkX�"[F+
ؖ�j(TjX��"[-�e�����D����JZ���([-`��J�%-��h�
�3.1���*�Ym����mIR-b�DJт6��QeZѢUV�kl��ƶ�E�+h��b�DF�-m�R"ʖ��P��kj�Q�,�[KlZ��*�-JZ����q��U��eK"6���KJ�K[*R,mm��-A�J��2���[l*�FR�����X���e�V�*TZ,V�[#Fʂ,Q�DQA�ZQ�[Z��aQkFҍVQ���DUbT�TR�b���m���-Ap�9��C���\[�JqΫA)K6x��!�b���*�F�67(wJ���s��ۻʙ��Ӻ��K��ڬk�r)�V�f፾��8�lJ�������`��M'.W�f�K;8�nR�8^-�Ao%;0�)�K.�[��%5u;g4u�cUC�4�<5ӫ�T�7������N}j���w�|U�$nvT$��s�o�k�*9���8�7v��l�ٮ/�����Kj-��&�=ێ+9H�I�WL;�u�3�s���7�^D߀kC��K�+�;ԧh��`g���:���#o����ow��y�e�nHu�CXn]@\1ՅnT�Qy���r�S��r�to�Y�5#��6���g)��W�>�6�v��K/��Tv�sP�޼�O�\��Z����o9DŪn���᡹����ʈ�7�����y�m&���^���>}��<�)�޽�&K��s~0c�hBW���M�cO�k{�2��������BYq���s��M���l�t��C��=D��bStr�f��⹕+V�
�cx1�CEB�ֶ	/�4�V�)A��R�ȅ��r6
@�.�N��e[ے��j�zRw�۾��`��\�c[.�-�<�;�OB��9� �SI�+}ɛr�r�3�"h$�v����s?T��ۑ�6���a��0����lY�!@�l�u):y���la���O�ke>��z�==��A໎D�1:�_$�Ev�l��I�V�δ\Ʒ�y.ϩ��*�U�k���k��@�Y����U=�}�SI�kK��O���&��Q�mA��8�J�r�5^�_�4T��:��cmĹ���E��֎W�:�J��oFO��(�sT���n���֒��~{T+ݰ��M��?G��|�~�bw��3�ǿ�� U���1�4*����0�p��sQ\s�7�#_A����kw��/�1�|`�\�����
��U��2�<(��0�~�'�Ļ;�p�;���Z�q#ǳZ�[��K�o���< �c�����ڼ®˷Ut���r�W�tn^�Vs�#���S����)�ddru�Z�k�~߷1Q?[��Iɨ!�Ѻ�������a�u��$5o-pm�}t����q�� ��Im�#�SO,�;���9$��X9�F��k��4�3���Eq�yv9�,!��4���Uծ2���-us��J�q�}-�D��b��{`�vS�`^�{h�y؋���{��W	��Ժ
��Z��Xa�-�췪ɫ��G��1�Y�*�q_7~����9�R;2�����B�B+yi���Ke�Ek�>(P>��=B��ޱ�ow_����J{��L���F�X�f��ٴ���Ҿ�G�H\���]K�����o����2Is=���sק����~-/%�	��ۮ���F[XWy�e2��߻�ry��S���p{��|�ʷ���r�v���Ahv�⍇������/�U�Ml���է˶R��W�z�.[�� ��ܵ�d���	.Jq�Q�Q;u1__%K(�����(�]�����WT�5Z����]՘�t)���R�
��?L`N����W����<=����ӗ:y���t떗z;Y;}�q{8�!]%�����G���=��-�7�.�I�d��"��ݙ�4�m�C�Y�˗�x;Cr�rIVEk�o9���w� �sJiyy��L�^���9�{�˓����%�ȂdU����[�B]�	(s�t/�ۣ�r���S)<S��x�s&��:�Qn�+q�a���ъ�ò�b`ب�z�#ѽ�L}��'�<��r�!9r��m|a)��d-wY�^���q���b���׊�g��<�G[b�j��|��JQ�ev�|a3w&��ӑ�{H8�vہ�����LmC}N����ʶü	� �Y��zfk����pk��{�vŏ{J�]Gjʨ���cU,D(�yAu.����E)�Y�:஋ި�O���;�,{S��A���,T9T���꩜���^{�~[^|�p�kj��җm柝�'�Će�t�.]��|ڨ�G�ů2L�}:Z}�����A}z4�.��
����ز��Dźl[x�_:y��c~��چ�������;$�L)V���}��Ftc��k��l_�ػs��v�藈n���T d_��\ae�ˑ�5ͫ8�_q�|u�\BM����l�O���;�6<u�W2�jS��o^v;����@u�P�%�g�v��=���+0zCB�t��pl}Cs��{I���=s[��뛲�7�}�a6�]Հ]�Ly� ��Kv:�Y�{9f^�ZA9Ҭ��WW�WY�a�qQ��l�TV�:3��׶'�����PkZ�8��m�q�PƱkMm���窰�\3w#n�Ȫ�]�;�g�-q*.w���������� ]�i�ɩD��G�]/�5��߇���}]��\;�R:�~��3s�t�j��8�ֻqy�Hm%�؞����~�FBU.a�w��ꜛ�u]�qpq}ݖ�t��u�;U�1�Je���/�%m>~�y�a����c3�z��w�]�v��)�;��9�[��;�z���s"➧��9��7g��Q���EN��<Χ6OM`y;��7m@�a���mtm�խj���.&ޣKm��]�_^'݁_)	*����N;���vd�cj��1��):���~�澢���2�/a�cr�Þkg�.#�]UfH��9����q`�PYo���K�t)�ߕu��͖��|k0�z@��"�f;�dT9���wD�YW��o��W����n�p�v�����T󎽞;V{���oܬg0�Rʤ��`71���"ߵ�<�v���������]7:U�1��Qgm[�@Wd��2�f��gHt&wJ�j�Wg,W�}��:�Q�BB�\l��弁�~�W�Z���:GLsٯ���kWGf�^����g(��M�x�_����� �&��܋�S����ne��P<��gk�mbڏ���Q����{�k��yp�����ZnX:�����!�c2��}q*�.qXǰqF+\�oa��(������N<IF���^?�gm�����̮�<�;��ó���rl�Э�6�Vƽލ�T��5e����w^?u7��6��ލZ�U��y��IheW�{9��!{��>��3�wE���1����h��T�j�;z?���؛�2��~�}˖Q�5�WC�|v�v�	pwI+�[Y�����k�>��gpS�����>�m�����yڝ���Ոm���~q�0�{w�R�b���"Em�b?^?9�����*'�|ta�"����3se}�]�*��z�3}�8Lo+.^���	��V%ƇOyD�{��-�6O_�R�.�@)k;����V.�:m�y�(��aӣ�4�Y��{o{�Ŋ*e1��ŗ�-ؔ'm�kx�k7��ć{��J�K�����aD��N����fvC��wS��3����������7��j�w=��
TW!�	�'�PgG�Q�m�:�"�p��ͳ�n_C��98�62�l��G�4n9;!|��0^�A���(yZ��]��ټ���5�[�s���[1՚��*�z�i�9������v�K��3x���4���B�Ɔ�r�\.5��=��]�+�1��:��8�}y���Y����䩻��ZШ��w��{�:!����z�;�T�)d�hP�}�Q�=/�WHݫty�]��}�����M�5%�����\թ���'xV;=���7ӬX)]r׽kGZ�ƫ�*�޽|�wi��4ڵ9�=w��o��K}LvQ}��/����Ӷ�	��ݝ�$�d��Q����z.�'��\��)P����#�I��ҟ�묱8�7=7j%s���+��G|[�A�%��ݖk�+r�dޝ �h+.G���b�'�Sf��N"��z��;釒ܤ����5�I`4L�ӛ8ʏ�ۙn0�w-��og��W�6�c6���1jcw�!�׏4���6F9p~���&�y��:q��(֛�����J�\e�
%��/�i*�AR\j.."w��K�eP��c�#�}��5xQ0NLj]ph��~�_3�WfU�px��^�=�73�>sX��U:W
��Kw�����]�s��>��O<�Ppt�K�~y���gP��[ɚ�ڶ�c�d[��s_t���OF�ˈX��(zm�$B�[�򛦨���m�_*+���̸���S�sGZO����EoV��]ۆY���jUu�ʢm�@��2�<ˎ+)&6�o����&mNGT'��V�]`5;=�r����$?�}F�m�]�c=�����cn0�Cvʮ�Ij�^���7٭�\����ۣڄ���V��,~�N�P~\�г�0/R�@�ٞ%��%�8���-�������kB�ߊ]�W�~�1W&��=�O�z"��[.�5�6v�׆]�|�j�]�MwE{�3(kZ�Ř�T!�\��onßZ]$q+�6�טnl��g*.z�0�K;�s�j5G�ղ����lV�=��r'yJTХ�n�]:}�A_#N�t����S���E��V�ڙ3c�|*z44�s�+p�=��؜�������g̓>�N��}���{]^5;�#޻�_�n�d�:{���f�5z��Wد��s�zu�N}�8��:�m����IӠ�c�B�[�U[��d��/F�qxR4:w�7ӟ5>z�~=6�����Z������8�5
w��z�Û>���x{c&��q�;�}\�QyꡭϼHY�^G���s����ք��~�����]����f=�R7I��,�_z��ɝg��p�A�vX�;�z_wf�[�m��BT�S��޿R��Ǝ�w�}�%I	N�Ck���	���{ y-%u�<F���(w���~��~��0�|�~.%b��N�g���w����7(oy��O����8��ʖmy�o�o\k���D�l�{���9�:*���v�/�8�Y�~�EN`�[������c�nV�q����}D*}��U���ٌ�>޾g�Y�vU:>�F�W������-y.��ѳ�.��G�Y��i��Lz��ث�W/Lg�k����#���@��R��;0~YB]�k'�b��t�7�k]e�z-����]���Aέ4�u�:��۾�&�=#M�λ]�xVԠ]�`��ډ��<2���Jj�Epst`��9�:�Ղ�Ea�E�*��P�Ӭ[��<l�K�zj�N�j�Z���
�b�-Sܛ���o�Z���%#�/l]"b~���9��R�%�n|��*�9<�j�e{r��^��� ��f}�Uh�������$�V�7P��xLM5[F���F�Ѯ������Q{m�ݻz�n��{�l��]�k@��$g���j>�c�pf�q��
���W����{���{gi��=��F���G���3���{����G���izHYc��ܡ��u�؆}��|��{F{w��3*#:X�ǽ����z��D�zG~˸�<�g��X{�9��E+�m��瓚���~�{��Y�~X�X)�#9��Q�����@��_Ѿ�����
��N���گ=щ��a�/���:vX�3���Mi\��]~�5߼H��R�lG�ȓ=�gտ�f6�����#���+����~�[��5k�Y�������Y�:h���~ͬ�����N��-�H.���ΐ���<.�]$1ge�c��+�w3�}]S͹5T$C{�e�ڷ���^�g���5s��<S+}~�.^+�y�V�
�2�#2X
"(�ϣ�O����� V��X��&�#P�k'�7yblr4���˼��v�wQQ!��f���OJ��su�\x������ݞٶԮ�j�HE��	�;�1�ݷ�rG^]^wTc����Gu��V�l�4�ˡv�[�E�	�6&}�}q�p{˓�ʜ����U�r��е��r+�M�����/vuִ��5+_ �0IT��]�[A<��w�`�.G0"�y|iue�af�5���NW0eႆL��`�����"��_l��0n4	V�k���W:��4 �ܺ9 W�z�p��ˆ�uǜ��*�o����3���ܲ��g��j�|�Ӭ�����f�x0����	oK[CP����V�B���S'��dk��J�z�`�MB�s��fcC�5Y[Hl]�2�|�,��rDu^a�#�w�n:r� �7M�P^'�>�:�BP�m��q��r�졃w7�,�J�8f��*n�՛y9 ����i�6:z	�(�����d�wՒU�����WS,��N/f��yɥ[QMm���YL��Lu�}$v���$M�ϯ�\F�8#/�>��qA�j��*s�
K��n��E�Ny���3imK���-���ɊI,�QX���J�֌j�4�
�>WhG;�_��:i��03��Ѳ1\ۑ���3�6�7�[R�\`�ho3���e���'*b���xm����[���n��9�gW¥NqM�V�����ŗ,h2�
#�RN�c&7f�Y����@��!���ؔ:���[�chwj)x���2)s�u���,��h�C�*�e��7�R*�ݳ(H��vs�o��b����tӫBs""�X.�G6�4����uh(nEJӅ��N����gKT]�U�e��T\����v�1�%�Bm��ƚ�w�٨\=�e�*�${���A>e!g~�����3�)r�����,�^V�S\¢�T�~����}��ǉ4�睖mͺ*��'p��m;�B�z��%/=LJ�o9!!�-[��t�z\<W,^�SL��w�AWk[da�],��݇���}$���w�v�WWN7V�8z����;e�pe�I�MGY�`'���vλ�2a�J�w��A}l|zl�#?.&���곶���ՃM���M�ƺ�+��U��Z"�]ѡ��nܺ���,xWn���J�F]mN����5��*��T�:(9��]Av'R^c�6	R^������]�/i�:w�|]cJ�9Kyna.�ە���Y�8�MR��a`MWn[�1�s��0�,���T�)+���/
��F1]F��V�b=�"�p�׵���`�7٨���՚���O��5m�&��Lj�Ӻ(�pW�{W˩k���5��fD)r��s���nӉ]v%S�H �5�)�i�;���c�ҭV�
��"	Z�D��[A�j+P��YEb�(�J�*�F�U��\eb�s%AG�QF-ZQ�J*�Ķ�r�\[-J�DA[eAb�T2��FZ)QJ�VVX�mV�Ш���(V�PE�J#L��`����k"[-�dQР�GWV�-�D�,Z�PEE�YZ*Ķ��kmQ���j�1��DF((��U�����cU��¢��e��V,�F��(��(��m*"��QT1b�%lX��UAj�l�K[UYiE(���UH�*�Q�Thت�b��K��������[J������`�V�j
����*�5Jҵ
���B�P������E-���1h�R���b��3-D+*���Ո��T%־���F�qo�) ��;u�s���2<J�c�n����k�)�MΔ�a�7z������"^��׭�sT�9���_Ne��9t����|��˟�1���W����^-��Q�Ǫ�K9�|�	��Ө�;�Љnem�)^��#�nz"��WOx��%�ڙ	�WZS�R��/J�g�<�m_�=�}8<�ǳ3��5w-ʾ�������������-�N3���ͽx��~tǸ�nǲ_��:��W8������ܿd1�)���g�ba���F��;�}���Ƕ�4m�ϖe�K<g���=�G3~ܩ��,�Z=L��jИ�}^ӄ�wu�~Yjj�>����I��SʟGq��\9R�g�%���� w�ې+��(���X�n`���!����2�_�����mOsKO���F�q�*}��O£n#�W~9�t�s��g�I��|8+��f��fn�ǹo>��`�}��W�\�2+�׵�)7�;s���{�c�vv�<$�a�>V�}�>��5��L�����S�3kC���Q���3���?]X��t=q{�G��S�b�:�U��y�ګ����{�� -��-�+Ė��ӵ�[��͚�f��3y��׫�b�`����8g8��}�N�����������1Nr�W���(�.��$Ouw�$��R5���*���73;�N.����N�*�̇��e������U�b��c]p��<Mp�{t����݌���_x�c$JM�4��/�[1��ܻf��v(+Οf������3۵��Od�����C�g���FmV��΀�[��y�IQ�������pк����qn#���}�W!�	��$�ۙc<�"�����]*���^v��-�S����>I��dk������v��r6���dw���Q��D��zY��@�S2���Kaښd��Nz�9άn2�~��~>�B�{�<W#ˬ���}Fe0n��e��Ig�<}��s<E�3�K�O���^��>G��ך��O����]���ɚ��*���z���3
�&Q�����"���7�)��8=�yב�y�]�8W�l�o���`��!#م�5RD�\x\)��9���9\Mz�Qn�7W�܇�L/�N�;ÝZ����}�?��J��F��1�+}t�'�f�M
��K
�/p�z����g+��m�\}��G\?RF����u�%
�_�FG�\�@-��,?7�Ǎmg��ዒ�� ��~�X{��g�7�7qW�����Q��ǷnE[�rQ6�A9��P�_��QbG�uKU����\�W]��QL|ysgF��[����Egw���9*��9p=��5٢�Ծ���t립��.N�'ٽU�V�{�0쮍&�vG}ys��-�j��+:�m�7ܣ�jO��OT�krJ����}+B��S ���W�-����������.}�P/}߅��~�u1~r�3p�u�>;��Y���R��]�J���}��K&��*��\ex�+�S�j5Ώr�'4N߅X*FL�^��o���Cn���M���N�h�H!0xi/��L>ܭ�
���j4���˭�p7Q��
��s��ɥ��Mf�+���ޠ:�n�x\9�DWн%���;l�/˘{�m{�-W޺�����_���ֲ�����C�������=ꁧ���/�h���r�XZn'e��ހ�ng{�Fl�����W��V=��S(0[�c���r����b����ߑ0�͎�zVT&�BG�d(��ڟ��qY#��~���#==�S���~�=X�~��}�뉯G(����+����}�c˦�Ӧ=�Mɱ�2�ߣ&��y3�'\����Ʒ>�"��*~=����	�U!qeߍek�wߕ��^��5Q낑� �93+����S�:�9�P��taF�V��Xۖg|�Nz��e���4����_��\K�CF{�*:�$OIwN�B~���^ˠ��T���I@<����*�,�b.�+��e�.�;y��ǵ8[[�u���q��x��jjJ^�K� ����ީN�q%���-^��n^��׷�\�<���s���:�]˛�ʁI���ev��9N�!LI �M>�:�1P�(�N�5{�w%z�g�=�\<�������lxj��2��&A�7�E���Q�}^�%�K�}��W�`��ߺ����>�|{J�N��~�_�B����@l���t[��l�/@'�g��U�|N�,{�rQ
�x�&���c�v�xn]:�_�3#�L�P�3�,�K�}Tpz>0}����ǽQj���s㊻�w�=_{�W��~����:f�<�
6ET{�y���m/��x[Lۯ��� ���4_����厔<�����o=�;F�q>W��Jw}H�!N�iz�����P5�� @�����}5�5��$ȨXlMw���=��h���֋Nk��Ϩr3����DW���j&X�\��\f�.��>������.����O�γ�R>��ب�~���΀�9󭻏`{D�Dq��C|_O^�ܧU�O�N>Red��e��BU��:�Fl���.�=~�n�{a���X_@�6��_���C���4kt��}?5�_�n���KS��+�V�\d�9��:���#���\��:{��;kḋ�=9�l��;�*ὧam>����fRr����Uܽ�p��-TO�%��h�T�t��f��|�ڧ8.�z�t��'{bb�P�.���H�V_l���S����]�eG8��kW(/v�G.���[K �{0Vf�ć0>�$�9�^���"�t�����5�h��0��o���9}q�~�u�Ċݷ�W��j��5[�j��QGۄ�=���(h�������}U}��~���@kw
z��#|n^.�Ԫ�����M�g�÷"<�G[��2#˅!�J;�gf�Ϊ�SyIN]_�g������n\��(ꙋ�����|���u��
�{��RQ��$	�X`�!�4�v*ۯNT���]|��F/\m�|T�/���xr�2�����%⸸kjY�!{�d�D�u�z�q$�&gҤW\�r�F��H��7�b�%W���C��oަ�!p\�ׯga�&kq��JOW�k�U�*��9\Uz��M�im��=|(\7�lW���O�F�s�Χ�p���l����1���y ��&a��Tb��,8KGّ��G�ߦ�j�9~�]��4=�+�~;������f]r�C����xթ��}^ø���"'�.{Ϧ�֣�f��j7��w��~>9,�������d�'"e�L<_tV��D���}s���s���E�6�������J�t����not�;�����;��Hs�t���<<=�!�wj��Sq��M77���e�#��^rsR�{]nTD���s19����!��Z^J�6��Xf�� ;�fB����$���S{�Wx�eq�Fl�{���7�Q�yUx���Ly��u �Ή3��g'���e�)Z��z8g�j�y�C�i�_o�|n��:�׍�[��.rc�������M�k����y����A��V�q�;SN$U�d�zMf��f�,c���A��u��φz�{��6|���-�l芈�	Vo�/���B�N���}�5ρ��l ���i���d��ڳ/y�\߰{�ꦉ�tT?eؑo�kE���h�ɇgs�UƓ�cE���y~�k���yO����xQ��g����Q��c}]R�8:�Ê&X��ű���3ޞ�w��[�-^m�o����f�vP�ƽQ���_�����=����j�����IHKFj���u�:���L~q+�Q_�����Ʒ��q��|V����_?7q޼������η�+��gЈ��J�X{Ņ�T�sjPg]PQ��8�3�Lc��Wyzn�RѾ�>��\nG.��,ؙF�O��0&���7Sson���^G��{�)��cW+�֧g��+��e�º��SWl��F�T��e���3�r��h^D+D�r>E��KfR@a+��,��y����)I�{�<�X�X�DMw�C�OB�r����S������D1z^��Vg9]@Kb>��ΈO>�h�Egs-�����7�����Z=�	��s��7�B�܈RM�w��FSt��¼^�joaD�5�ox{0�h�#=�\?��|7}�4W����/"%Q
�	MA83�#Є�v'��t2���v��rT��F�\j!�Wn�i��A3��£�n�\?Uz��@Zgu���5p)�y�n�������U �xރ���~7~��/ҫ�W��Q������n܋�΍�2Ū����}�o�'I�I^=s
~��&��:0���@�����U���~��DJ}�_�3t]���o{ �C��ωD�I�su�|LlEt䚌S��e������[^���{R=sy9v���}C����h��*dp��(���u�w.��t��Ӄ�^�ɛq�+�n��}�����'��:���7���xc�4EB��r�X�3Ƣ�*M�����,NoU��Y�E����z}���g:��������[w����qp�M����8KT�
��|_���u�UzF�7�\�d�l�'Q`,w���zu�NB>�Q�θ��=��DB�zz5�zy�eq�;[A����7,ʸ
 +H�㙁M��J�5�k���NDp�/���#��tM?~�MsgOB��#S��4�*���RA�JcB��>+;��#��x��̊wLTvuX3%��7 +u�m-JJŗUQ���u)��\�
�O8��&|�oy�`.4n!Г����g�r���p�ɭ+���k����j�;����X���^G���$�*s���gs{s�]��k|b����rl>�CۓZX�ɝ��@7ު�׼H���6R3ӯ����qbJ:��{�գ����n=QJ�@~��q�~�g����c����I�EȖ����D��{�Fߪ�����z}�u��ǔG�وxo��1�A�!���5
�W�_�����;���[K<�^�۸l�yTy��{NG�X]�����K�lb���g�@���7ӹ>�W�S}�o#�-J�ǲ�Z��E�F�j5�~�c�6o�T��v<�Ey��-NQe\�8م�9s�T��䗀�#�ڠ�ex��B���S�$aC�U���:{"*})e����WP�7�觻JK
�*�Tz���՞33__.��=pRe�6*̟�2�e���_�s?�y����!~��q���4��/����_�����{��C�7銗� �/��m��Y{����E=4������@V��)�.�������\�'�x�#�m:���>����k���l�k!+���jT�8v��'�� �fE]�ب�;ub������)ԭ��������מ���О��`��ů�J7WE�.9+�	�r��ڐ*z2a��x��f�t�P.fp����W���W��[:l�܏_�8�`]�+GC�׍�]�g�k@�d����52�z��c�p�������k�N/��S�[��^�U�p=>���.�QQ�E���@y���ǰ=�MD"_���Ń�2��ۙ��;aȞ>��q�Z�d�Fl��eq~+�̸�R��r���3��=8k++����f��{�����~?�������ۓ�O�r�^���s���`RW����E����[�neeh�ݨ~~��А�S��3�j��iB��Zn:����{*e��K;�
Va���U-Y#ЖR�r����A�����+�)Y���u�X��~Y����B�Y-mov9y���3=	]��z�7�|;s�;�������H_љ%��,��QCŹY�d�2cg�}�<��}�g�VV�/��wߩ�{�~/��:<�����VF���
,ߺ��m_�$f�)���>b)�ǯ�E�����R�QJz��<S/�_��*�B5GT%q�Q�Y�����J�:_�r��OH�|T�g�G�mԏ\7�CЏ����MA�{$Ua����K���ZZ�-CtwTA��Ue ��_�X[[1�����u��u�s��r 9�ƺ�O{��n��x���P��p�i���^V�ʫ��@:��u������Qٮ��ė=%9��`�YBMُt��UR���q8 ��K�'3��#�0��Q�2J1���)�I�l�py�GR��!b�GNz���n����InnS��K� V����3Ӭ�{ ��0��ңW�a�%��	�g�"�ܩ��}x�fڤ/ў���*�$q���#�dp�T���°Z;q2�Lu����:���^�++�ϔ�G�`L{ƽ�.�~����� ?)#\��j&P\G�}p�����ޓ���Tz�y�"i�i�ҼwN/K~������G>u���&ߙ�fe�M{���I�1���ѷ��us�2+\���S�Y��s���ӓ�r㽲3��ny����ݗ~����ɨG��	�麎��V��zNk�z�=o�c�s�h87ՠ��)�'��y��~�G%G��mX�<�#c�%Y�/��D�B�Nፋ�����u�g�2���}"���w:��u; {��Ş�Uy�:}���C=�pw�Ӥ�r�r�ῳ�P�s��T��k=}�0�Ż�����呪��߯�����ᾮ�ފЬ�9�,g�������T|E���͓��p����D�U�
)5Ts[7�싨kC3��;s�Ei�jEdv�v�5k�[z�s��a(Ģ�N�v��Q�3���)w6��|)`�M�;!2�o ���r�Շ$Q46��It��R��U��]�1�S)ä�k���}k)a�wE$d�(	�]�/\��k�����I�[O3)�5U�1�
�s��ܬ�}�������1�5�E�GR�>%M��^[}XK�<vK���.�=:a�؛t(���u�D۽������8�Ү%RV���݅��N�E�2����O5�;l�bW 2�_%�RKm�u/N�9'��5�S*�к�hx��n�tiT��3h��0ʘ�ז*]�iu*��c#���o�LUNߏM��K�ψ�~$5��"ᙔl[�^'��d��qQTt��c-w<�}�.���J$�;�*��I�t����ٖ�꽷���YC9����h�97Q����,��6#Vy,�w��+0.��y�Gx1��H�@8�t�(Ԩ`�U���t�R��BZL�������g��eF�4)u�ú��Hx��ǕA�����}f��>-�!Gn&F�0�٠��ux�i�u-)�TN�W�qQ6ˎNZ�b#�n��ݺ�e�C��,鬧٪��el�u��y$Ș�:|zB�V���.���51��s��8��'#U5���k�3�۷eQ]`��*U�k�:kC�:�^+^Vƌv&+ 7N֛�93���B�Go{������
�*���tN�ن��a�j*�R����j�ː�c��
NiVQYmVQ�r�Ѵ���M�&��^�A�wk"ư�p�{�V)|�W6.�����y��+q�YQ�� ���P�>����F}�f�F�V��Om@�Ԏ�u�Ә,U� 4��+Qh��7�6�A�cÌ������$ص���0՗�85�Qh�u�R%�w=��옶٥����l�v�N��&��L#bW_ɰ*�����j�:)��qR�M]���`a�@I����U���2}D��ސꛝ'С�=�������I��M��Ֆ��9R�f��ŸC�q���8v�K��Dp+�FN�Ւ8B��`��,v�vQ�wU�l�̺۵�{�5�*�B��L�g[����p��]���F��OE;��>��]�C�Y��!|��ڕ��V��s�=�v��p�-�d��x��C�&� -;6��J�0gk��'Y���$��U%lzhV
'v�q��6�%���B�X�6�R��z[7�����<�!q�ѻ�����_j�u9�|9���n ��1m�F�@����Z��e�-|��Ʋ�qWϖ*��W�T����c��1+��VoAD��]8tT���ko\�s�tf��&t�(��GC�{����w|��<fZ��E����EYhQE[�LFj* �AJ�b�KkJ��m#��*Km(�G.31
�E��*媶�*�,DT�T��V�ڪ��1b*�W,�2���QTb(���5�AX1+,Z���j�[kU�V���,���lDV"��X�im��QQm����5Kck�D���[mV�F4Bҕ��֡U�Jыm"Ԭ��V1��Z�QQF*�F�0Ke�bƥ��R�cP*�D�hUR�Z���F��V��&4��2��1������(���YiDX[X�AE-EUTQ[kE�*�h��,b�ZT��"�R��J,b�V��lU�,�e�m�%J���1�"#m"*"*EEV0b���kDAcjUV�(������*"�"Ŷ���Pb�VQb�������,��(�DAX�i(!kh�E�*2�Q�Ekb"�T,EUU����u��u��ֵ��k�9�3���L�b@s��yNG|�"�6����]���E���a[J�qǚ��g/I+4��=�S�9�쭸{��Sѧ�5��1��^'�ޭe/z�Qi���eN���u�zhG�7s߯��9��&��ѿ�1�į��#�ޫ���/=/�iط;�Z��N�354���焕����7�������a#R���Sb�X��~<��\ꃱ��t��G��h��Vĭ�����ӵ�:}���㱪,�\dL�(w�"��5<���wn��7�����uX��9��P���zxx����|%����+�yP�ƫ+/���o��J�������*��7�-=F��_��?Gu�f���#!�[7���#�u������A[R� ����t$zui�$7�"�g.Y��c�^OzǠڭR/2!��F�%qN}I�Ñ���<+�n�[�W����&��g�ŷ��0DL{20��9�����~7�7qW�X�t��Q~>w�s�t���Y]�@�G��>&���v�&=5<Lҝ�ѐ\�N�2��~����_�+y��U��0Qe-�|��{z�%�������gĢj$�*��_�^&&�rMF)��d#Lmdxέ�_�]rg=]ki̵\����\���/�#FXO^��r�2�H4�����rlp��z/�7z�j�@Q�۽ް�p�:�f��ۄI�ɥ�C.�/tPr��K��SJ���-��rb��\����>���|ǖ1\×���t��2�B��N��M���v�)ql0"�oF�j�2X�B�U��M�󝓃����RbxTA/��"n���n�W���I�{O��&�[�|�ϲ�1K�+���~t\/m���:h�^��\��+���Ɉz��<6C��M�D����GmǅCy����Ԝ��@�O�s#Ё"~�{������듓:d���U�5���������,{�TmK�K_��dzu�M�zF���uīs�AXVWwf_t����W[�Ͼ��}���l�1�5�\FO�i�·zr5O�\k����:�Ja9�^{�7䲫����B�x}�|k>g ���p~C�fz�Y�z�𙮀ב{,r˙�zA����
w�n��G��Sg��}��_�]e�����/	늨~5�����|�q݈{]���}����;�wb7>\����3����/-���JH*vK�桁~�ܳ+=1�U݇7l���y�<���Ϻ��Ŀu�Ϡu;�����G���J�-NQe2C8��\H�X���Wt��_q��d1���7��wjģm�\{�6}��������^�:�[^�$�	<_��r�w�fpS�RBk��u_��m��j�X��*�YB'�:2�-F��dR������8�זW����՛3I�Le�p�d>:c�ۦ��z�=d\��\�݋��|r�9q�X���Dn���qfܵ�L�Nr�����|G9K��-q�Ǚ܆��w��Y�M��O�E�~�_�ϜV�oo6/����zѯ>̿\,����_�E�D��w*H�YE����^��ة�	וVd\���f�|���X{���D{��w�ȑQn��|G�baz��D��^���@{�x��;��7u�^�Oc~0��5��r����*<����`��K���ِ��	�k�T�%ؿN<�ٵ��Ǽ��
g������+���*� {���~�D?ĩ�]áR u�[2}�w�X�|����l��K��6��7����~�eC��	�p�Tzꇭ�T�}wZ���)�3�}��S�Eh�77>
�kG�2w�j#6��3p����̏b�Qr�Gz��dp��߮������ۮ��K��}��8o�^/NDI�:v|?vN����:���߲<0���C���9ky7��Wu�7yV*��1]�;��v���y��,(�٭7��@w�r����Z�<���X�m���-��I�{M��Z:��hH��h��N�/�UC�Y[PքO��"}n�ھ�3�oRʹ�h�����'%-/�����:�ק8"T��C����4��|�b��J7��9��iԔ�2�����:�ڱЬTo�܆lgSȶ��EQl5�ޗ/ta��;8�kw�z��K���]��3���P�J��9�|K��Nx���;���-�����(m�2�����������i�C�#9�*��c���ɝs쭪	���w�߯�r7��_o���q��yl�z����Rm��9]Ң�=�u\����)�}t�r%��{8���؏�׋����'ˬg�w=��m���]{� J5�;�`LT�����/jd{��և��3��S��g���L�}
�hǬ�t�7���Ǳ��v8�Dq��W��-�M�^/rY	��w��..��ʪ�є�װP��Lz#�f�+~��������!N��<�Cs�3!��&2
�,5z̢Dl���ܥ' 籜~�u�Hп�z�9��R����t-��7��@l�5�O���t�s���j)u�G�/��p����D{��U��ߎzv�߯�{����I�ίm`��3;�fZ�J{�xy���Q}DS=�4�r:U>95�Q���s9��*r@Yټ:��4��_wy)��>#�aD�.+bn���=D;+L��;�،������n�naO���=��9���^�4i��e�Ń~�h��苜4uG����Zp��=�QA��L�@��xD�of=j��3�ו���%�͕���]5�|ܮ�ZB�����I!��[;H�%��4r��uIB��*�2����8�tM��ײ�Q���!�QԞ7iW*�����D��2��Y��I�®*���&�Oa!��DM�5q[��O�I��]p2�1䩨��"G���m9�~`;�]6�l�=��Տg��Ew��$>9�;P�en�w��+��;�r5��U�v���˶��v� W�����^�-I�����bE�i��x�/�)ڇ����cE�L�I��Lꥫ��8�B�]��>g�:� �W��>�\�R}郧����p���Z�:v�܀ף}`�uVwsU���ї��d�\�,���z�����7��g�_�9��W	���=Pe��yY쾝���h��#�T�X;����}ig�S��w�C:�������(;�ݗ.*��7װn����هѻ��y��QQ)�8\U0&�X��g_�+n�y��?'�%z<�-�\4���ў����ǚT����^F�����ό-�Q�>EM�0(�>'p�]�\�+���ͥ�9��^��t����D��z2=�����ȉ��F�S�W��j	�;�X�3>�������4O�O�[�낍E�uǲ�6r#�%���#C���0��e�!�	{�G�or�v������{7�0�u{{����1YtLaֺ�Z�ݸ��pX� vN7s�@�R�+>ǳ}e�`��`��(����}Ge܏�-e#������*�^����Oz.���6��Sx�#q�����͈*�nu1C3�T�7in$��#p�+�B�=��n>�h�r\j%qW����:�2������0g�-��'�l׮O{�@�)�����P����2S���q^��~�L��:f`�~:�n�����0��n\A�o��mq��]��|J~]�#gԸ���TC~�=Vo�)1!uz�yv��y]�z#�u�L�z�@wv@�s�x���W��C��+���MVѽs�ݽ'�wލ���]z�.�o�u���t\su~9�t<�!�����H!0x����7P��+t�� *�ɳ{j<g�ڳ|��,�=W�0�:�P�TQ�^��Wf����%��;[U�^�z/��_��.����Bx��]��3i�ޟ"f�n�ǽ�~�TYG>�\5�wσ�8W8�/&�g�2���Y^2p���;>F:��'kg4��Q��z���(�N2���Hf}���d�y��V��}�Λ�D���oӴ�\d֕��p�˝��>�_���
b&�T����5�r�~���k��ύa��g �\��y�*��3���ɝ�t�p�s�=���k��W��a�\���A��	[�h�?)��]�w;]J&8M%��.�������+u&�z(��׶���GT�FK�s���k��7m-��\<E�f<������\���X�k]�����\lvrk3���4��AyN��eN�R����//�^�y�����.��\F`���xO]T?��t�/����z�`A��=v�K��z6���;1����9�u�{~�W�.��p�DlL�_Ia)zr���d'���t��U���E��~%�Ty��W���es���;R�}uK<�o�o����2�v��w�%�0��xSQ�Iρ��L����S.��<�zR7��>=��}��ovGm�L�@�m��㏔�_�_�j�f�; r��Ш.Z&�X�;�>�<W­?[f6�>Hz�E�U�gU^��ߟ!���}��YN����^��-�0a���F�	^+D+�5σ+���x��<�׺�_�Rg��(�q퓥[ܸ�~�i��똘^���11O��S��+"O/f>��z��n�g�y��<=*k�G�i�����ˉ��*"e�W >>��=����+���oUn�|z���7�#܄ǰ�k���7W�=� �|� �f���,���&r�*��˵��K�x���ü�!ߧd��}��n��:��h�)��:۸���*�J��*xR�2�{�2��:�p-�ӓ�LB��JXR�0^K�\7�½�5�Tv�q;71��@BV�g4i'����L�Q�YW7������mgFU}]2,��	�T�V���Z�י(E%'��q��T���أ�s�����}H0<���n&��^mhw��3_v����"ǟ���'v},�ՃJ��q�/RHZ}�ں�&�*8̼='������;���N��f���S��P����}){s�.��U��0{�]�r!:w�4'>^۝0g������=�#�-���y�~-;���u홭{��]�����W��h�߽$/d�K^����N�N�/��;+u3�ؾ��۸�u^���F{��;'T���j�f;>���9�~�ޏ:�����P�'�1�T�X���W����^�=2,/F+���L�dV��D�����~�K�}S���{^x~���N�����c˒V=az�.���=uL	����_C��_����}OK�~+��(H��'8���[�i-C_a��z�Rږyl�(��޸�`LT����A��6�G��և�۸�/��2U�.Ky�<�m����Q�G(�K�Pz@�q^�D�Q7W���=qVǲK�ۚ��ݞ��X�_��}x���vǐ+��u���Y�U�P�����n�*�؈{�Y�l��CH�-�tK?�f�k��=�qs��Ò��B�$8:҆fTˣ���1��tY�@,*�v�Y�R�'=V'Kk+���<]t��\=���7�S� ���&�:������T��C�*�Ӥ��J�z.�M%`�S�����,��؞�ԑ���ؗ��ĤVd.y�RG�ïRG!����yd�.=�����0�>E����܃�*|fڟj�}�����E�{�|j��k���~*=;\
�~� ;���ȻX&�1�����>����I��f��-Q���wNAR��7�q�U^7����NŹ��5s����%���F�nI�Y(ј|Q�c�3�C���E}�wǲ!cm;�y>p@�����e��r��'��F�%�<�m����&�d��/��L5���]��t��5�3I�]U�w�>��eq�U�[�/����b�s��3�O^uc��Tw��$1y�P�q[��"}N'I��F{�f�x}�|��|���2��Rs�@s��	�gGzO�������F�'��<�S����P�3j��������~ c�W���#��y�>���ﶝ��q��߷�1�L湅�` V��c�8����v��s�2��M�l��u�1o���5�٭��v�X;/�>�ݹe�#p��z��d֗y3����t���U���?ᯨ{O���$� j
��Tf�=��,B&L|C-\����f�J/F[��Su�R�1л�;n(S��X��q�+�.L&��J���˦7Y|.nl�R-A 6A���B-\�V���U��c�R����z4n3�ж���.�{Bj�tX���SO��|7c3~�������p�����6p4��ϗ���������{���7��'`ME��c�����{v��S:=������>%Z�������͉�H�*v��G��'���k*���6��\����n��c��|ǽ�ё���~��yh1��C��q.��w�H_S^7�=�撯0��i7�#�����yd{a�W�r�1���{��cmJ>����5�!����o�^S�'Cf�+���@�d�}��
5�+��^��?IE3������7����.F�=@z7i��� y���a�Z��#{�X\w~�~5��+��n�z����*��e��6��uK��;�i:p���}�良U9RA��&�D�9��ڡ�9���z۞�~����H�s��Ay�u��r_�Wީ�	�*@�>%Q%�Wu�+���5[D�j�I�0���W=�j�:��)�;�jN������'�x��6L���눛�}�ǝ�󪼧�k����t��/O����Н���Ϳ:�!�ݏp��%ʪ
�N�w���[�� :��R=1��.���;�-]�]��F�<��ʥ+ݷh4��-o��%zޜ�F^�b�e=�Ռ�{��M	G0�<U��������*ps�;�*��[��0D��iv�C�7��!Yضq7���I�i$r�f6n�ǆ���)ND�M[#��n�MU�}�ۗ�V���Y���si"Em*�I0%�k��+�PʈNyI��;V(���l�t�\��,��@�_t��Vc�eԗ-������u�b5�Y��qW`�ƶ�b����pݏ�A�NgT�`��M��7��#�vN�Z�,d"l]��y�1C]�s����۔2�簬B�N�q�ˠk�"�/DgK�+��
a��tÜqs�pL�Z���\�u�m�tr�,��a!��p9��9+�L0�!� ;9��^I�W��{�bs����A��/�1�n�-�JkC�EŪX]tMDbV�n�F�����n:7�Z������Cl�R�����#r��qgÃp͸��Vʰ�څ��K[+-������a�߬��т���D�L���;r7f��}��p���άݔ�Xj��n��/a���v,�f��P�n��Wu�PE����U�����X�iLa�+*����er˖�lz~��9���/��W�_u՞�����_2Ґg4w��#��m��.�y)e;:��q�*sk�lF���M�s���(r����t>��wxn���C��d��o@;�����|��Z�[�݊b0��`S[Q}�(���,]N��ڍy��މ�t<:J��u�A<7K���X1i�P[�$ݶN�������JC�葻
+,6�'�JAX�����NCeQi݌v�z\Om�4MXT�o!��r+�6�x��_aM�8�� '�pZ6$$���7���Y�;"m�z/v4.���Z�6ak���tx�u��o6��^j�_Zwۑ�-ΡÀYk��Qn�#c���+)��uY�Zum������ɼ
�9�.Q�I����,=u�6�ؗUo9�s��i���fbT�l����W�3�|�Y��93�U��-QU36:���틅�\���`t��i���)�p����Jn�}�V�c���m��*R]��ywt�-���D�r�˱P	r�U��ލ8R�p�5T��D�m�[W��0Ԧ*w��t���l�u��E�ƵWc�oBV���Z�MV���1'��jT���Y��-�r�yi���.0`̍� �80R�B�1��t�{HY����q��ͫ\f�!��47N7IP.�̮޼n�T�d��*�D�����u��3Q�k��lRН8V����lw/E�h��\��Ư5�	���c���g=��|�X�J������Xk�1��H�m���ȭ2���q� M�6	ᘹ#u�� 1Τ��)�o)Co0��N�@+�ڬ�'+*�R�f#2��Ȇ�9&e���zw�M�|���n�{���!����Yy���v�ʧ2O��P���AD~DUTE������[j�EX�Z�*֪��`���B�PE��3Aej�	�sX�&Z��Q��U2��*(��* ����F)[QTAT���U��e*�U�UPEV �,PUKkV�""*K[�bV�5YZ�
�Qe�#"2(V�km�ai��[`��ikKh�*TFTX�ł�E�Z*�1��X�,�Lj"5���1������V#��-,,���2�U���0Q��������ŋ2�e��"�RذTR�Q��Q�4Q�+���mJ1b�,.`��k**�h�,X�U��m��b5j��-�X2+*��b�UF*,X�S-�6**,UTb����"�bTF�k���TTT���#����D��jUDUQ)�U�8�V5h�%��F"*�",TFE��J��Q�h���*�
 �|�����5�ұc:]�Zz���%v("n�G��PQC�;���e��PΫ�����sm�,�uv_K9H��M=:H����-K~����;ͯq����f��~7�v熿Uzc����G��3Q�y�l֮�"��z7$��<����8E�WNic�2�T�1ׯ�w�Z�&��C��0q�3�z��Mzt�y��}�뉾[gM��N�����;Le�5�vυi�r7Ӝ|4����>����{��ח����Q@��j7�i��r
�a����ʷ}ic��Y��,b����ɒ���cU��.���;}>�!��u�{m֎~�C{ˬ��%"C�{b*���,�=��Z��V���1�e"�"�fD��tc_z����י��!\{�lpȏ!(u��=�=J^k;�VawA��
UR����f�����}UĿuC�r��=ҙkb�~j�{=�x��جվ���?F��xs#é��7��v��J7�O�"����'�i{����T��k���}��ݾ��i���٨= r��Т�n2X�;���T�_
�iį��=�;�d��j��Z�>�I�^�w"��E���7S�\A+�a��xẘ��fH����־r��c�]q�%mvӶ����,���j�655�'KS��ь�ۧJ.OKuK�*��1�q~��y����u�m��y K�*Ӳ�Y{q۝-�G��oi<P_S�������u��;$���<��HA(�S�+OJf7[�.U��&�I3٢y#��ﺘ�'v�c~��.o�$y�{s"`W�ؤ�GL^ۤLy�XH~�d������Sv|J㻐xz�����>�*��
P�|��ć�x^��z��pr���ݳ�4�Ϛ�6wA�}Kմt/ބj�O¸\{ʯ�7��=�8 U��6D�G_0UW�_��H蔖.��$���44o�h�Q��5�l�>���5	ب|�F��=��U�U� ���<ގ������E�ڒj�+c�M9Fmhw��5�Lq����_�ٙ��ޡ[T2����uw���w!����Q�q�ّ�;��̽9|��Nׇ���>��tV��5��f%����o�N�x.K�[��`޵��U0{�0��*�߽�:c�a�-���yy^�Ļ~�;L��[}��y�9�@��ڭ�Q��ޒ3��h�^�q��BE����`��C���!��My�<�}��L/Fuu����!���쁯��s}9�ݾ��u��v����a��D�˽����;�_xѿDΌ*d ��Wq댙�O���&r'��n7������~��3��n{��Gz�<�/�#D8XR��b���5ΑQ��o-M��v�X�`b4�4�j����Q�Xf-m୸��d��B�Y�z]��)���zb"���]��p��N�*ޗf�T��x���L�
����oDC����p�"b��d�Y�7]�����]G�f��a�T���\;��i3�R�n%��<���v��˘�[=��VbF|4�>���o�J�o�nYy J5�ze��S��o��A���G�
�ڞy��{�sK�{GzJ�ё�����n%�=���f9�rF�5(��Ш%��͘����y�Rγٯ�1Mr�w^�����!�G����ƻ�?H�\!�<�G��$��ԣ˘$���n��|��u����n����u/�ZF���$_�P-����wB�~�M�]�4K���s製�vy��} y����Sß��ϑ�~7��{"�"|��o�x?M��r��r}$�����Ҵw�EϏ���3�#s�Z�%�Ý��wN/M��Q����M8\���*���|��i�>�m �=�&��Rj&a�W��1��!�\�25��o|������0(Ca��>��O�C���s���	鸆�T3u$��Vv$�>���j�oC������q�z�y�ݻIw,8�3�ݴ��>�A�\?:<n!{jǲ� ����:vaz�E�b��>ò��K���,v�z��fy�ih��<��o��O#[�7�%�h�"�z�����MϚ#h7@cF�\�}5�y��+T���K/b�a,� �U݃�4��&+��(Hf��5ut���]XV=�x�K��vg��H�u�����cT/�X������U�F��� ����s�>Rr����˱B�	�Qޓ�#��o�j}1�k3�~sq��v}�P�fp�/ǧ:� �����sޝe�<k��g\��C���*�9|+�;=�]vf�ǳ$��>��φd�B茟+���`o�%�X�?W���ӈ�y�������^��.몝|��EY�u{^D��⬜8��z��}�Z]���`�ʞ�X��Ckf�]'7�k���*���3�?���WM�:c�������(�8JD�`��T����c	����_N.�4��r�.��-jW���>��Y�����|�����ļW~��2��j��ND{�^�Κ�
v�&�����w�]y����Ͻ�Z<�>�^Z#��o9�q��b�Nc u�&� ���x��)����_E�uǲ�6r#�F�ޮ����Ng�6:5Zӷ�gw��oӧ�s�xy�����c6�>��]�TSu�H���S6�G�*�u��{cW#��׭��ܿ]���E�����U
���9���S���Q^�@�͏S�,��"�3��6أ�tiY+��5]�7��v����>4��w[24-]!Y&~���{����m8i��^mG��j���[��f��{�)lS��`�vG7n���A�45�o��,�/Dy|�L�U���Z�4�gB�b��9����f����J>ͺ�Q꜔ND��\LL/U�&�����;U�-�U��=۫r�V[�>�[�=>���{�9�_�ے9�(�����S�+�ği�UJ�Gg���m{�q�:>�:X��i�����ߦ�WޗC�s�S��2L�_�y6#�E߰t�9��t���C��=q��N����_���x'���@��9˱ᐧM��&�O��YW>c�;{/UW�U�ѿL����lyܘ�}�^�Z&Tv�?��/�>^�,���ĵ����-�l��ϧ�}��p��IG."g�i���2���u7�|sK��:X����%�'��Ի5p��Z�S�8O�}'�ouF�/m�6���'�ߧi���kJ���6���N(���O{n<{&}՛x֛w>B���?���xK���U?>5�������h9/�U1��ZX�B���VUy�۟yv�S>��X�;���:�$^kw�W<�
�~�C����H�����CSS��^��v)�6}��E�οNV�Bxz���������3������CF}�
Ane�U��Ÿ=I�YĈ��Y�t���X@,�P�E����!5?��{�Vv������ɹ˱����t�;w���WY����M�mM���7'؞���tI�b�S�֐�w�Y�N�����茻��8an���Q��]���&s�,�t�o%�<
�I��n&���u�,�[}w�!S�ȼ���N}�}^��ᔁ}�w���Ĕ�^�^���@+L��C�x)���X�m�+�`^��Ny;�"�'F���=�C�hw��gкW����rK-|������B�����X�;���/�)K�t���g�o5پ�^�K�i\����f=��d8���/����&��]
����L98�{h'�;�V�Λ���ÿk�*��\���R.}čj=��"��6��Z=s�V;��Ga�%}�7�U{��}^t��-��|=^�$X��*��*�`�����??	@ݐ�<9~���-�9�����h羙3W�b�N����{��zS����r�9� ,�'�m����Ɯ�>#�Z�ɩ�@����!W���5^�Q�Z���:\�fϭ�}i�ّ���J�ڼ��um�ta�x#�~�c�n"nXW���N��}�O��p���}�dQg*~�-���#nO*���g�����Tx���ǳ�v�����I�:v|?wٵ��:+N�Ôv���1YcdON�qN�A��oi���)m�IS%���hI��✞�@���� Uet��ֆ��}]�P�$̷�����`�9M�/Z=I���]������-��+p=*�:#�c�B.ձ��]���%W�KDb�j��ST//V��^�gѾ��_�<��H�Pf�}�bo�^۝1q��n$�v���y�#ʫ�{3����=5��|����_�$d{�M�/V��e!!�	��X't���]�Ǔ�>��>J��sfaY�V�u㮳s��5��_��k�x��վ)9�˼���zk�r�w$�ƕf��$����=7�F+�w��T�}��!3q<��Z�{K�K�}֪xǯ֠�������}|1.����U}2��*�޸xS>��O�"_�ǶJ�n�Y9�>7�7�|�-�+�"���Q���ZU,��d	F���;��SjyzM��e���m�����v+S��"����y��oG�������/=q�ϔ�f:�K�_�9\Uz�|wNQz�{���=�J}��p>=��Y
�篅?:aǐ��d{���~�dxdA[�ps��s���罽�����n��Q���^Ä�}��om�a:�6r#ޔ��6Z����R#��K�k�ڴ���:3����թ�E�{���j����U��ߎ}��{�zbd��B�e�X��ˉ%WWB<M�L��-+&��b���N�4�ZV�*ruks7kw��5.u�ԭ�v�"��KP%��5�t�vShaW��It�k���V�!CPO��S\s��4�cY��MIJj ����e��z�uɓ�UY�>�UD����/F���DM9�;��ӟ/M��n9sn��u���.�ܫ7�g���Rm)T{�rMC>%��0��R�nz�vV��wǷw�7��şn�Yq|�V}�b�n9�71o·�����9RM|�'�����q����2�b�F��a}?Xοog�r}�~qW������Nǲ3|�~ɡ\�D����I|w�:^��pj}ۺ���ݍl�'}]�=�/Ooz�3g[ T7~��^�-I�H��v$Z����f���YT�Һ��񣞙�t�Ǭ�����mV������� ����9:�7���r9�}j����������+�U��f~��q�Z�q�~�"����s�k�_��~&��P��=�ƿW�ǐb�8��O� s���S������ZgZ#0��`�\?g�i�����ʢ�>�K3�#;WwAھ��R���3��Do���;q�o��=���VQ)̓�T���{Ň�Y�b�����ŷ�˖'-ϫn�y��<>gF}μ�W��T�W��Y�lL�Q'ȩ�����OĪ�f=趋��Jӧ�(t�3)^1z�"F��fԏOuw]7�P�wL�� �,�{��୔�3���f�l��⽳#o_:�u/����k������n��1�ۖl�+i�����E��£[hh��%f��`-��Uq}�	=w�rW�Z�3����Oӑ�0�p]{����$i�����t��)���A��YysU]Q��
�������k��"p/�jo�q��M���	av}�4q���]���3k=b��x���A:3� 7(-jj�}��׭"H��s{x�'3�����x}����~����`�ۛ�,;S##����|N.��'�_�1�ŏ�p�lkP'�ų���=���s;Ģ�N��ۗ"��S��!��/;VE3�8��x=�T�˱�!~��eh(g���g�ؙU�/�+�:����ωD���St��u׉������W�L{���Q�ޕǳ�e����'E�~���K��9�tz�r�P�����;�8�;=�ݧ}7P��en�w��5}��m_��;�z�vYϼ�u�wc�ڒ�)��u���瞷]:��G�~K�9��20������?�P{�ͣ���̿^�,�48�:s<c��kv9�e���=���?}&��� ~�%%��ge���8\�t�l�'5K�@u?{1�o���3���Rú��(h���蟼*m'�-�J�UkM��ci���Y���A@��R]�{�����I�S����C�������nnT�k����r���:,�z��2�Ύ�$>a
1���+7��շv��/��A��2إ��׺�8+��k��I��~����Vt��{D�P۝�2�[��׈y��3�<�F����j��2}P��=��7�:�>���7�Wz��\,�Hv|����/�u��Mτϳ�y^\X�L�n'U�Ȇ��;#]{ċ�:�=Npo:���F`���ە1�@�+}˻Њ��}�Oz*�<kׅ��:ϲ+n�<R��ֽ~㨿w�c��YhhU�/m���rc}�Fʅ�.X��.H��&a��[�PT��?�_�ǲz��=ҙj;��*Őo�;4�#ՙ�Z;�=��z�¶��� J�<zn����L��BQ���#��ڕ��"7_��oo�v�8�|s���>�~rJ>@�٣�+�]
.Z'g7�~�O��4Y�׳}x�bY^#={օ_���AW3�'{-�;����,�l��10�}t��ݤ����1��+��_)�����M�ޟ�T�w�wkō�yS>�����>wpDש�@d@,k����j�{������oz;zQ0��{ON����7K�㼹���_7���������B@����	O��	O��$I,! BI��$I?�B@����	O�! BI�Є�	'�B$��H���	&�	KH�w$��! BI��$��! BI�B$��! BI�$I<H���
�2���P�-��������>�������үS&�)M]�y��SJ�h��n�M�K[FV�{�||𓞝ֶ��۸�v���w�@��-���զ���I^إJ�ڣ÷4��ۅ�o� �=+��݃A�7`�^��]�\�{��i\�h��r��v��{���e��v�n�����ս�RPm�9�-���ŚDx{�uKۻ)�kr{�     51��RI@d4 ���d E?!�*��� ��  F�JU(       �O��)R� 4     �	T�      %#@$� �B��zLMe6I��忏�uh
 �'Q�@ ����PP� U��  ����oġ���?��Ú1�Ed AꊫD�C��� E
�R��J@
DP 1�ݎ4��l���ϻ��UW:!{T�hJ$
�}�+Ƙ���ua��Œ�B�|f�w��߫#}�|V��ʲb��R-nR��`{L	gtAx���T�Y�� ѱ	��d�m�˙�C�@k�{A��A��ҙ!��(�l���9�����Yz��e,�m*3��(��c�쇪������c܅u�v#�LZ�h��%��+INͩ6d4����x�s.�5�ӦX�қ��B� �
��ai��H���蔴��
����N�4�V&X̼	�1慅#�5ސf��&7��$R�*�u�FA@΄BP�I�C���!J��^��r!*��9�� �)�2��#fmՁSh�@��gs�-�[L��6���*�wr
PJ(m��Q6���\VѳX�#$��4R�)Cgp��O"X�%�(E+L���ê`x��!��"Y��,��eJ͘v�ῌ��qR�ga6swN�#vJ�ZKŮ��#e+�L��I�ј��%��'>������W��HE����F�V��1��^]��Ȼ��U�L��76�J�<���R���)lv�,$ӈS��L�nK����_�T�n(�v�T�f�[���ⴛԉ�gH	J��P$�ܦ%ˆ��{��Z{��u���`R�;�d@��v�|	K���r)2�V`י�КX�"�U����*������Sa����n�.E���[�kI����^c���6��Y�0�Lt:b&tɶ���a��O�3cP�o6���Źh Tr��"4m�2U�ŷ#L���z�a���.��oRm��)W��L�N�� �bc�O(�f��� �]i̹1�Q�͡�d(��\����6�2-��܈�u)��Rb�t��5\Yb�l�¦d0i���h���-��Q�e,�^D�t��7��=qc�Fۃ�.��~�����RR�g��X3�S �Cf�S^� ���i`�a�>�����@���2b�.��\�[�Oqr�
2�.�ګ��2��b��PLNM
�c�omy�jc=��Iә0fS��AzZ�$Ol=��qд��B�vh�� b��g��E����y@!����$şw�{bO�qȻ6���}��[�a�f����1�-]H��떻�!��j��Ns��u�5:	��7�m��6ν�|�vh �=��f��;C�X�ī����{ �X�0�e��:��-��Ӆ"vY6��[f��|�	�
����jy�
������q���C�ޭdx���U�a�W0��zw)�̾��pƊ���rn˱��1w�ul|���ՊH,/�<��5��{���l��g8�
C�V$*=W9>U:��o Y�_ǵ,�녋��e���ʅJ�r<��_u�v��?�P"����s9b�.����7�R�ƹ���U������;�;�����-�� G�:���oq�g��.\)����-
�9��wi��ѧ<"��u}֊��
���4�3���nP�'`y�*�'�P��Փu��,-ćN� U�����K[W|���蔚���ن7z�����a��Һ�B�u���ʺ�`��pI˺0��Ļ Q�Ҝ���}��'wT�Jm���H���)M����'wwT�:����I$�K��_{ڡ�L[����>�>�PE�Iˁ���W��,�Rj�/�Ǽ�WV=����mI�Ȝ�宻|� �vM��g~�3�����<v��J�) 院>�ԩu�(^��m�5�%����[
������ټ��q�I��;-�w��ݶ�;�٨gU�ӟ4�q�ݲ���*iM[���Mv�#[���O����.�Vb:��-�l����R*
�9òxvʼ�z��	z��%X�����s�{�6����n�Y��EUWv�B��1�E@6努��s���,
��G2:��3Һ��#01dP��^ҫ�s6g�R�[�7����p̦~�&X6{a��{���թ]��t�&���u��� � ʝKd3jpl���JŦ{z�ʎa���g�����z���Z+^Ib����mvTx;��V��:�gyR)�:i�·ox.��F&6.�K9Z1�ru�޷��%p�6wIe�ι�ΪOp��U����Ŕ�Ψ�R��
�m�|իҭ�uN�L_��5�fj:O��t+��cka��(�3��<�N8/�}���a���Ͱఔ�R�Is5���mu�T�W��dx+p�0Y��ޔ!��'b������#��Ĭ�U;a،�Ǚ3�%�Y�o[��;���H��m��g9�`�}4b��wxwtbY�w{�.�yV��E��Ⱦ�m:�x���E��_ĭ��եv˽�}�4c�1Ծs��t�r�ۮ��Il�I|M�\��6X����
��擎�pp|�4F���y�����s�bN5���u���N����n�ts���U�FCK	Ӫɇ��LVX-f�.�uL������#�I��Aa�-u�gQG��:�I��
��S��:�;��ss[0!���4���JJ)�)�8�ь}خ��xN馺��f� 1�&�c�X�ӦQ&���8\�.�\��&�[�&���W�K�&+��w{pN��Q�{yGVHb���MgIS�*�}�+���w)@���	��n�z�L_�\�������Y�+�Y$%,�7�j�f��Syn`����%�߁��.O5*���"�Z�ۓ�T�r�0�cKd#J�,0)�P��Q8x��kh��D1��e�g;X�v�~��.�����sr,r�G���^�F䫡��M����WgoK�Ms8&���U�Kg�J1��t�@լ�ص���nTUX�	'��)!,�	�p������ĉ�~�M3�����YT��
P㻽��!�p�i6yvGպ�H����.���vf䌳�]A�]�� �~<�lt�2I��u��o-b�L��L���Q���"��Q�F��*z<O��A&��F#��$2
���(%EG	hY�K8A�@RH�#QY"��UB�B劀dqI���7TInDl��yӜ�ך�}!�5wm�U�@G~��p|]mJb���#({i˓q�֧~�N�,u�Ҋ�ʺ�>�7E�����8)�����QG��q��s��_ޢ������\����!Ö�g+�;���H_1e��5p6���v�ѱ1RK��ދ>�7[�+�ͳG]�xQ#�mn�<|+ً#��+ޕ/�T �rS�_e?;�k�{o.^���C� �S��=�_�*�rg��IZ��z9�͓Q�=����&hSo�X��d��$!6P7O�4��UJ#׳���ڠJ�zea7��T��S�**�ۖ�Mޟu㩣�b���"�B
�*���C�ouq��	�{��L��,-�zR�!�|o�κMV�g
��Yy�����ː�w���.-Y&��;��Q�$|[�����;��e������B�j�+	ւ��l/�[7>N��C���ΐxCY�~<r���Չ�{��n���tȐ\;i6qY�k��Z[�/k�lTw&z�7����a��@zH�ޞt��㓨;;���]���D5���F��r<b.[�������Z}�|��֘�5bwdi�ݗ�'ӽ;z�X�~Z��(b,�n��ȗb=B�lĜ��a��c/�W�p>�?[��	�y>�|P����^MM0��Y��������hN�t�%��g���L4tW5`��{���49Nl�v�ܕҳǆ/�aZ��%B
�J��O��Xz�T��Y��@�J7��Aʙʆ�,��]��=��Q��~����P&�䱾��� �й�c�HR���ú��>�*i�9p���w;�	]m��njS;[L4�E#v�i��ʑ`8c��9x�2N)�Bދ�m��rT.��d�>D�b��R��B�� ɊC2��,�Q�E��@,*�̶q��-jzkvr�x�zޥ��̠Eȫ5�w ��2H��,�>�syg���D���r��6�,U�eAb�D2��e!$AKZ%
� ��0:�6͚����X�A�3T�_]:� ŷ���/z*�q�A������k���;�2j&�z��\��-!�i~�D�2iX�h��Ua�g��vdl�����3,xW��<��v'��vA�m~v���'�S�f�������q�C�{�:�>*sd>ls���5�l
�qk��\/V�n�{G���(06I]dx�f�f"]�w������F��>gu;�yA�G�s(k���D�/�Х�c=F{�>�j�/.�G����Q�e���d��+0��g��lh���n�4��~�5[��_�oF����i|&�j�T�j
5�.p@�Y�\ub�T�%  �k��k�j�����1�=7�]�йRZf����y���� �k���bk�)�Uq 6ARAB�A�k|ee�CT3����ARE+B�JX����;"�����
�� ���L*Z-�.q@�(X�--	�/�Ȧ�)� q@TU���M�x:Z@��I�|���-{�9m3:(�3¯����a!m*��>���;k�뛳����w���9�������t?����e:w�X
-����uTU�.v߷��M�UqV�+� �Z�v:f�*��b���[qwZ4�����;��ʍ�UF6�a�4�4�T�n�	�DzQ}��<��5���֜^ê�z�k��&2���_��]u�j
������6����o����;�5-�QW�&�mڠ.�;U�B��0���^�Ӕ'��P\�c7����+��N�y�u̱O���?����͙}��K��w���6��<=�y�žAȃ��҉#�/�-��B��`}䏜�6�םv��ǀއa5ue�c$��2����w'B�V�<MM/����?-B��3̚�gQ�ju5�VJ�d�f!.�fP�i�5hH}�.ٍ\l�f����S3|Z�|�����-�;��+�J�'1��+�����uNd��_ob���iG������I3�h�4����W��'�:}p]v�1¤����-wl]�V�v�r�YVfE�VE�m,�0���}ѻ9��B7XF�[.Y�"��r���LRxr�2��1�B
���ͭEa�a�I�U��,bt��^�q�i;m���{��h���M����~�S������ Q@�K�%Q9l���AG�B��V��K��� %� �ր�Z(~&���)H$����e�h}s2o~@����¾��`O�ǳd�o��d�3�w�QI'{�q�;*�={k�an�w�]����<���Wr��.>��I`��k��p�P�{�����Y���X��~Ȟ4Q~5	ó�T��[)ěz�!�����
Nr���=.٣0\�E3m�axE����dj=�����S�sY��̜����j�-��x�Q#`_
W����j�$p�s5��Ks�;���b�՝� �U�����@��/pZ��վږ�eS6mL���K�<<�~��?W�I%��F|o������)����V$�M�&�n�9h_r�];�%��m�
����t��]R�7Y�[����M�=�x>�	���l��b^$�P�שޮeiWsgɵ��~~\햝�DPi*~Q�D������<���N�2���SF�Z|�So�#hݔ��g������g��J�ѱ4��5A��i������^8� �%��0c�}#J��5��rS��o.��it�U����Ȭ|N̚�q5�c#	w�=��alG6dƫ�>K�)�I��\t���Kؔ�}
��{̆��a+T�ϱu�˺m�[5���2Z^3ո<ZN�!�ui�!����<Ss6��\Z�1
�����4�KE�kI�M�2ϲT�۵��Е���=%'n��$��Q��bk&ۀ x�1��7K?
�͸�4��P
���!k�᷍B��5��M$�����+�^��!��dΧ)�3�_/�9+8�6��3tk]������.�J�Z�cLU1��K�kV�T�s�
�Z����Pl���)�l3�}���ϰ�9�,��۶z�U�~6�uۣ���X*Ǥ�VE���jycI�rwVQ����aǆ���g�\�>�1�ŵ�6�K����jԆL����ڵ?
�sa.�k���L;����"�j��X�=��i�������R@�I���0,���n��M�x6���H��t�����߰>��� �F�
���8$���X%D��B��BptL�0RF�b&@н�	j1Id�Q!�**T/�\�Ç<���r�_a� �B����:&{�4U��v>�p�Sx�4�O}}lU�
��7���*�oyG�61=�N��"Ѝ^���uf�����L72v��*.=��xpr(� ����\��wW/J��M�9��d��9y��4-�۰��: �7y�x}.��5)q�~���xc՟��������m��AV���_���y�8(����V`�i�*k��u���J���|`64l
��皽^����U�m�jIU�,���]��;�!���r���7D}C�}�g�_����&+�*�~=���-,ּ���L��c�g��8�Ս�̊A�����xЉ�Y� 3��l^��?�b��]b'R4������)������{��/f9^�3�d��s�h�n�g>8^��s��d��6���0p��������#��`K߿a��1�]e5.��5�eg�斜rj�D�����%���o�ɫ�6���'�:����x D�+Kz���q�٫�hSy[w~|����ɵÅ��|�+r�{(+�L��e%��-+^�q����w����uɉz
�2��Q���m��;t�fօ�����PF���C�?8�;�<��84G��0KD�ע��SWv��Ih���ٚ�5�&�/��.��Ń���]�/�����>�𳖼��NP���^����<��98�~��h��*Z5���������?E�"9�o��z*s�O>���N��K^�����A訝�jƵ����s���GP�r�Jb���{��%��4H�!r���	~|���ob���X46f��=:;}�~%">#� QQ���('��'�~�����K���͋�pn���|h�]��	(�ѭ���J�	|7��7��8�<�*'���[ظ&��F�����ҹ�����z.�%E>��^Eo��F��V�B��e�����0�&^1��sR���]�zI�ZWs 	��6����Yoy=}�/��4d�$2�	�Գ���Bƾe��b���Փ��R����V�`v�éi/���[ٽ%��um�0��jg1�r<����ܗ�Ɠٵ��!����V�K^i$���Ē�K!�X��a�:���V���V����Y�����`	oe�ʂK|���X��nWm���QZa��f@�EEd�H*���M6��V8�#v)�	3CD�1X��6��Ϟ��z���3y������(h�	�4_�;����Ӣ�pt@����#E�n���kèfE��_r>	�{�n	q	�y��D�/}�j�Z�A��z9�sb�c�@���sq����o<;������
��>5+P�Q{�c���n�ݗ�?%j���~�������,�ދ�:7s�@~�,�5�y*�ѹ�T�~[�~�a�׆	���LTT�bS#�WbPNo-0k��
�(,��N��ř�.	pM��h���4�����dG �:9զ���o�,�V����l!��<0p�ц Kp҂_�|Ή�Ž�y�ѯ�=�|�ܚ$�)�����E���,�ȸ-��.!�7���*%F����39<���h�>�t�ߦ/��9��ң��|�S���~�3�y�Ĝ̰׫mn�뙓{�K@� �AH�0�����~�lMz%�;ʸ'��4

���|4Zh�$�"F����=�5�E�T��?6toEE�%��/�[g24A�S��K���w�V����y�9�z'҉po�1;��2K��g�2x�ᤖi;�x��V�}�<X?���~z*|/��|�.��$X*Q����
�o��?\��b��w���D����h�M�j	~������x,\�yȒ�4]�K�w�k��65����ٌ�>4~~�S�h�x�w�!�'���lSq'>6��go;	oc.6�p��(K�q����|����\ �VE�ʒ	���\���b���gj�|�po�����+Z��AD�Ur>��z>j쉠$�"~��x.o
����D�G9��8{`n�(��M�����̦�R��x3�ϙ��ȰX�D��.��s��Ÿ��S�5�]e�U���	�����t�evl҂�O6��yѿra�� gQ6;���^f55$�	R� o�.���]�{��Ưq��9@#K�^$[�R�^��sP�dW���>��n�SϤ�5��Cn�c��W���(eg,���~#4��C?	Z���X>QR�y���;�e��w��+�E��������֎���^m��Vif���p/
����X��B\��79ˊ���X9ww�ν���]���z�Z���"��v�R+�1�`X�Ɠ@���	d��f'��Yw����y�����xZ�������X:뫪�)�65����|h�5���\��n��T`��'s89�{Muъ�p�O Ɗ�k�^څv�u�w�a_?��7����3W,}t"�/!��qr�s�4�pݏ�NV�z���`�4陲'�F�e��J���Y��sE$�*l�+*IE]��RY���:5��ub$�E�2�y*���w�}�L8-ܺ[�U�dT�lPJ7$Q	$I��	�PTrF`���@�$Q ���?���.w�<u�Q%}S�e�[&�Q�P���Z9�w:��S����S�ۘ �lOD�<�B��f3^
����������Z�]�]�;�w���ͦ'ǔ���;r4+�&�q�󺻶���ޤ�n7�=^�F�=uB!��h[�X��'*��켠
�Oh�����ʬ6����˥� ѷ.x�,G��H2��陋0���C�k�4�ȨS��*�vα���lk��"Ҋ6��#ʯ��y�����:�bX1gS�2�����+�Ea��9u��z,ҝ:�vp/޹����0��Ў��c�ϸ�+x���vk
�+��k�������O����U��0<:���X^O����e"ѯ޷�,�G����,#���ۯ�>��l;H/Np.�'�"�q3��G�7���jM.��lW1;$t��u�%u%���z��ZS[�u��Y�:���QZ
�:9q�yL������f�si�vLǛ�<�u4	�ܯ:D៾�z/K��!�����C�L�J�4�O���-���(Q�L���޶�@a��jq�qb�%��ff6t�~�eoa�0.�S��ޓ��@lu��}�%�:SУ�uE��U�y����Ej]������^J�e4࣬�ö����&T�4+g��9��6�^{{�ً�d�W���_L��X�Pw�|�od�hj�6�5n�#�̙������Nn�䏳�� �v���C9�����I���W�|W�쑭k�i!g�7�w�
���郲��Hpl�/<������� 񷃍���r1�����^��r_����v��µOV�8l���s�G���CXu�Ӛ�8%f���G˭ef𕤙L�yl�DvU��v)Z��#SM:λ�n>'��;�e;7���I��'ȶ�R��Jި��P��-��e,H�n]:�ʰK'���6�K�z����1
&��D����Xm�˕k!h�l�l���cV����Jx2���kB��������/,VUBȨ�A\��[d�F��b3r���Y0[`!i6%FXlU�r@A�I��%X]w�fo5�[7Fq�*��C�O��x>����(���0�r.m�OM�~�n�����k6���I`Y�� u�:';�>����}Gl�Z����z��<� �r��V�S�[u��&��np�	�l�A� �Mf�����z+ā���<!�OD��ꬪ�{EDT,�������0��þ�&y�G�=�K�~��3��d�@���ݟ����M�TX���f�VN�*��`��.5MK�������z����M�S�����F���]q9s�&��co��뼙ż��H4-�a�gesC��y�Ҫ^�� �9�[�gn%��}]^���փt�{�-�[z`��_n�4BJW|}�'�fg`�e��v��G�`�8��m�\3n�ܼc����]D3��J����B����+���w^A1� ��3r�P�eI�E/��Ӎo�uF��%�{��юʟ&m�E����b��Ʋl�N��o�_Os�c�˝]�t��#״h�xX�	�f��O��x�"�.����5Q�����y�y�iR1��m�o#���B9
���]���U-CG/eѧ=�l�YO;��^�N  �K��D�M�{�薏]t�p��Or����`0��{]��5X3|ˎd�c�E��X�@oo�:�Ip��.�9mMeN�p���|bB�u��;�V������%�U�T\�^�I����K��t�{�b L<!n^�K�����lh�3xM��f.ҁ�r�$���Y ��]'6��m9��Y/VU�荡c�V��ZTl�����Rv�����b�7��[����_k����$l4���*�)�j��b���f+���L�X�m�jF�Gy� �1t-��mX�8]������a�k�7,�N�,V�4w]��~�u_A����*��s"�D��e�� ���r�S& ��"�iF���ce� �
**V4�$Yc�n	h��T �o1oOX�'%g��﷕�3L��ӱW���'=��������mZ��������`y-�ZL��	h���S3�ʶ���M�K����$��n��0����O��.�)��Q�L�ۣ1Mg���9�;=����w+2Wd���Ф�%��7��i�s��1F����c�M���^�1�~�W�X��K���d�H��^×M>j��Y���
���r�1�2�����h�a�3��ٸ�KDxa�B�6�Կ��_~�Z'��~���_�"������׏ѭ�[Ͻ��������e�=�'�=�3��M�ג��p���@o��YwCn�B{�Y9k��x��������<��ËD�F��k�8��_p4�y_��1�>T�Ls$-��F/����U��D�U�y���!��_ ��3FY7P79���O�utq0��`l�qco� �L�;sVt�n�}柱���f5w+�#׳�F�M�fL���9)�ĥǤ3���?>j)j����Փ���^�0� E��ۈ��GL���*Kd�J��2x�M	��R��Cw��&�����L�!�G�s.������Ͻ =�-%B{���<�QjtU��o���L�Oo���NUy���礩���c�ii��Fd$��E�{y8J&�u?q�W���:��a༿\�TE��-`��f�|�kt�5���Ɖ����^^ђ���kR������º��!Nfy�.�ù�"{��X�@ЀjZu�5pZ"Ɂ�W�+��f-p=��yb/nP梍k�q�;�+kz�졲�^��F�]��E}��G�HΦ
��!�x���ɋ2�9(#}x�S1b�@���4�f���+7z���M�����x��;x]�N�Z�:k��V�� B 2dK�e�n�ʦ�����$ �T��e�R�)l�(R�"�H)>#�?�BY��z�`�ݾ�T���uw���Ә��yOwpO]7�������l��6c�e�~�oK�^�A7<���=ަ\��w��3jo_������3��W&u!r�M�H�qO:���K|��E�F&��;�X(U��%�U1��p�D#i��_���o�W��K��v~�gi�����Z�4T����a���zF{�Z�'�fc��L�Rzmq�h��lW=zdi�+}M�'r��}�C{�?r9�_W]���1�"u�+y���O�%#�2���	{$�w����ĥ�3!u6Y���.μ;���(���ukE�ۏ�.�����P�T��&_?_(������+��_d�"*�u��^�(�������CU�/k�hKS���J��&���|��/�5�n��o���|R�A|��۬�f�l��^���<��J�F�#輽*�K�LE�T�x.��y�Kf,�u�/��Dt�)�\���	����N�=��ͭ�He���V�~Ǩk��#�~n�ew����|�w�N��>���F��v��w�C2�����|/�5�.��SeHi��SEX6���*�g=��)����M�D-�������oW�:��X��*R
������N�4�>0��o&͖V�_�N��&:#���������Wf�yK�Y%�=���ܣkrv�߫r��b���=�v>�� �x��+�~�%��@D=/3oP�Knb*O5[v���KjykI3���K�*{w0�'������[g��*V�y@m��b�]bhj�L����.*�3,K)@*9LѪ����ԫ%?^V��]���ڻ]�sʒ�iX��:�m���1����ۭ����wy�p�}5c3�Eh�+/{{[��B
^o��1뾹������I�{xK���ץ�=��G�[y�V_'�;��o�w'�p�]�$�<sy������.����e���
J��
e����R�%�PˈXB
J�pX�Y�2l�m%�Kl�c�R��)VErH�""�M ��������6� �J.��8�;}�����k���<I:B��G�Rд���w���on�{��%zǵ��\y*�s�X��ls��T�g�ѕ�u�dJ��S6�泌����EN�/�6�N�����b
��!jY�Ͷ�
�R��)e�̲�n�u,�������w�¥�:��d����`\���O���ס�^��^*:���Q���g�{
�y�W�x������{tU�C7�b���Nv*]�\� �[�H7k���v��s�&�H2@������*E�%`ח�{��U���.��C��;�0�X���?o�\:���Zd_v䍹���Ю��&m��|��|x;��=m�:�؉MeU���f@��o��s�U�b��ӦN��xr����mpX��S=��e�PWx8��f��s��<�%
�����S�8�q�x��r��>�U�l!C5l]���!��աNmR�a�Y{��r㾃�����>u�|��R~R��V�D-�1k�>��ˀT<U2pK6Ԋ����U^ʂD7���~ޗ3=�7&���d�{�w�����]�� w�\��5�GU�r!%�-���:����1��М�
�Ey�eé�0�t��B��#G���ӯ���	]�W���龋.'��ᵦ#""�f�P�H�C�,�=�9��2��ͫ�4hH����Jx�Q��E��gJ��d���__�B&���I�B�]*-FTM;pQ�-tw,Pepp����=;7��y�0����������o�P�qB   =)J ���(t� UW��Z�U�-C�BL����F����LS��c����:����A ����/�����P%�Pv$��(��a��U�A)���7ŬTU_AM�(��M�:q��}���t5�ҒT�^�+��H�;.G�fQ2�R�f��ZIL�.	A%J��۹_.�3�U~���z�{m��'�R.@sEU_�`D ��	�S���Kx* �b~�пK�?}�3���_��.f��(vx���g�e>u�q$ ]jy�Q[�Hᡏ�����-5/���)�Z�Jv�
@��'|W{ā��[�C�+Ј}g�LUY��\Kj�+�Vz�ʀv@E�zad�����DWB�J6�(�*T��]�%�n���U]��q	����y�Ⱦ���P���HB{�Q�7�'#p���Y��y���C��>��i�0�����F�*�~�@�FTN!�Cv9��}��S�T7�J��(!wm<:��uwa%ǂ�a�4�6�ا��I����F󢢪�N�$	�/2��=fˎy��2���4x_9��A ��w ���>�fB��҄��P-��
Y|�Q�t����yª  `0��$`��I�����d(�-�w ��NA���j+�ְ�i)I2��Z��<��iA�d�lʦU��
��j���Ϭ��VX�9����v�:�?C��?i������S�nQ^���j�O4 T��<�ޚH�)���W��lrK}�iEEU�;��p�	=KJT�����OEU��.�	�S�>��GC�O^�ܻ
���ѭp\r`aH=�*�T+;(t� ����= \�@u=<}>�:�A�X[�6��۪*�9��!��Ҽ�����0����!��x�@�(e׊q̸D�z����.�,EU_�`������s������{�Wf�UU���w�L�����`/v`(�dB�W©�Z��B���@N�l@Ӄ���ܑN$1ᡀ