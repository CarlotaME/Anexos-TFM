BZh91AY&SY��r� _�Pyc���߰����`�_|�>��� ��PP���h��&�	$�2�I��@MM4�چ��j��?~T�SF�      T��*J��Q�4��@   O?URh  h@    %jg�0���G�� ѡ���QE1MM�?T��i�z��=F� ��脑���Ba" �H|~�	#�t!��xr�;�M,���,�[$�#H�Ͻ�J�SC ."�Y
͖E������s���	�� �JJ @ 	(  @% ��  R@R@��($  $�D�J  R@$$ ��RB�  M����[�0�ŝ�zB�����+A�O«�0~&o�ˢSn�X�59d� K�ʘ���9䟈o	�7�64�R%b�R�l��(����Y���9��9�;��Cr��ͭ4�d�Ne���0kM�*�ce��LW��[/n6���,⭂���Af�#6v�T��jqx��b[
\��cF���uc�]N���"�SZw���ty_�χˏ�߉�w��@D��<q�L�I�,VXWi��
����$�M,�D��I�>�ݴ���j���,��V�WJҪ�YUUUaʮ\*�U�U�̪��mUr��W
�UmUt��������aWKL��*��*��ZUWJګ�W*���aUUXUUaa�iU]����*��
��[Up��eUTYUW4ZcՀ��ɐ�7�~�_1&��UYc�=�R��p*T�>�oy_/vwo6�m�    wdv�b�L�C��N�t��TW<��v����1F�s�jT�R&��l#q
]ƤU�6
9uv��Y�n|��jVf�ܕ4��h���j��Jt��{:c��緞<�~�N���ok�w���j�F9�=���sf�q�U@YUU� �1�0ɿn7�ѩ����Sۆ�*c������LGI�mM�tM��[}����C�u.ˤ���_��J���v��T;׵Ț��w絀��b0��뚛� h0E^O	�; c�y4�)ɥ�Ŏ��1�Znb�^W^ݣ�h��r���t�c5Ӟ뉺��odV�3�҃����   � <�#x��Ȏ�Ìw�΋�w�.q'�j��x��f���@6��bz�m�ʉ5��a������`@�+��򲰸�s`8�S�,��}��	�ώ���֔�r��%���v��ݶ����x<�:kw��z�
DF�&�=j��]�4k[8     m�y&mU��3	F�����X�P�DdL��ƶQ��%�VP�;`2_Q=��^�1 #������	z�l)̜������uc6�pU	7`d3Q==��T���V��S�d�^x<��}n��w����F�f�$�s����J      *�9��[WKAѐ'�9��l�Z���(ZFV;*�dfP
0���w@#S	���:wH����B�w2�*n�U��<�&�Ƣ�<�Q��Ei���&�F��4�Q[�.2�Z\�.��5�.���F�Hs�Y�ow�_5��Fg2f1u�L�wY�8�      ��3���z�������87g5�����`@�B���v�=�Jon*;r����ܝR,Sيbh�='y�e���^F!@[����V��Ǝ1{tQD�SS���V��>��������C��,���z�2������m���    ��щ΢�Ȯ]T��ʹ���$�t4E�'2B}+��޴�پ���wRہ�\M��O3r:���'�{{�%Sk�ԙ���N$��@H4DtW�g� �T�X�0�
St����Gl:�9�c�m�ȕv���oX�3]Fx�\��     6������OneFA���#��ʊg%���"aۭ-;@=;�l�K�h�Ȭ Fu�ݚ���)���S�O"o���3 n��*7�:n e�� :H����
�۔����譬h
���v����s7I�����8��L�wk��     6j�#Z/;/�� �oU ��������TI��&����ب'Kʞ}Yp�K�)��R�����`^9<wX+d�^OR$���3~=]~	U+2sl�}���y�nj�Ԁ�;3�K����Ѻ�y�f�l�.��M8  @    �,C����q\��o����zGZ�H���6�^oFZ=d�p&6��'��7�1Ci����*cR�Ÿru�莓�{��W��������J	�6.b������f�>?���)$��!�#�<tK�m-���n���ιewh��$4��JR��z`���)JX�vFe)J���)JR��)K��M�5����)JX���,R��FJR�)b�JR�)T�,\TbR���R�)e,R��E,�JR��)e-,���K)b����JR�X)�"�)b���YJR�)J���C�R���Մ�SK=���X�� -[+��$���������y��ۉ�a�����í��n�,�m��w8�����tK��0�.��wvvj}[��YmZ�'�q�fתcM9�B�B�Ǯ����"wF]G�<�'U:L�mE9(7��;�s��Q��T3�������C��,Vu��z��UZ0�����0�m���ũ@��_���i�̭��X�0>�K�����P†fb
1�B��z[Cdk~)��f"�R0#T�����&Ʈ��0�W���[9os���Srlϡ��/���?T��&��	���6O�<Lt9���=9�4���9�8q�H�����HqBCլ��}��XQxfD�W�Kw�E9`D4�|�L�L]��7::ڹ`qi<��f��5r�7�D�* �u��J�l.�Ƭ�I�)j���V�wI6�V1cS��$��o�%���I<���	�b������;'7�ɇQǄ�߾�C��ì��}���TR��#{�o��d5:9���rn�`f�[I2��bp�Ι�K���uy�}�E�dBA��=MY�n3���4$H����n�º�W��S)�Y�j��C�<]�*��[5�G�Ȳ�dd�y�&$V�AlK��p��ᄙ���t�w�'�Կ�.�p�!'���