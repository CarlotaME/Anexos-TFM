BZh91AY&SY�i%��_�`xg���&�����   bC��           ������ƫL�(���m�����n��t;fN�kU�uSU�N�wa-Қ��kN����]Ӝ�mҴ���K������n`
   n��o[+�q]��U��vukU.�m��W]١b��������1�m�횑�[lkl��gf��Il�)�sRv�5� �	4h֙6���J!5�m�]E�m�t�lڴ=�;^;qYm�kT�z���bʭ����s�k6ʖjq��c4TͶg�5h�丬�g�)y*�ۼ7�ƽ�6Ƴ�IGFum��C����fJ-݀ �   &�_v��[�.�[;,�]t��=��m�ïLK�[*�dMP�u��U]�٩L�wu]����lc�]�v����Az�Gw\Ġ��h6��y��|   =��QA@�ӆ�F����pP�:��PU 7�tS�!��'�=
�iz<(�@v���t�(ouo<:���x� ����UM5Jl���v���6-_   ��.�h n�x���W=�������W�{ԗ�+@f��ޔ��QWE���ۣy�UR�C��k��".�ϳy���<��}��;��[SZkn��ڮ��  �s���k˷�����vx� P�Ϗ�ݏ��3���� �F޵��P����Sѐ�7��y��z�)�]��A�=�5Ej�Q�T�븪i����F�u� � =�>�t  <w��v��]��7q�
��wl��M�-����T�������8;�m� �\�n���;c�t������b�k"eh�P��ڻ:�  ݹ�j��;�֥=�3�㭱�;���zt���}�
}����뽝*����<
R�y;�t+l�,��W�h���7������[7Z�ڶ�;�B�͖ٟ  Gw���Q��� t6�p t��@��Tp uWvn  7Wp �hj�;}�  s�\  ��5VV�q�ݹڔn�Վ�Z� >R�+����k�ڻu���Q�h7U�B2�BÝ i�x=�e` v�P: ��%lj��ѥ�{�]V�Mo� wX  nFg��= 9�n�!�8 q���� (��� �1àt��w� �/F=����Μu�e��K�  ��4�4z u9��F��� Z�� \�v� ]]�  �Ը: !��[���P |          ��R�Bd2h�43A	��F"��������@E?!)UM�0   A�  ��
J*�    �@ T��AT� �#@  Ѧ� 
H2�Bh����d��M�6���j4d~wޯ��a�P{��}�z�>�w;��{�[��K6os9�p<��<p����y�"
������@|US�P������
���O�?����������������������_�d�UU~P� _�DQz�V���������?s'����l퍲m�l�m�m�glcl�`�`���gld�&���񍳶2m�l&6�M�m���6Ϭ흱�v���&�v��&l�a�;`�&���	�M2m����l�e:d���D��al�m���� �"el����d]���6����`Cl��6��T��`l��T6�&� �(�=ev�&0��6�;a]���T6���E� �`Cl��Q6Ȇ��ۂ�Q�"0��Wl m�v»aCl����&U�(al�D6ʎ�P�
�vʻd]�����E6��P��Ȼdlm�M�������
��� �
����!�*m�����"el��U��v��l m��� a�.�l m�}dl"����U� �v��� �v�&� ��vȆ�@� ;d �
�`l��U�(a]�.��
e]���Q�"����v� � dSl��m�v��Q�"�.�l+��"�����6ºe���l�@6��@���`\a]���Gl�m�M�)�E�(�M�0��l m��.�l��U�*�v��@�eCl�� 6�;a_l�m�M���6����vȻ`C�T6��P� �e]���@� ��D1����� ���6¦�U�"a]��l��U� dCl N������ ��d �*`]���Wl��Q�
��.�l�*m�v»d�!�v�����A�
�6»e^�]�)�E�"��;e��l�m�M�	��m�fU�*��.�P� d]��Wl�m��6��Q� �`l+�@6�ea]��Dv��Wl�� 6�;e���D�+��"�v�;e]����vȆ� �"�v0��D�&�T6¡�E��m���;alm��P�
;al m�v�;eSlm���2��Wl��&�6�m�l�v��6��v��M��v��cl흲흰m�����;gl�`�;gl흳�cl���;glc�6��1ۆ��cl�Y���cl흱�6�0�`6ɶM��v��6ö��M�m�loY�0�a�!�CN�Sl.�O6���N��L�lgl�gl흳���N��m��m��`�;gl흷��q�l�e���v��6��靱�v���&��6��4öM��v���gl흳�v���;`��d�cl�lm���6���m�l���l�3�6���;clm���v��`�`��6��gl�Ӂ�6���;g�v���;e��6ǭ�L`�gl;cl퍰z��6ɶ�m���6޳�q�����v��v��n�m��.��`�cl흲m�l����d6�v�a�6ɶv��6��_��gLc�����~��<��c?S|~������.�ſi��82+j��Vd���$��[Y*̷kz*y*���o#��UwV%��Wl���5������]>:�4	�T��y��ddL��fvnj?&r�!�j�'iiUw����.�sf.9u0�r���Yduא��>���EřE[�ѾEeDg���͚��� ���:�6YN��;��mD�5��-W�WU;F�3F��&R)+D��U��8��`�Z����x7һKGL�X�;��$�̟J���S=�#O�D���)3`Dt�V��"�H��w��+'`�],]ԭCɚwL0�tR�{uǙK��;�k]�Mm�w�eW#u��F��Jc#�����Om�N�%R��ނ��"�W�2D�+e��:���[R�u0�V��2�1�>@b�{KeN�5M [��W)��Q�����[�^E��,e�LLC�72XU��f���t��tΡX�J�u3Wk��%PI#i�&Zΰ��e�f�.:
�'YٛPe쭑��<2+[dd��J6����B��v�!Zm�su�4��l���:��;ږ*#i���C���M�Rp�j�{Q���o�м��/��;��ڕ�#�Ue����ͮ�Cȴ�c�V��{�	H�M�ܺ��%��ĝ&�%VǤ5�3kW�inR�%	E;sFe�Db���*ǚ�Y);7ۖʞEV�Si���hkZ�Mn���d`�΋��v�#��kcK�w6+�̸	�*Q�,��pUz��r'.�Ձ�ԁ��]=�n�gB�cr�	KÔ�L��z �a�q�m�zڕ^�Ǖ�)'3���u�h�XD�`�h�_m��rw��=�3AB�"�E�J⌗y��VZa��j���*WV������{Wz��v�ٛ�����6n�-�a����ֺ֦)���pr	m�YVI����9�J\�(�(�"d&p֛a�pnҫ�X��Ka�X��vg0�EK�Ô*+��7I̺8\�lKf��G�YwP�Ja�I�e��]�pS��R��
��:�fԦ[�fV�B��Z���}��VS�yv�h3��`��i(�$6*(�P�{`֒+^8F᜷��j��ޝf�5�eg2�&�t�No���B�w��h<D�0�c�%��pc��5�v+l���0``�gg#�+,_Sd���N�O���K��N�f9c�0���c�b)��1�HV�f;捊��k�a`�2<�P�]�&n,�~ئ�{1,?mf�.�u�kH�W��N�r��.�3u;n`7,����@fM�iZuïh��U�mde����`�!V!Y�ȋ�}g{V��R�̸�0�`�bHFt���̡�F�AӻP)%GV����|r�l!�"l��%ft�JXV�B<�'DxUР�Ъ��+½�f>;�=��V
|o��FI��I�T�L�WI��f[arf�Nb�Ɯ�9��ҍav��WS�=�T֡�L�����w��{��Q?&{n�Z��v�,^6i܁=�;��9��Uا�I�4w32O*�1����+zA��U��IbPf�Ř��nF�Zj#��$�*��Gr���d�����b�za���Δ�.T

�� ��i�e���$�Y�2k ���6��������;f��_���I����(��f��b��$5��
���G�s�Phj���]��ef�!S]�V�	��ঊ���
e.�y�M�׳6=ڰ���B�F�F�Z�1�^��]ɷ4�s��X��4$�W�-�N8�7PRJ�F��N��ݬ�E0Ff1x����
���ne�lZ�E���{�솃v�歧�<�v۵�cIV;cx�]d���B�o�n�&�*�µ VS�=������2ҳ`�G�ܖ����`U����q�;-Y5zT��2��6�h8Wk��hz��Y��3�� �V�hSt��{�KDx���G���m� �wϬ-:�۰X5���fw�	�p��{�*�
e3�k�Q����6�d�Gf��IAO%Gj�Uu�l��E����T���/.��h�ȏ�S��O��kfK��J]#	h�<�|Jݶ���=���F*۷��fՍ�?�`���x����"��Nހ�ѧ+Ve��e����R4-��%�rhyD�L��v�["���	TR�l�"��*�foڛ�q�H�7dOc�L[y�r��M�ܖ�c��#={�����r�y��4��H��1� iU�;)f޽X/B׷���q�v*�8P���'��2�n���D�%��:S�$#S7&;�v1�SuM�DF�.`��x3��Vۆ3Q�Z�Zl�U�:ޛ��)��S�����H�]2�:���{�C^oU�<�in�k{#�uY�72�����-�`b����0աK�r�΂��XA��9n�#�>�����9%h���7f=���l&�;xN�2[:�L�����潒��W��P(�YxKʬ���N��{.'��������R7����{x����@�J�H���ʭbԝ;��4m����zb��yCd�7����L܊K�2(��d���ˆ�R ��X��W���ZB+]h������8���+���Y��F���+L=QǢ*�TR��Nbb��8�:�2U�*!H��vt��̥G5WS꾦ȥkv�y�ArM�g���H;����b텱��*�9��(<�NW&���z��*�����g�廥�]w7F�x�R�A!q�~^ۑ�G�2A4��y+ݕm`�j)A�k�,ee�4�q��t�����6�L�N(Hm:s5+��ĺ�76�-V�N�:Qm�Y��K�xZkF��Y˸�+�dˉ���<��m^aPbK��8�V`ɨᑴh���ҡ[�3V�-�"w#3+*P-��׸n��";��J�4	M����gu;J�p�۸���}�V�̫S���|�	��y$�f�Z�me��r�d[X�q���m)F^��aK!��c:�ZD�?��`|���n�U#)ѓq�%"�E��d�"�ڣt��m����PW�W����yz�R��In��Q�wh9t��A�B&��#�I��!l<j�޵X�6�[��f��DǗH���&<�N�7/`4���	8���Ǵ������ku�{�T�,֪``�c���[����l�_U�dC
V��J
�Ӭ�/�vЮ�
��3�[݊Jݴz�	Y�A�F(�A
s.�r+��nn��][��9�+kv�V�Ҍ�,wN���kMM�Q��R��v2dBe-�Bo7p�C��أ�U�Z�ۤ����*
<�,�u-����$h�9F�AXjU좘zp@�L�y3(��2��2tx�Yϭ��v�;�.d�y��]�v���G'���Y���^��mj)f%�ʭ婴u�W��)u��ZE!�T��1�03L�LQ�(t,ix�w�`�J�ʽ@����;)치�
P�p�n�yЪ��C�4+���rӹ��C-W3[ ��&�RlV�6S'z��QM2�[���Y̧v)��Qܼ�d�C��,���G�� ��Pw��n���7���ٛF�&��V�mR\�����h|u0������:(�7IV'��c��+2
Q�C1�XL}y�1,7�V�n]�7@wL<T�Q�܄��1b�6�#�/0��YI��+M���ƾ�Z��L�I��yb�lI�rV�(5�+��Nf�"`�蛘4:��h��7�f��Y�:�I4�5�l����܉��m�f;ͭ�n��ðN)LB�����ք�)�G%l{R����2T�T���JU�*ͭ#%�xf�F�I� �NTD�c��զQ�݆"n�ܬ�rf�W�J��V*�V�A�s[����T���K7aʎ։t+&�g\���Gtԡ�NЏ5mlmn�cU��h'N�m�@���R�U�"3! ��P%��
�XZ³r��)�oa�p��j��eP�w�k�]��Ҩ|���Ji��w���lb̬Z�v�+�@F0��|7e��n�w�9�5cu�5��u��b#Y����p��&�Ɔ�K��.��"��!L��ݻ��׹���\�M8S�'kt��2v��T���z�;y�vI+^Ң֝ǔ�v��C{t�e��k(+-�6�qk�O#*�R&�Lj�yVobi�F��h�(eW�u���	�CAf��JVи^��K��O���Y�-�ћfL�NȢ�X��%@�۱:��a��[B����v�*�5��h��I��{v�+�0��)Z�c�vc��P�Y�ȎIH�N���jۻ��r�L��6᪗�˄�at��;��7q�B��F�W�n�0�{V9�޲vł��.��t�.)�L��7ZHlf����a�-�ä�wF�分����FmJ˗1��B�w��Xa{�4+��&�:Z�/(T�6��Z-�m�=y-��"ݬha-K�:���蔻�u�^R6� ���~����ΥBZ��U��e5����(��:����7r��OU��6Z�BΪY)��`�$�M
�u��$m�Ul)Z������oݎV�mc���ZΓ�,*a�Zl��o�w����LbA�H��I��Yz�KUĽ��7��k�{~��G�M��՚���F���֩H�)�eA7�29W�M���Ȋ�Gl/��E����񢀫����+�
Q3K�l�i�©�%�.��!�Qg������	l�$ූ��Ɋ@U�A���Ͷ�S2]X�:9���3E^�h*�幄�cE���\�N��)�ݭ�f�ù��1]��%�����ہ���庘McܽI��L����u[65J�-0T"�A�2�/J�( �7E�r0pc]�2Zۼ9[��2�v�^�x�l֒�BX�^��3aUf�Э��)�t�ӂ�<T�{�	��}Ζ�������]����^��j���S4�j�od2M�Y'c�^l�VQ��Z�Wd��1XA� 7Yd[͇ye9�0b�+KҒK+;K]A�Y5��|3�V�u�l��]��Wp7�TW�-��*�f4�H*�w��sc��g2��B��nd���K�V�n�Z��w_�d�n�͡��?wD�tXx��t@���a:��0ǖ�4��r[�Phݺa�ȁV�-ǬC3ki����@�w����Ʊf�r%.�Z65��ێ#S�hF0�	�fi�bD�L��or����w��=�+bY�z�y-�9a�fkm�����ÈLi
��F迴(;-"����vC�p��	�uh�4
�X]V��|g��Z�FK��Z����ʓ�;C)�i>"b��s��7��6Yx~l��/jX�D7��C�'wN �y�X�WZ]����ԇ#o���0ubV��1���[ 諔>��4F�.�,;Z�[ ���M;�:�wu��]|&����j9��7u�ִ[SR�chg��KE֮��k��^㒕���JTB��!���-�z2����i�UU�X ��{-�k�[��P{�`��);ڳM��id�V��ۜ��Ζv�u{|�Z
W�)N�:Jl0�f<�����dztU�8_�b�YX��e�L�	\�����0��j��bk�v�i�-�S[��]9��݃*�f�`�s���i��Kv����)���@�Y=����X��WV��fa��.� 6�U��f��fam�E*닪�OQ��=�k��47&^����]��Pz��gDy�(�(+v�8��-saٵ�U���ն�.ʼBaA���b,�{�T�K2���
�F���Gj�T<h�;v�剈�C#"1���v�U��vR�����-��Q+���*�S\.rp&�H��\Y"��e.�JW�R�+�	"a"���P���Cw}����ypj��]�� ۂ9��������g|�(�
���"f!Vb�#��E���Z��uŷ����ys�ĸ�Sh�~����Tdl������f���8�[����[�.;��f��h��>���3��\�ỵ�41w^�B-K������A��>'�]�.e��1��7���H0��zZbp�5�K�
���&7�:�C�]ɯq��ͭ�47rN�Ҙ�8� z�� ��b�Za�A�Y��u��)l{Z�㭓�B�;�|\�}i�SQXDZf�Sv��^�;ըO4d,�E�뵁��p\�n�^��Ƀ������F�h�6�5�EٺW��XR*�gt�s�����  �w��������Qh��C!��H�}z�{V���\"�G��cS�4s��49���~����S$�|�b�`"2X���0�N�o�j1�+ԧ{&+0p�L2ʄ�1��t�ޑz�:��"g��&����V���-L|�M	�E���p�[Z8�*\��(ǥ>��&V�PhZe�Z�sO�"U��gR=+����ג�`�� 6F�nah�X ��Uz�Ø
��l\v���+�6��)y��_����d�� ߪ� �����}}썺���}�w��PA}1<��%�F�=ZMO�^���X�U�ឪ���&V"�@e�aH�9����3b��>) 8uo�ɝc�b7v��s/�	d��Cx�[���pD[7��M�s�`(m��G����G�q�f��=Y��&���!���2�	�c�^1�L�r-��bӸ� Yl��n�Y�z�2Y͢g�ݚϮ;Ը�#fK��>��
�_�SYos�C�,8�S(8)e��ޛ�yI|���s����ܲ;�P�X`�v�[�P����Ѩ]�}�ׅn\}0yO:`�Ո[�A��Id��	��D�Y�~�����ﲢ�K|UdVA�Z�[&sۥ������;K&Tn���˕/n�}�����dֽ��<����$�/�S��z�G�F~?��u�'�?���rI$�I$�I$�H�S��^f�'$��K�I$r��II$��$�ɣ*�C��X�r��U6
ε�-&pb��%ngLF��l��IRi+7�ݫ�Z|h N�͌��`t��F�Ձ��f�tj�lw�㫗�h@�7\q���R�t�|V�Sw]̏N��sܺJ[�^wy�L9>k��cU�Ӽ�O��2n�S\�cQ!�ܘ�-AIO�W�&���1^Ś�9�Ur|^���y�JD���<��v=�]4ܪ�U��ӓFߩ|v�׏��r��dm.3Cŷ-��	su�TX�n)��~��đ�����A����[c��Z���f,�� E`@d�1ݗ�͞����*^n�U��5$z`��.W�A��1��5��X���:.-T�w�$����D�ME����g�0�3���9`�V<jkZ\Zn���$QW��UdpS�x]T3��Z��K7oyо=�7�sy��-�<�(`OyY��|�S��y�ׇ	����E&ͥ�cQ�;�OG{�,�7h��5꯶oM��,�qh��d%s�}i�a��qK4��^�W�1��J����]�&~�4��ywh���`�ɋ!�r���v�h�t�*[Q��.A�gwnpt�A�^62>=@�_*�q�Y�	�/�j��Pr�Ah�tQy����7-h�Oh���F��S$��F_9ܺ��:�WWuw�J��{''�+�ܶw�"�"T���:�
|�5.��U��g�}K�X��E=wX��qG��*�~%�G�{��t������ֲ�
�5��tjck1�Z��0D�34<��ݍˀ����v�[���6r� ��=>�w�\�k�S����u+a�*g9m���E+��1:��ʒ���yul�m�^�����׼��B���}�	�\��W��"E<&�b�7�.�6'sG�i<r��զEC<�m����3���]��ʼA�[��!�n���-6�Vӎmhy�t��c��}�i�D֑�J�۱L�����g?t�<�ɾ'��yζlij�i5O���}m��C�"�X\�����'�P�4�ԥ�:��Vs9�pE��vK\	һMB�m]r�CHʂ�ѭ[��:sK
KpK[/u��]זA�輂����Q� RD�њݕ�ֲ+#�³��!���WΘ);���{�*ѷ�C��/o���䠉b�Q����m�=�A �3���X)��x ˛ד��E���*���V!�M'M�%X0d���1m�x��6��n��^d��0���$U�,:�@*����8�UVf�'blV��(�օ��ӯm'n��dq�W���u�ty�o[Yj�@M�sq+2mҾ�cގڎ�K��r���\�v�[̋ޣGk&�c����)Y}r��ȱ�m;t.�b�nS�4�o�J��;��Y���6�W��
�z^\�8��fP��3�x���Ĩ���*g	��j(��DԖf����Q�7F�0׏m]�{�'��"��|����<�wO�N-�Ets-���y����1�uC"��R�0�mm��Z��'J8��-�wA���"Tu� �H�t��֤��]ooCxݰ"�=m�pOn��K��݈�	x%W�l�<�����p��ozx7չ���4t�}������W]��Ca�}]�(&m��=z)!硏h���~!j>��X�Q� ��̳۳0�,�.��F�3��{�9�@o�_���w����
���0�����5��-D�Eo�eGp��wZ}C{hvh-���b�=o��i���\�P8v=������6��K�ބD�}��dk*�P�\I�3v��S�$Wu��7���i+�5N��Kkd�uе���RM&+�ٜ�[��j�5/��B�~�F��+V�<�vȏ�:��y�L�2f�l�ss[��cyř�U/r��k2c�%�e0k�)��9ػ���٠��N$%�S����*��iṾ��1�_�6.��Ⲗ�-����%٧� �r|q��ʔsS�2���A�3p��e��JU��N�Siڰwɣ���ڪ�[h����rnC����tr{��^��TDeԺ�3��n�	pɇ���k�I�g<[)博RF�E�9�L#�w������b�u����s�$kmr&%g�P�=Lm�����b���7����dsQ�.aQKo�Ub�.�u�Nټ�޺��a�n�.L�1��}]J�6�B�4�����m�������Y�K��K��!�Y�U7x-�Ȳ������<�r�b��b&9�j��y��6�ӯ5�+wW���v�4�E�(�]^`�eL�R%Y�k~Yr�Vظ�ٺ�v�W}К5�?%i)�;!a��܃漼��>�0K��������ɧ�W�o��I�2�vtKu�!���gSY�D�]�j�i��;��F4X���T�j����8��́����;w-M�]�����HB����bۚخ/��;oxD��h�As*A�7W�;Z���f�\�K9�oV?�I���=QDU�7R�Ӵ� �gm�s#��wZ�aΐ�I3���t���1aI�N�yŽx�-!}{ˍ��Û:6�wjKV�ɭ=I�]�hˢ�hC�%e,N��N�&7s]��K��D���7O%�BJ��Mb��%1�{�ӈ�5�Ѫ'M�w�<����ʃ'��3��[���i#��t��Ot��� ��ݒ��T0�s7e;�y�jq��!�����Y��"��L������6˸���u���ZO�c�8�36����c!WMaCQe��m:z���>�o��V��1v���6{Qi���r�'�6^i����1�wy'w\n�-`�|JB!�1�w.8ٕ��&�Ɖ��n��[nkT��:���6&��2츯w��#��eP�9jۮ�"d&`�=��ǹq;w���wu����Mk��
��FFg^�3S.�6u������Y�%3u�����\��k׈�ĬE�&mGz邚�[�D�GW	�m]hodޓo��;�0h������VD�WS�h�i�T�7��m��}���.����KH�`)/f%�٤��9m�'ι��{�X���Q���z6Wd�$��o-��T�J�Z�L�����3h�w.�19س��s4��q޾Qi�����x�eܦ��b���M�M��-"ս�hE�3&�{��q��ʽ1b�7W�Pc���̣m,�Oe,�,�S��q�E+��}�m0�˲)���b챖�w(�f]u�\�<�ӀVa���Xyys43\�Q����*+��'v�R܊�����MK��g�5A�l>�c:�1ŵ	̓�bq��QXB4mW����-�3�;���0u��ǴN+N���� ���J���=�חg1�ͷ��2[��|��ks����91WYy��6�c�:��L(@��7�n��
h`#���NJ+o��/m�i�]�63G/��f+�So:����^ѳ��ild���+o�$��J���W("�e0E2��)뗨k���(.��	V>��D�f&|�,vQU����nr���Wv�KS<D�h�I̑!���D��(.Խ�M�u(�*i�ykV�A�	����ə�M�F�
���5s�^q謷�Nn;�r^ю<�}��r���'\�:�m�t-^�aa�'.�3��\Qmm�6�Γ-���0v�?;m�	(97Mّ7���F�幜� o��zs�즱��m��Z.�݌�;t� C5�����2>����w��^֌�����a�E{LV���cJ�^�L�t�du��By��9�}�3;o��1�����!�l�%���>"�^�\�^"&f��nG����2�;.���W}� ӡky���F�I[g"�s��|����6����=Gm�9(�����8M^����T����;ю�)�pѹN^���Ae��5"}����v6Q螅Z@#_ �#��u�v��I����m���L!���:V�=��xZIU�|�|��#ɹ+���;&�|��Q�x�Y�­��w,�sǵ�j�#RFu�0�{���<�W¥-|�0wlX�x<��LyLe�5�ͣ�����C�5�^L�����'aV�����f�,�υK;5�b��v�L��F�t��ޡ���+4�������㩕n���iV�I�u�pȻa�P�m�[[A\�l��w��9v��+�pP��Ǜ��ɨrj�h}`c*I�e����Z���|��ba�Cjs�Kj�>G9U���3v��RK3���x�YR��J
��:���wnħp!2�M�7c��s)D�♼��Yٷ��FT8��,L�������^�h%�s�5�N�BF��I���D��4�)y]�s��Z
n�dzj�B��.�.�/%���G�����,ĈF�6�C#C�P]��cx��p��K�'dC�����'
B��4|2�ڏ���y�����N��)G�5&)ٍ���<��H���v��O���M�t�V��z��i����x,�]�U)�.K9��9w��P��-n��)t�g=c�k!gJ��vn&c���&�:Oo,(�������ڕy��E���a�)�\��T-��������MY�8^M�Lbκ�7��g�ъ|m���l�svT5�r����H�����M[����0i�F������w�Y¶Mu9���������M��!B�Z�Wfvh5w]ox6����j�#.�v{g�zd'B��n���%��q��Tf+��o���E���3mΕn��<1�*�@�tþU������d�Ǻ�����+�[ZsU�V�?e 3�W�sf
�T����XW)qG���[U-t��	�%���@J���{�Һ%.�Y�ɷ}ԌJ7�8iS(gn�׺6���i,�ͣU�ϫlnn�_n�[]�d
Rʧ��+*�PN=��w��"��ޘ�9S��8�Y[����tZuj�$TR�y����[����IH�y+C��r4��S�]�y��e*�c	u�A���YiP�*��6lEֲFzҩ�^�w;;�:M��]*�V��ueb)�[q����Iy}%X��F�q�{
&�5�MU�� b�GigS�Jt���z~n�-�rGx,"��iZJ��	9a��r7\���ٺ���(��;�h����nwzX<YZ�WaQ���ujv��;���,�j-����ͷn���Ο��N�U��o6�t�-]�ܦ�erd����,7ɶ�!���`H�1@��bQ�q�+In%�݈V���bJ5�X�h��5,�XF����hG	ӂ�J[6��g�{�V(���R�[�S����u�fY���Ú9}�p�������]FZ�EM�&M��Ǵ�8��ɗV"l�?2Mv��R�K�s��[C��.s㱣��; r<�O��L!���mX����g��:,���\�=�_hK__���j��2��a�,�@m#�$��+M��c`E0e)7OYpivE�ҳ#���3L��I���U8^>���)}�9m�m]��-.��l�{��ewp�Ԥ��u[�]B�FCMDHi��խ��0+�C�/�Dl�bjĴ���K�]���TqX��f��RV�MK���]4��&re�i�a�u�&�]K�q*G��bc��@_��5�c�>��1E��(S�Y���G��͛�+�:<w]s�wg+<��N�\=�
�*�T�F�5dޚ��oAo7w1�2zI�JXE�am�=�r��;=.У] t�;2�1d��č����Ō������e��"��r��]o 6����upA][6�x>��:���J�iC�/v��{���n%�8�6+�s�-�@6�C�7�X�7��K��W�Թ�RB0��\b���-�v�ZOeX��[��-��pd���	�:�J׺�][G�E��r��a��k���B�8E��ڊ��e^f���N̘ƈ����.Whn:���W�AkK��krE:$�\�9$�5J�I(�I$�6��҆?�����{կ5u�NYuo<�u�5�kwdn�x���c�{��1�hK������F#^���w�k��D9វ�R����nl��ϗ�G�n&7P�GY��#��btA��z�dw	�����O9��f>[�3;�u'^�� G�Z� 3�cM/Y�P亞u�{���+�Os�5Y���]�eN��B�`'�fF� b ��]J[��q+R{��]'e�쥓�/ l����zǅ�v�J�%0\�� 4�<|�/x���?���{���~ R�9X+� _0�� /5�߆����8��l��2˻��՗������r�_���s>H�r�b�E�s�5�n=���_d���Փ�Xx "���
�����>��E?�����~�@G�?����?�?��j���5��k[C~[�2]j��N�<y�HX�k��D�])vKHմ �7r�0��ϐ����lCv�E鎦uP�V;+L������P�r��
�X���W�����Q��N,u<��"�;¹�A*�������nf&�Iu����V99�ARs.��(�B�^�ǎ���m�W7�j�Z�5�!Z��o��X�
�� �P9t7;�*k�a¦��P�}
h��mm��n�S�4�Fŵ0�vِۋ���C����[F�'V��u_r��nkJT�8eY�G U��oaG���V����r���v��Y���܀�a�ͤ��+w˴��b�'�V��T7$�w�s2j���M�
5[�۹�]��7ٺ��HÍB�4M�G%숥�p%P!�2��Ѳ�V߉��j>�48�ƻ�4 ڣK���uk]c��wQ��gG�)��gOR�-P�M���e'��`:�C�����H^���Vy٨��Ȕ뮖�Js�SM�\L7#��l��ή��e�u�Bp��R`����ƠA� 2Čp�	��������S�r%�!�wr�lf374Г�F�Z�u�ݍc̅d(`��iUp�b��'��384�5����i�֎u�~��\�|3]>��}{g��N8�<x��Ǐ�x��ǧ�<x���Ǐ=�x���Ǐ<x���ǏO<x���Ǐ=<x��ǧ�<x���Ǐ�<l�W��\m��0Yk��j
2h�Φ�61^�N�w�s�'ۘ��Cj�w'd=���TK��=L�@�ƧV�l��{�aJ�����q9-�uƎ�ݷNb�0���5&���
K�1��vƤa	jY��=�+Ղmq6*r�T%j^\��-g&b�ќ��%�xȵ�X��$�њ�^�ݤM�B��pŵ�]�Je���������-�Z�$	�νv+������]�y���X��Μ�^$��J�t�a�֝:H���������K�Υ��3�N���,ӄ�ي ͍x{$bv5ы��	��0�Źa]l��e��K]��A��F%��Tå=���8�h�ٶ��f�Kv�Z!˥.� RJ�.匼��:��e9��1�;���ޞ��ר�ig>�Z��7m�Kb<��Q_v�ӄ�]&^����}`]��o�Ձu�c�z�ʷM9��0���͙]�2:L[��L+�	ڂ]2���a�T���z�{��x����oP
�!4w��z}�����ĳ�BҺ�_h�6���'m#�CYZ��[h&-�05G�97���E����3x��9]�1�l��yg��gQa��뮕�#��X�Ĕ�ك8����pO��E�g�ۇӗ�,<t	e�i1��y�����R�����I�	�UF��>�Oc��]:q�ǎ�<x���Ǐ<x���Ǐ�<x��Ǐ^<q�Ǐ<x����<x��Ǐ�<t��Ǐ=��}>�o����}>ߧ��J׶1i��p��o8ͥ8�f'�9�a��oqR�x��bʓH�N=�fA�R��ڎ����H����5f��NZ����₷Dw����#��:��P�:�4��Pyj0j���fq��r����5���Z�5�hLbt��+YB�h*!�
5v~�)X,�<#��"�m�2gY���W��z���:�is;B,붗�'lL#�Q^�C#)�ZۉgA-@oZg��6me4�=������U��]q���a�ح>�,"٠�y��n�K��81A�4��p���)NZ8��}�9��a߼�,{f��6UQ;�{l>�nR�(��̻�Z�뻨��i)�Ihj���꧚[����ܚ:����	j�vo�c�}_�0P�+2��P��9L�3�	+�i�ڬ��	L̓w���tS�↟mS�=O�6��t3J�{�o]E��֜�X�'˕\5��݀�� �z��#�Vw�UGj�;M���6U��F�k��R4s~��	#��9��Kh����bsm(5�aJ(�����݌��0)�7�M�ok6
�k�j^ �`㲘]��Y�w}�Q�8c%�=uYzwwJ�����������)���'pyE:o�1�o��ƿuN7��Y�m�s�T{�2�]	7��ϲ�gN5j���=� o�m�5ު��}��g���fX���7�<k��zrH7���w��-H���z��g�@F�k;%�1P��/�����|�ϱӧ�<x���ǏO<x���Ǐ:x��Ǐ<x��<x��Ǐ<v�<x��Ǐ�<t��Ǐ<x���}>�O����T�|�#�\F;�/p�3]4�!���fؓw��8*�Ef!w�o����h�Z�u���x� ��la���}36H�H��Յ/�b��W.�կO�|��t�r�b��*�Z����,Ja��폠��;�M�1��X����`<;�y!�aՊ���y�֪6�mc�@U�e��Ohϟxn4E�z-�u%jQ�4��@q�UגK�r��|hZ�2��rF�S�{$X��[��!J�ʠkFh�Y�s�
���=�N*�n��Q�;n�YvA��U�0�}�H�K�
5x
�Y\ �"�1�� ��i�y���﶑�t���%T#��c���s�έ|:�O�&k�Y%�D�!v�R oa@´:T���kgKM4�bڌ���CspT=���R��Z��y���v�m5S�v_:��0������H�:���
��]����kz�[yj�\_4G�Tl���&GGK��Fu	�*�6;��RZ��3�w*q�#�[u�U�T&�"+���P��L�k����NƗ(�Wс��'��XкH���x���m����e?�d�I��-��gh�I�����y��|��F)VLMv!�\1����W�9�4Ijp�4Լ�(�s�XR�QX2�w�=cJ����vn<r����3*m:b�k��Y\a�U���M�;Y�(GPU�M"��u[8(赕6<2Y/�ȁ���+]�?ot�|�:�{��t�����N�;x��Ǐ�<t��Ǐ<x���<x��Ǐ<<x��Ǐ<x<x��Ǐ<x��Ǐ<x�㷌��Ǐ<s��8y宸�γ�齝���V��K���H�9θnHr��,r��L��I4�3+��wq{6i�8N���+M��Ǌ��d�{�W�QU��@l�j���^C��\�<���+9v5�bŇjɤ����v�_	Q�oF˺U��j'�,�-�F7�52�+V�`��L��<���Q�雜a�ﺝH�NѮP�M\<7�i�`7�I�45�9i�P{|�r1���"���:��C�+]W4�5oEj��\s�LS�5�:rb�b8>&v'u�ps0�6���o3���F\IXn{(���x(v�!�e'�<֮�]�13g4�:�ٷ�Z�U�v8��C	6J(Mp$�w�|���#^���k�E
�%7N���t��@�_.a�uo�l�r���#�ܞ�9B�m鏪w�QKmޕ+�8wvu;�Ӄ,��)w�س8R���7@{���>�w!�'w�|)�U�)9*#����k�(��n�+���*��c6�s��撏;v��UUS�`�S����������E�wqI�ܒH:ͪr��O��uRA��܉qѴqd��z��5��=�M�Ɖ�׸�Rj�Qp6}��o>�3�&V!V�2��Z�2�:��^��З��ĞV �o������ۧN�<x��Ǐ^<q�Ǐ<x��ǃǏ<x��Ǐ3Ǐ<x�㷃Ǐ<x���o�Ǐ<x��Ǖ��}>�O���cJy��I�x�^f�R�Wek�{'�>�����ސC��p`꽴.�HGa��a�(�<̄��)���=R�ʵ<�@b���1Kkt�S��<���v��!����0=�.t+���7�V��nl���z����ރZ�'e�z%��U�U�78-��d���.���>���,��R�2tAN[tlYꈂ�[0�ds�X������sE�4�TT�#k�S��+yl�VỴbvN�ܺ�I뉘[�6>ǅ�*V��N�U�	fwB73Yz�g3�PU�C+-���v�'9���3�]�t��9u�V��m�]V'\��5��--��ꝚFo,�8�
��x좱��J���=ghI{�!������"T2��v՗(ê��o7W���kY�x�l�&<h�l86UU�^����4�<<;Z3��[�OS��������b�F��5�O�l��{p=g���1-n͓+��MW	�bӥ����A�MV^T5���pV�9���7��k�tƘ3	���w�1-�����w� ��
�����٭E���X�*|����W[��ާ�S�Cb�"�#yN��r�hSB
R�ڨr$�#��.��uaR���m�jޖf�Y:Y��c��H�'�'�gY�,;��ۧ�{x��N�<x��Ǐ;x�<x��Ǐ<<x��Ǐ<x�<x��Ǐ�x�<x��ǎ�<x��Ǐ<<x��ǿ7w�����8:�F��
a
���V��Ę���E4ۛ6��li�q��Ұ±�؊F���v�Kzf��#aB	{X1�uX�Vj��\]��1�y��f����\��GN3���V�\b���3xz9���S��1�L�8vcR�)��އO2w^�k0I��	�5�	+�ݫL�q�<d�o�+�Y��-��ىe�;��R��{}�z�^�$�0޳�ccv6�2�I2��|1nX5qn��gY6��
�[�H)m�sosOe�R�{@&>�9�Zʙ)���̥��~��&9�@���n	�S�3J�w̯VK���Y#��?-��u���
2��"��j����)J�cN����*ꂄ�*�1��qc��hĬ��8n�!S.��X��+C��N�.W�����[%�(2�U�l2�*K;]c�⋻�+�*����h#I=Է:�^<�x�*�[	R	d���X���JJ%�_qn�CmN�c�,�e\)�Z�mf�"6�Ɏ{�V�
!�mr�|;��#�QZ,�,F$0�9]YS�u6�C��]��<��^��4��-1 W\Vq�n#H��hwQI�M��:j���Θ����ޮ)�(�C�#!��\V���j����}�:�|�۷N�:x��Ǐ<x�x��Ǐ<x���x��Ǐ<v��ǎ�<x���Ǐ8��Ǐ<}x<x��Ǐ<x�_����}>�c��n�j����r�bz{״i���6���cq�Ku��5ٸyR��m��qJ:�w�y�K)V�c��eW����ɋ�N�G�noV,X��I4�Ga�/Cٮ�>�����|ܕ���kO��Uw���ϰǭ��ilO����grK3hgfܖ1+�k�u����q�g[� \�����b�tN�Sf�ō2���?ݭ�h	V����K�(l"�,t��u�=k>L;쬉�W����2��#=),���mwY:�w�M���5�R]��e)�՛B�c�Yn�㣹�A ��h�tv$VKy�q��+M�\$��V��|2J����\x�vw E[Sf�T��&��1P5,��.�3Rʮ�f�'m�#�\']K�U��c�5��X�j���=0p`|�ɲt��Me,�ak&����\�-�Y]o+-n����h�؏oU�g���RQh!�4u�����"�wc!H��-�� �r�� ��7�td]A5�y�]h��Z(��=+��V�b`�^9�LJC7��G9����ԳPR�ۧ,�;6Z�{Z�7]#.o/4]�ڎ�j{��_:�֧^�]y�Zך�3����Ƿ����8��Ǐ<x��ǌ��Ǐ<x��ǎ<x��Ǐ^<x���Ǐ<{x���O<x���ǌ��Ǐ<x��ǎ<x��|���T���z5�X��{�ڂ�|{j�h�a
]�0��u�|��ԢOP�k�p�x�]K����949��� �iWs��3��SD�GC�4�1Z`��Ӟ�fk��mt+�\���mD������j�Zoc8��J�nHK�@���Z���ق%���g�M�Y,�.���0�WPd��m��7%�Kc��=[G�ٽs+7��z�gƍL끭F�1.Ԟ��Q���9�V�A�by�$��}M��Fw#�#�>���0jH�ru-^ϭ丨閄�Ի7di�F��"���B��/vk��l<�Ҡyl���x� .��,O�$�]�O�䁭�&��QPSz�*��vw���煳[r��:4Wm��ؕ��E7K�h��B���B��}11mg����d�c3T��[$s���o��w�+�����t�Q� �W$6чȳ����cOmʵ$[.����7�%�6�i�YH<�6n	��)��-Z���b�	Sj,�G�*8VD鳋��oC���ʇ6��y�<�_�]�%���,#�Z�u�����V�3L:�ݻ�|�3�Wz�l�m\u� �s��=k���wZx�7��\v�C��_^�]uz�������$c�<W>���l���n�"�\�sU�5�z�����B��7W]ג��U����!��'�R�nճ��T�"���̽-;PX�Ucz�^J�W^4�En�`���Va�٪���9r�{��a�˃4Gc��k>u�\$�y]��FN�)�w���J��t�U�O:V���/��n�Y�H�Զ�S�W�SKz��[�����A������$5��윯�]�˺�6���6��[mM(�Ž]ʗ��V�ݝ����j�'�zi��HB�wuƭ"V���ѭ��Bc\�j��	�W�ge����[;�pZ����	�qa��>���!.�⥣�������&��K�Y��� ]��PZ�yv��Y��a�{%��tv�3�"@A�e돕݉�ei���|��u�:��n���Gi��)%��iJ�I��8L��r�.�n�A�1uR�	#�r��t�c����η&�كr�oz����ʴ�e'�os�8�׊���Wo{I�A�-��h�N��sY��K�n��]���:�hݲ�>����0mU4���kx;�6֗b;pT���v:U�g�h[2�tTE��у'.r�\�i�	�"���5��v{���o������� *�2_����~���|W��w�~�˿ٝ�F�>�tj��]j�!���DE
,�T�� -6�^LC?ɪ��F�!�c��p��e�RLA
$�19��gR�Ji?�	G
,�dP"�����D���-&�,�n�N�����(	E��
��RP�&��vX��?W��ꨯQ2��1�#)I$*�1��)�*2�.
P2�q��!�m�|A�牀��^-�K�����d#��aD�M�CM���@Q���]��_
E���xH^�V�@�N��q޹nJj�6��aK���!�(6�t�.Ů6W>�֏�aʱ��\m����'%�h�U��{c��f5�YZ������:�e4gv͡���̔�ygS���k�.on�>����##��,�,^�Ֆ��Ů�C�O`O[�׋�����#�}�vtu,�5�;Z�%�hm�R���Y�8օ4;�/��Len���u�gj�l��s�:�O��&�ڲf,�c��0]j�|)k������A�\M��=�R�[�I�V.�.���B�:�9W���r���Bnu(��-h N:O�˲h����Nģ��_[zweu��IB��і6<{Dn��(�c�&vLL�uAT�Q�p�хܟb�N�y髶w0���z��Č�6pw^Ɍ�MfK��[�5�vQ:�ڲ��%�����[a�+^��z�gok�zܢ���Y�51�"ε��������|w�Z�b(6a�#��es�`f�z�h����wŎ��7��u����HVR�N�`�Ԍ�.�+�,l�f�u��O�Z=�E��No���ٵ;��ww-W�Y*�C�-D�!"�e@(�p8���ף��4S�%E$11p�	Da���D0\
$�M���p��52�P���	hm�&�*���"ey̒4JP�$2�0H�Q ��А���D�8�b4��F�"�0��*4��#h��L�eS�4�l�*Q�Ia"qKa��i�)i�sւ*$�s�2H�($|cR�1[$��D(�ؕ)�d���Ix�,F����:��A�P �l�IN�-��N@�a�m�x��&"�x6aq��ԣ"����
��dj$�A$mF�0��
H`���+��*aMh���h �~a�\)���AH�!����".�3$"F�m�q����DePt�y�ף���q�["$�r�d��3hB�$/�!��I"$�� ��!
(�:#Ē	 �E٘�UK����SAUǎ:z||x���*�/3/3*�������{pƪ"��aE�Cd�fV�Y�jի����۷���=,��r,�h�p�&�莢��̲��
ݩ�U!�Ff%
eM�Z��ՍVF�T5��d���-(d���E�֬ �̲��hL3�����v�x�{9�Ff�ae�Td�Y�f9eefNNJLA��C���VUU�+�3,j��302(���,,,'Z0�Y5R�a��cd�fU���ǏOO^<x��ک�"�,�,��13,�2��ˬ2-Y��`S������ ��̦̰��3+,`��ǧO<v���>�Va�YUc��gQV�&���0���*�̾f���5�s,r��v��U����ӧ������\�ީ*#U�����"�5�y�R�QK���r2,����3�a�����������MG�5���"��(2�,�Yua�٧;̚����.�
��j���D���^<t���㷏~rɚ��(�fT]�Qu�Dџ3(���e1ՍMT��
��γ#a�u�5��Q3k�h��3��faTUڼ��Ñ4CEƣl�a��#��FC ���(8���Q���/�al��©�Cr�u��5�ZH5m�\	�ܖ��Q$���h�ݲe�:+�,Z�sͥp��H6e�?���FB���	$
h��M&�%��qL�ʍ�Z�#���HOB�p�b$���@(�E�i$��7BX�E DE4^%��	���*3���i[��t����~����0��S)�~��GVq�}7m��)��{G�G�jp�,��5ST�ܱ�=S�xL�&���Ov�c�DvMn�9W��u]>�s. �/�}�[Ծ��|��;�ח�9V������9��z��D�x`f̝���r������5��Y���Qq{�*"곟F���qߔD���=ez�錯{���"�'/����U��۩�>k��uv�`�ER�`���Z;v]�@n��w4q7�g�}>�������K�r����㲞6R�y�z��=]=��p��秩I�>��}�y�_��_]����e�Q���vWp���p_{�<V>X��Gz=>��$�u���Y���!�ϱ\�3�~�S�����@�eb�	]�(o���N�k���"��cx?9�-dQh8e_ʑֳI4Ҫ�F�O���A�_��eҴ���WI��d.���;ӫf�*n2*�x�Rx~3��W�TO�os+�vswԯ�����{Ci���*�ݬ�R�������@����������������t�n��\�	�d�������o���
�1Fz��:�3}�?C�y���"L���sh9��q�����}�,�1�F"3�&���df����\�?N����yB}HY�B��_z`�� �M�b�,7��ˆ����|�ϳ���Ca3�(E�f�c��ȱ���bғg�Cw��rx��z�(�yS�����z����m���~�����sƊ�OmSm���`�f'j}F��^,�p1^�.4��~ba�\R֙�ܷ;��/��u��hO��)z��2/�󿌶j����uG�߫�<��
��p���wս�v��jv���\=���2h(%�,'�ث��u�W�=�ka�.�*I�N�Mwp}�"�N��Y@yT8�Ez�x�b|7��χ&�ȶ2���x�^���F7���������^��8�uZ?߁6]�>��L�0|4^�sF�rU7�z'�>?|�S�r�t/����?F0Q�����l��o%�ΤG)�`4o4n��r�:��+Y�yG��b�-`�Vs�4'�]K޽� �rP��vٴ6Vms�J}9v�Z�+�ʱx��r��nNݲ�P��m��=j�ܾ��^z���1Pn�y`wh_x�P��;�6,n�P�uo�=�ĽV�ߏ���k���n��ޙ�秺���z�����3F�{�{o��D$�����R���:����C�${~>��։�5=���w�������ϱ}��U��3
���f�����?�Ց0��y_m8̬��Y�B�|>�� ���'ˋ���3�|��-�(����9�MYNu	>G�Zʷ��%SŬ�qO-/��o�����1eZ��]e�ϗ�7S6��yj?{ެ�����S^g�/S���֬U)�^��Qp�f���Ψz���o��=���=h���? .z�\{����ug�P�~�4~qv��oH<A�3jg1���k���ۄ��t����{��^B�t�g�٧��������_� `Qe�(��[��1��s̜;Rh_f܉}��i�'hjeMJE�EN0�5���%�}=����Jg(ޡC=6��{�S��t8��[/��w�v	:��v���4��ە��,��o�G��vsb�4~}�Ys{�b��t���.�}�2� �{>�~�U��&hw��/���D�or��Q{|W���g���U�瞃����(��4��|��`T���e���;g�Y��X)_}��a�kg0��'l��㹾ƳW3f�q���C��]�}]�q&��穹KDy҆����ϳ��{�w�\����K���v+e�z3�;o~�2���1�O�׽ r�	�{$6F��[��}�5�@����Vo�vo�$Y�(��WŴ�W{�V�E����;��t�tRs�ѧ�p<� G�� ln�q0_Z�&��1��-�덆�ʒu��A5ձzX��8)�O�pȣG@�{�_@�rF�8��X3Eemբ���J�B��.�5,-3����z��k�a�r&���ߟ�T�;��ގ�z�/ncs�}��Jx�������o��S�6�׼{ÍڡfAX�\��z��
�bƱ�=щ.|�=Q̧�T�'h���-�37ގ���o���>���oqI&X�Ny�:��t̜��T���VN��m�د�êL�����̛�����<���sis�H

�6J:`�A���{]��D��5�<��Z$�M�e
�C��R#�3�׾��/�%�?*@�N]��d1���b�r�:�s��%����(��o�<3�׏�)��_Ҹ|�w���fa��6�;}A�i�A������#�l�/�����>Vz}/ �_V_�����2�O�wi��O�_P�w触�oXY�9$E�sn�Ϻ���[�q��^#*N��W������(��Ѿ�c>c�~��}Vj};��V'?�ƤA��=3\�9#x�e�]��g�6e��jM�b�g�mV*/n�Y��/�����mr�}Fo���Ƕ~S��'$l�f�s���V�\�i�G��Gb!�6���&q읯�2���>t(�m�9f���8k(�X&�&����uv��P���ݷ�N�rj;��C[����A��@7ٵW:��j�["#A�"�c�"��$;<1�x�.���%��i�� 讍�5eq��}9�P��[j�3/�RnP��@m�������`XO=MM߶]c�/�v�%�H���﬋��'��ku���Lo�D@@��ǨH^kj�r����� >��fܧ�j��Fg�4uE��jn��\�������mL����wݘ��Z���'�4�47���]�QCx�O(<�����u������z�O�p|��3r�A��1��1ٳZX�1����0��3�o`��_�K=�o��x�����}��_�מף�|���i��?x m����d��T�;=WW}��u=�X���Kz���S��U�g��n罇.u������:y���-o�>�����
�^�$4�a�ƕU���C`�W-π7V7~���r�t�¦C���\=O#����2��kh�#/����U�s���P��W��-*Uqq�>�\��Ng���!�=�3���О�ޟp��}��X}w�4l9����׋;�=��� �6x�a_b`6���]!Pz���þ��!�릩�u��oe���y�sH.а��ս�ز�CV��`�t���2�Waʓ{$�)�n���r˻x�x�(2C�p2���k�e��9,���oLz�sh���hC"Ŵ���|��m�5�P���=�UU���қp�q�w��`[� �|]w��l�G���=�y�
ܜ_��^�r����)�:���K�dͯjM��UW~�����:v��f;z�$�2r�NO��8�8ߞڛ�|�m��D1W��k7�P�E�x����Um�G���>\�*~'"�yPj���=b��pƦ0��O��g�*FR�"��ꫛ���NUE?Z�oLng��3z�~Ul��}��ا;�n]�tW���F��ǏUٸl=�E?_�x�	�=g�8�{��!��׮����K���C�a�[��SYe�Cd���Og���DT���a��9��Ա1���}xl�������>ln�����E�5��+�nS���Z�z]{*�iy�(�7��t�U��*;2�Ơoc���X[5�9�i�X�-t��s�e^�	�b���L��l�B�΋]�N[wP�r�5mk�V9/�H醎
�`��2neN�fdS3�q84X���WwI>��ʮ�Q�ƐT��e�����.�@���^�]�^�Z5|7���έ�,�Pr��^-�j��N�t'IUw�k>�]��{� �o��#�}}P�{�O@�4Ǟ���8w<۾� S��k��{��
�n:���]νeh�d�AH�{<���[��;�H|R�>�n������Xݼ�ӿBbU���r���)S���x���Y��>k�4v�Ru���+��^�[+kwEB=)W���6)JAV}D���GQ��� 
�����t,�[����U]D��ʛ�'��'�N}���s̙[cmz箖��~'���\�Ů&I�8����^���^O�]ܜ��&������Q �v���7`K�;��������w��e����{2	*zL/��sk����S:���](5����P�9���c8i'&:f�H^9�y����P�Y� �ϼ뤵�7�4h�Ϣ�����j��'��܋��֎����q�4�0Mq=^q�}���뛯3~�+�h��E�1�d%����/UXs��m�82,�R����*�m�Y��u�,����2��L����妛A����.��W�o{�Q
�-R!�E���5 -I�
(����Ϳ�E��_یw�s�ה������=�&6L�}4.��%%��L����y�{�?��1K�yI�f��g��<�tz#��вe.���l[K6v�<ⷦF��bNez�Y#Fh�=t���3�>��?^����}�~̐p3(�<�h���<߮�,��Em�3C��/�EQ{}��������X��w�G�P����/7�s���op���#\�3�a�͠�����U����E,���u2�K�05^�7�1Ѫ+ՙ�y�k�6��˾5~�xÆx���W.M�8����[��h�{d������k'�˱Z�U�ogǦ��l1�������dEv]Ǫg�����.ey���B�rǝwe����I�8[�-�>_:���|���Oo}��S��H��Ҩ�*��ht���qq&�ua��kv��&��oG�5���W#l��:|�}X)�SL����6�A�4��op��|y���z�~#�Ik����:T��&A��]����c�K5�x�f����L�#�T%��8��;:�%�Y;&�-g~+�a��ڡ�;�9���_<���F���{�5�WsZ�rm���0�պ�bi�J�u�M���s�����N��m=oY�B��l���d�-�N����&v��)�����+��eo�qֆm��ټ~�~�<Mzll���{~Kꐬ��m�|=��1c2?J����.n�~��{W���5O��{�6z�Q߱+]��+�;n���A�{�Ϲ��g��0�Ǫ���>�:{�wq�&w���`� ����ٽ>/�(�+�7�e\>��#x�Vx��~��莹[ju�g�}'lS��VM��[�B�x&;�u�$�+� �~���.���xȽ���nO^�ѧ/y�U��U����mc3�.��.�r�Ydf5��/�~�{����v�	���n�%C^����?Ho� 7�o2�E<�����~��=M ��̛7�=|+U�ܤ�lkn��gS�f��B�ҫ���Tkd��Ih9aC�4ދԆ,}qn��V��/pQ��k �ul��1�͊jor���*�:��y��o;�A���Vw��ޡAJz�^�ÿ[dڧ6NS���A��̃Y�Y{�j��8̂*M��kK;�Kڬ�⋫�j՘�wC�cj��6�@�F˂���82��éD6���'�M������kl,�˝{��8��kz����(P��p�K���*.�g�������Il���:�'�W �i�q�jj�4�%o-u�������:�zn[K��⫞�w����>I�ݟ1Zj�eɬ�����2c�U��rX��0���}q�`%�mԅ��f�:y�d��Q�$ӝ���
9�����yf������s����(S���Z�T���]�aڦ�̔43�)���v�s/z�l���!W#t�No;Ĝ��Dp]�Y�掙�R��|c��D�3�d]7�ej��fl/�`9��h��}k�
�j�
lm4�R����
WQ��\݅��v���bS��^�vM�9�*r��2�G���u�se͒:��R���ݲ�ewkRݓ��s2�oq,ש�Y��Q��l7&�l��(C�ub֒���9�B�1��% $[����7 �����B�B�3��Ju�~D}�����C�_+���0bn��5kiȌg��~r?-��c�n.�D�@�k�SJ
�ltݩz��l�Z���tm�������|q� ޚx5Ԙ<��k�;eq�,�έ:$��ަs%h�j�r�(�m^N�I�引��L���5}�v�X3���!���`�:6��ywdJԣ�u���+z��۝-8B����鱄��֦��Et�}�zX�}�[��j"�T뮴����������tT�(�&�dw+�Юj���=սY�^ON��=�Y���L���;�`z�WL�fQo�V�L��P�l�o9�î�b0w�po��u��[�uu` ��U��."�i�H�{x��;X�0���eX��`��I�Yc���N�a,=����R�up��&�߭^������ԫ_:��9.2�\b�yڰ�:~<����N�V�~޹ՀB:%�1/�Y*w"���ڽ����ᇌ-�"�J�BfY�÷��q��K�PW"���nN���#�/�;�#���n��D;RTV��aTŎ�Y}�!��*-}G`2�h�K�\����r����p�k�6cLPU�2���5"�ާUJ�.l�4�K��L����<���M�&\|x�j�g3$�ܩ��k���Y������ͱU4DU11DEUAf9W�)"�J�0&*��"o^�ޞ�;~?�a�D�U3UMMՅQ�4i����2b����
fJb�fESD��|zzz||}x���&�!���<�(����������<����*(������"$����*x���ӷ׏=��U�̐�fT�Q�3�dIED�T�T�U4�A{�|~>:z~>??�Zj�1��)#�Ȃ�
�,��ë+�"���
�VSQAL�$EǷ�OO���>yQUOy�S:�"�̂*h���i�j���0�".�0��$�ǎ��;x��E�TPET�Yda3��Q4Twd�G��xXPTR��y�����o�o�o|�*$��&&Mٖe�E�Q���LL üȚ!�x����o��8eT��DQI_0��:�k*��"j(b���*݄M3�F`�a���d�3F`d��L�׉ �W�$p��.�|vT��\������iE8��!� ��w%��3;Cü�s2q���{�o��-���d��5�
�yx�u4�]�;��L����gͰ-�Ư>�-�`����u> g��,��A&H@�<�8|�����hQ�֒�����v�+�}��b_����ۣ2G���k�� �"E�?M��6�{�nlF�?*�!����ؐ����@����/y���v���c�j�
���<F02�e�[[�'�s�G�N�=+ƺ=��\����a��	���OBj�}P0��2���b�JAȹQ-�e�ͮ;ߊm����f`�V3'L��|����E��oq���5 b{w��SVZ�Aܢ ��j��q�%s��߶-�qWnK���y����^��t�n��-�VP��8�1,O�<�ӎ��!��f�	���գ-���^oJ`�ڑ���i�L&\�� ���<%�h��p.ʝ�o�ge�ǫ���h�E�m��9^W@	���b�}�� �)F7�|���� ��%	��kh^�ʶ�֮W9/�@���|��ڧ�.=���z����x9�O�pf�fC4{/�CP㑀+�w�i���͋L\K����g�ڜ�7�{5�͉]PvI�+��x`as��76o�k�@�C�^�R/�[ԭ� ��c����9m%'�*Au�靵/���R�³��O1=�SW��&zm�;m��wE�1C@�E��޴]��3S4+���moߢ�b<��7����/���	ovv��T�W>�U�!�un��	�}�J\eY4�դb�QN�I������{��`��oTw	\P�P��W�O�� �X]t%���=��_��%�sԸ��odO<[� !4�զ�]�t��n@ޏssL=zy��c�e3u���+�rd/�jȽ���Ò狁Q�H��|���G0p�y�0�I�D�a�ru��������g�l�S�H�폳�f�`6�nmRa7)S_m��s�m��[�V='�T��'ѹ�~qxH��7��	𾞎�(������l��:���R�g_7j@33�&s.�ˠ8eNi��ChO��ϧ(Pރo@���ʃ6\a"��-�}];l�1��"#�����^����ak�����*�(��y���Q��>�u7����[g�<�g۬�g�po�\���_ +ܢ�y�Ɩ���ɄG�Oc)��@�������/��%5�M�y�����Q1����"٤��O��wU�6�hޑ<�,^�Z����~�)���@S��Ruf���#"��yN4fd�P���� ޡLo���w:a��x��V2�"j��3z���a���}�o���Aȶ(����35�ӯVa6�WB�ƪ��1t�>k�:�E"��-#DT��$�<�EҰ^��� �jϫe�������Ϻ�V�>o����߈��9��P2I(}�a��l�ո(������p�q�pT����lQJ�����bv�B5���4;�Sh�1A��vL�*�v�^���<D^Dx��>)y��xI�6#5��+^~�[�r�r$�2I(H��H����Γ������<�_q�D�Ikk鎽1I��ܡ�E[���g]�Ж��"��[�q�@V�C���E����ۓ�ř.��5�W�dУ����P����6�k��˛~�咽����yA9��Dݠ����@>�����fA�.��k e��i�cEUX��Ԯ`��Ƚr
�c��8��z�oP�57ٚ���L�s侊�{�MoOI��1�N��VAC$�t7�N���q|sR�oڧ���
�څ��Q�6\U���Ѕ������>y��
sZ+��-6��%�z_G����ǋD�s�-��0���ْk���'�sn�ڦ`�ݸ.%�Ғ��<Z�w~/ʣ݀��+�pE��OA.��?�ZRXb�{��Ԩ�9X�*�7\����ͯN��^�4 ��aE��,�<���*`<�LMЖ���)�TyK$��y���G��X�^ |zC��n0��	�����qMM�cH|�N*V�������J��.�[g>3ӯI��Cm���6�>y*����̟`���g��켨qv&�V�Ew;�T,Wc���L-+�}v>��J����h��:�MK�rl�t���3i�5b�y�j
4��0H�q�K�(bm�T\z+���*!-���L��{S�4\��;�v�u�\x�;k5	������o3zy��N�Mq!�I��f��} ��X���d���hx����G�2����{SM&���WY�-y�^.��Y�#���Z�������]u��jtJ�틗����}�Ze���z��\`D���`��;S XÑ�e^%�d��z�\=b.2�%[���mk͜����4���x�K�gMm"-K'�q�R*)�ҟa�8q��C�Ьyͻ��2��feE�����w�(��,�,� ���Շ~U޺���M5^�b�e��d���fKM�ꇪ{U���_t�8麟��o�@���FBHs�u�4[ �H���5:�*3�a;�>��;y�c����c��y*�<��6�J}m�(�̘��Ƈp�jE���]
���z*�I��ա́��H���z��It�ҩM݉U�PX�Zܔ\>6�����.� ��i�ERŮr�ƫ��|[B��^q���ݥ+�c�Nb��YQ��B���<��(j���f#�P�q��G�	^�.ZĨny��4����R�d�v/�q����&�u�v��_f�g���=����Z�X��cյU�[��2'7��8�]U_,'sR��^H^+U����K�ѐ)�|ƿ�d���]t�'k� �ڝãhgS�L\7)M֠���w4�UuZ��[��`͝�[�VsAr��~`�&7c}X�4ӧ��{�����R�{ko�˻�L�\g��M�o5@CmR�->��u��E��`�n������TB�xn̈́�Z#5�6n�����b��������P�:Q�'���M@钓���e@^o�H���l)f��4�.D���g�g�Bt�@�������D�][��վTĺp-�=��Y���}Y�U�P�ǁ+$N��aaI�U�k�����[��h�9��Tc��%��>��	�so�lI/Iu0R��Ԑ^�����Of֕��F8vP�KP�R3͒v��3E3;;����48�'��������xL��a�.Qvo����ZZ\ �9���3b~`~1�g�^Oq~�q�0�s���7]���'UX��X�|!�vٴ�j�L��h��v{�F���o��'asĿ��QM��O�9����^��Ӎ1�|ϩ�� ��1`��,SM���J�&x�`����%`�V�����͸����b3*��ռ���[�f�A�c�Q,�,���~�YB��<4�zBm�VS�|`����ߝ�\�L��}��@�5{G{/�#�LW��*��ֽ�'��{�z���9ٰ[9r4Z���d�ή�c��4u'�RXյgm.�����}6�,F�|r���[¶�XYy���t�6�IV�`0l�{�;���:�0�o��&&�]�٪�[��&���烏��0_�E+��2)��*o�ֆ�w�ZV�MD���|�ٲ����=��F-�iO�/w8�+!3��7]B��A�m�s?~d�m	�����7/+z�P��e;�Pfk/N���Hm�a!&�AvO��f��щN���F��o^j�SM�H��J�t]v�O �׷S��v��l��0�_?ث�~$���,خ��C���J���^{U.Pg���:ӧ_�����4��B\B�	��Ȟp:㔰�PC_f݉�&�dv1=G�Nɯ�,��q>��Ϯ�>��1���?l�epT+�����t0U^� ���:�M��Zg�e{�u�=Y���}8�0/p'�o	߻iذ�g�mLT��&s����r�Ǥ�dO�`�Ǥ[p:DeU�#�b��G'b1\�W���F��AݘǙ�8��FD���G��gP�z�v04+�b���3�1��F��;nv^�K�o�#6&5�Z'@�:����@���U����6{'��VyA��������*8�)��ˮ�*�VK�w4�${�̕L��b����Tx��D�|�����nbC�pco���!�\I�C�ݝK.�s���򭥷��.>��q���̒i����N��Y��	�<�w��
��l�g�'ReW��4}��$ɛp�$�L�q��^���6�ɳ�_��_���#����BD	���I����а���'�E~X9D��Ɩ}���V{��`O�%N��)�0���9�r�7r��x�n8������Ds4�tI�wU�G�TO�<�Ϟ̉�S�o[�����Q�s"����[���װ�c.~N�a0!��w@?}-!=Ѭ_Po|F�UC�I��'gkuFf7^�0%��;�u�oAǬza!D�x��O�sE�Y�{�q��n��8U��>�w-�����_��jeg�[����P���@-cS�hޯ��]��6��.��e�z�N����^����ra���z�-�Qm"�1��',ңHfd��WI������w��`�9��F���K��^J�������VN���Z�C=�t������4o�	�R��QooV��Ⱥ=�׮K�ٝ簌S.~*=�Hݍ�S�w���8]�d_<%�m/B�T}M|W;x���~��{�x��-�%�R�<�z�v�0{��a]0��ۚ��ƨ��*V8�0��_b��;��Yr0䲳��,�[/}n�Ľ��,�lPθ�q�Z��D�dw��G�E2�� ^A��c�������6�:�Hv>e�a���ܹ�cF�"�g+���%�� ���W��z�׳�#�^^�VGx��z�Q#8�Uu[*+[G� ,���w;9��׫	�YB\}�u]g,sA���Eeo9�Z���9��[�}�<�{s��e&�2La� ���Bc%��7��+#ı -��5�K+���DD�_ەhش�\I�t�Ϻ�Ɏo��'[T
N���{�dS!��z^��f/��S��唊��oPEH�g_ ��ƒi\XU����6��<��dc-QL����հ
�|�`���������D;�^2l�dSr�R�Yվ�7���\�j��>7��ŴcѨdD7_�6������G�>T"?�w=�1����K��W��T֊�iw�1�Oݞ�`3w,� W��j�2��?����q���bt�a�O����OX�"���o����1%�P!)�#��3��:a��7S�t����9���x�/Q�gf���JDK+�<��@�߾b�����\�-�y�2��Hp=����<혶;i�^�s��lD;�v8�&�$(n{iǒ�.9���o�۩)�V�:�C����|G-u��_U�~���ٓ���q�O�ۗ��zw�f��n1L�!��MϹ�B�l',��)w9��*% 2�5?yRN*��x��p���L�'՟��n�?��&CtZ4��\�5Z�<���q#���V���Q2ҳ[PvL�q�����5x-�
�˯f?��KNX�K&�
2>�s����"�줲�n���  0/��w&��X�������D-kn���Y�cl�����'�(x�Ck!��q��t72���� ��w��2t����jd2GV`�`BdCR���Ng�/~}K,C&�ag�3)�n�����M�N0�T_L�uQ��� i�Jsc$\Y̡�|�T�]���&�]A�;#K�}
�(����)�~�Sm��B����|)2�8f.���!��A���J�A>��F�ۄ����vn�5�QqF�{�m>���%I�Y�3i���l_V�����q^w^�h?��b9��J�ן[��<�¼L-�J�5m�2�j��v
�wv������@^��	�Z_��������X��u��~a~����*e�mH�����~:�k�1���1���Ѐ�qOP���Z��ÿ�A��`�����/˾>Y�L@���ٳ��s����ƻg��Ԝ�T�)e�<�c#[x�yڤ�֒E��Aø����
x��~K�Y��;g�a��v���-��랓���AN׷��`��/�{7���'$No�)n��v��͹����A���m̀�1@�����F)5Ŷ6>�Q�$��A�W�z�E���N���ZJk��(t;�Rxf1���n9������tfW�(����"E�c�xw�O]��d�}�ht׍�up�M�%f"z������y��������b!�YY��̘��k��O�ϙޅ(�BH;iT��Jq����N��<dyXNۻ��M���X�s5��Ipe�i���.uj/�Q�P�_ʪ�������&$L`�1�9.��d2d�2�̔%-)AT�4�ST�R\�����.��q�ur��Ryw֟;����G���FéL���\{���v�wʂ��ګN�U�n��`��zC�	K��~�����_N����1W�B7�UJ�`�P��f�����.����3�^�p)��=�c6��|@:�}�7�DFb�"y�z#�P��[5��-�F���˷_-�Nm��m�LõҨ����1�b�F%�+*�J�A������;�0��N8o�3]�I������j+�r�;츪P9���ml��F�&I�9M��q�
�/v=V�0����Qp��E,�#u�b�C���ԝ�wH�o���Jr�0O�����&�Eg01�"���n�������ME�@-�XlaCxϥ�2}�.9�_Pf�T�
���r�\�-dNŜӌ��f��_uׄ�;q�ʉ���5�b�Xt�FЌ`��:����u�/����~�t��nL��G !7fB�\��?�lPٌl�.�n��������5Gs�&�2Dj������o��+�l܎P%��gy�&����x��`��[p^K7��3�7�#� V��{!�M<���w�b���uC1��,fpvW|�.1$���b�� �Ԧ^P��3�]1��*2P"��G�I�[ʓj���ۦN�N�ۖ�BK�)>�&�N5�./�0p�=�{ǖ�v�Vz�����l�5ŷ�i�r&\�M�]c��W}��J=�p��)v@vI�s)��X���$Y�
�s�D�>8,k�-�r�Y�|e�n���gc�<�R嘯c�S>F=�]��*֛�m���k��MN�������f�>l�ϖ<$ÝWҨ��U�G
�z��p;�vrgG|6�t��F����a +m�	�p��6�J�'�w�b��ʆ�[`�uu�1�/�ς��4"�dL��MA]��;2X�w�f��nR-��T	�r�׽Hέ��I�c��OyM<��դedz��q[Z\���֭�Xc��x��-�=]�fC{}�  0y�����[YL���}���;^	��d�,���P7���9/���0elf�v��,-�{;wP��w���rU_aN(��mH5]�˴" c�ժb�fd��27�(�W%�
M����7Or]9�ݺ�Z�&w!�{pN�Kh��|����W�;��E��M�xh6�W�l�W*�gV<��*jq��+u+*̩g�-weY�j�8��d�7Uǚ���]E����\ݤ��0
@��t���D�V�wbމ�9X�[�6�@:�~ޡۚ�a���L�V:��������,}��^��Ӓ�
hy.�[G_M�"�2���6���K��ҕ��c
�U��`�";2Lf.�����f��W*Z�ܢnZ��՗8�ޅSQ��v>q��C�`Y���AT�!S=���=J����x���/���������8��cy��XoP��(�t�u��@�vb;�=��S]2��v͚)T}��q�K�P��m�Df�����^N
���0nJ�<���!�5QJu���oIܝ��a������{������؝C9����o:�p6�k(k�8�«�s�Xy��Z�gu�1�U�NG�`	'�u8)S�.K���s�BQ�(\�;FwO�Ed�W�c�ס��4�����;w�(�-��뫦&����w�����ڶ᳏��n��ۦ�p��a\H+/��=CX�$��r�Z��;؎���v;;�dfV&[u���E>ެ�V����5�˨���I�����5�h��d���w��hCr�XvD>��1�8�
�Gyw%����F2x��(�u�����'�"����G{X�n-�fyi���p���/%���dT3���Z�0�[#i`��-��M��u�7k�`c���=������%��IV�f�sS��A.U����=��e�XǵN��cBRL��%c�Eҿ��i�&&� �(��0*��b��i��2*� ����$E;#��)*����}v����򨆚J�j�*�h4c-%'# �*�k�ȵ�ITS5MEMQ��MY���=�=�<x�{]�DTQJU,�SN�$IM��M3PTEo2j������ǎ�>�v������2q����"���������**�)����USDE5Gx`g��>�}x����o�廢s�CT�5ULIQDMS�f�� �h"(�)ퟎ��_���$������2���cC@���XKIQ�GQ�Eӎ;{{v��螓@Po�����$��Hu&HG����3�(�*CPd3���۷���ت������;�i���)���L���pkI�R�:̧�q۷��n�}����0��ʩ*�f���2��7�M%%{��ugq�fP��UI3M!�]�s��4Tya$EFC]FE'��#��|�Y�u]6j�3Z��Q��)��j��i$��6m+I��H��O飶`p�7a�,�'jփ{k��i[Ȫ��������G�7M*�V��1eQo��v��T�Z����RF��IN	�����"}�Q�
I�"��2A�.2�HF�T,p\&I$n2����ؒ$�	T�JTˣ�~H��3�*�!�(�ʤ�$�������ٻ:����acZ%��q��6(��� I|�)}��PXs��o����|+;���G��3�"�5?����ot�dY�"�m��ȶY��xmfA�����%�Q^Ǥ�#L��S��8�j<!�)�vcN��k��l'��4�B���pt��!p~g䎏�S]k����P����ۓA����e#�����<�Т���S|���"ɹ��k�mx��h��{C�R.��mO��߆#V&��Ҿ\���C���:�XnSro�pc���3˿*x����A�\[rt�0�����r]���1�v��μ�<�M����=�E�IWA��u���:�.φO[���a��6�*bL� Z����qmWp��]�e�e-��(7X0!�G)��DP�Վ⁘{r���?��n��4QY;���w!M~aɌȧs9=.�����c��^��m3-{UcKSt��%�B�Q��TwC�;=SәwkL��'��Q-I�}�FOx3U<&������+������c��f�\�r���?ߦ�(�e��X.J�?>�{X'�O~_�?L?\�L�ߺ���+-q��B��o���LA�J��03�MS�twK1��d8�xs�	�}�AV��I�i��9�d��Z�]}�d�eP�
y��5bu���aQͮ�U%:�+JF�X��uy��y�Wg0�[=�����+�PL"*�ʡ2&H�2�x�"L�
�C7ߟ[�ϯ>���y�nq����q���������|2�=o�)���"Dr�gd���*q�&{V��7Dt��Fv\
���tS煨�[>��x��M#v6�NdG0�{��.�k�����LZ��� �7[���P��S��_����cJ��B��1�����b�^�{�����z�j�T���z�FD�1��q�\��2Y'���+�׭K����ש������4��8�`_YX����	�_۶�
�S>��ǵ�=���-�8�H��r��Ru�/��%�'f�!�h�x�p��������%��IoH�EXۣ\�z����?K̯���'�(D�D��[��0���N�t@_*"�	�'�aQ�����}q,��e�ruo��Lbk�435��PΟ��܅��7~���dw�ʉf���4D>�%����Np�1W�-{��j�l��a!�lٜi����w@���_�m����C�;>?dG�KTfe4jjV"n!&`���^�T>8���k�Xh,������8(ߦR�%>��
�uF������MX�f�d
��B�Rq��w�W���!���<�!%=r:`������ܢ�M�T��.��9�
U��J�]�Z�����J���ܪ��Td7P������d���@��f٭�C�ڷS)pЪ}�9߽��=�G�������d �2"̂c(d@)�UI�dQ�&P2D]���N|É\;���C(��\��Bj�E���.4
�,a��Ii��[7?FЦ��t���%��:J������v͠�9<W1��ʄC�OW�d��@ɯ�&�<���'0r����^(ڌe�-��z:x}��_՜��F?��F�2�����і�%
n��ݫԯx/ �t��Ω�׷�6z|�RʡX�b�ٻ�|�#�� @�ߌ{�??܆U�@�>���Oj���.��پ��@���T�}сt[rڛa���o��b�����x����
і�D�4��L�i�1Ycױ�4xY��=y�$�oK�t������[l�6�\�
уz�Y"s�ņ6�{huO�>�-��6z���`�6
�.(RSظ3i���a�)F�zI}<�����f�0*Sǌ3�}i����ȥ-����hE*�y�`�A��7f��+����AD��A�梹&���ھ&�|C��;�R�_�!�5�|�:�2:s��@z��4���t�J��)���_�6k8����i�|���k���C���������c�?V~��;`���I�&��ڹ]-K�ʞr���>�Ϫ���C�|C[�lS;b3v���>�R��x��A�2��[O���I����n�Gh�j���85���ʷ��4{�{�>�W��\d�E1�P�LaҬ#�D`T�	��7�vs͝�ξ����ss|#�MCw�e��s^8}~�z��>�\M��C-��q/��PT�Y���ڹu�~hJ1���6<1�>G�����ڂ�'�z�kMpG�������+��v�ӟ��l���HHRИO�����{kd���m�
lj�<\��A�/�4R/�բL��{���G���#Gt�~�?�E��8Ј~��s@��/�n���u��U��:�c�MgѶ��sT��'�Sk�urx�GC�Pt'��m+*�ypB��#�c�ΰg-X�
�f�����#K9�R�-����Ժ~��wR�'m�T�Q�{��k�p�}ގ���r�^�>��
mah)���a�/}�[�۞�P��� �����(�V_�ߜ���XL��uR����n)�	�/"��י1jbY6Y+f��^jȊ���pܢ�$�o'�����jnA�τ��8���|ɝ��/�G2籊)>��/����b�	OP*5�#\o^Zyf�a��������AS>�5�RF2�k��9�J��巅V̇}�>{�����$�v�ʇ��W��:K�DR;��b�����Kw0�6����a�YY,<�fa�7hc�}�eu���|0��7�*��0���:6�4�v���V��ٛ(ʺ��M�����o1���˩��Ns��`����Ͼ����ʁ� 2�2"�)�
�� L
3*����6;��UtZFdk{��Y�h����:�&͢�Y���u�|Q��u�-�Y�b�4\s5�l����[�diǵ�SWn�.�d�|�Nw=�P�_��7�p#ù��2A�C���L����ɋ¹�m*X��ە�gYr'I�8ǒ辘��H忚��]0�0��dQ?ܷ3���2���៟:�sp�/��[�}ZE�{�ɒ�t� y b}%����"0���equ7wփ����OR�΋�./׿AT7��2�&��P���.wɆ_1������ul8t�$�]�+t��n{Q�`4P��	q��4���"F��Om��SQ���V���Ȳm�1d�@a�~����AӉ��{�D��c�~�ox���BƜ�n�5��m��]�j�tx����*	�w�2����_F��o�n���[&�/�v�a��5j��ke���3;W��~i��5>�*���[:z�]��OZ�%N2�Ge�5� '2�a���խ3W�zAa�.�e�C��<>G���i*�4�����>gQ�����pGlQ~������8�6���wIE��;;v=��fz�CKw,ݍ�������	��7�úR2���j@�Gؘ��&P@�!��tcxe,��v;��v1�S���־�.�9ٹS�f[\�6�#�����-�ڽ�5�����fA�L� �E�V`E�fD�"��^�g9��{�\>���M8��p�÷�c���r�%�GD��C�6� �y�"�ǻUk��;�h{ff�C=HL��%�<ӁL#���g̒K�^�ϰUЬI۹���N�N�=���|tT���g�h�VU��$<��O���H���F��&<�l���M'�R�=ۇ�/v�M��3x���0��v�Oo�ًgb_��0;�jQ�~�g-+�-4���+�	�i��}���q�ؽzY�ơ\�r^��&�Ê�x�=��/��g�o�m�y��S�K��X/�*����?U�˟�>�n��o��"��.^C���Ů1=1e}�ٳ����=.`D<Cz$�R�5��t�h�ye0���_���~�<�EJǠ��1��K���46�t_C^���a�%���y�m綄�-�<\X�j�����G��aǈxrո�;��x�-��[c.g0�!���y�S	�p��h��7�t	�\Y�t�*��B�X��NstB/�W�O0��y���f�!�p�r�����3������ݤ��3�������*/�-�Y��wKY��"�I�J��D�V�"�����Tn>�dѽ��X�u�K�ZE4+,�ֹ�;n���#���Ty�U�ś��R�I�.��Uq�h���Ӳ/.��[�+�E̞���ʫ{�Ҫ����\8u�K� �x�d &d�	��Uq�@�Tf\���ߙ��)Q�(ёM��c�!c��j�i�{g/X�;�'�a`����Ez����g�Z9�fX���%����`%�Ǽ'�8��5�ύţ�a�����	ϔh�?�b�Y��lld���J�S�%�^����7�	�A�*��7���c"K�]a�S0�5�1˶M8�.{���{���Jf�G>���}�
c^��D�b����|�ۇ,g����IN0hi�0+��Q80bը0��x~V�N�aӳ;uy���PTS���-���"�|q����C`����8 d��m�b9�n��r�G�߼l�)���C��O�Gʄq�SQMӒ�+���%���ke���C�Gt۞޺��,i;n^�Wy�����F�����×=߾58�IQz���/[ �&��3SR��Z��U��U勿	ŷ�;2�=z-�]��O�ݴ͑<�W9�ܞX�o�� �Wl�w3��2�n  J��:�c7���W�O��@j�aO��xgq󖯶_%lq���tde�ͺ��CE��#Tz~�.�X	T���J᧘Z���F�>�V��\�t�0�������H�و��y)�l?�a��-��]N�kzq͎�H	�1��˨/.��g��D�Z�^BW5Iqr��d>�	*���ɗ��@�e��6"bl<^m���Nb�7+p���J8�v�B�`'���y�s޺���ڊ���̇�d�E&�F`^���7�����¾���p)�_��[T���O)���$���}�qR��1��9�OZ륲�<���6��4�K�Z��������@���e�|Do��Bs:����3����ȉ+M9W���
&�Fw?5b�������m��ö��	E��~i&5���+����F��]�����"b"y�Eo.فM���Q�]Cz�3��c����^�ٳ��44:���č��I���+�!�3,��yyd�*uU���Mt]u�:���H&u��"�~�Pl{u��dU��0�u�����~K�h�{�	����W�����$@X��w�=f��� e��C�z�k���B:���esM���&�fmu��L$C��(HQ�����ض����^�P𑑹{����[^"���n6��s�b+���a _�"�U�S���,}o��~��D��o�vQ��{W���֯e����ؒ��4b�j,O�M�ܺz�<��K�6�� K��	��nW�^�|��T��������sܙ�ˑ7���x�s��O�h*T_���N?�s��j�l��ߓw��?~�N�������J]"p�FzwJ<�HĻA�Gn�\O?�����P�帓�����H{�~���`��7��K}�]�����f�+�TF�b١�f����ݐ�/3c�Kp>5�̍��߉���b+��l�]Fy�Y�}���(��=���(3d(�2 ̂�" ��<=ul�3dD8��S�.H�����d�+
4�$#��b&�&T�E���1�:A��e��y�	���Y�t��(� ���|�8n�*��#�jMR��čJJ�o
E3z�/U�%��,�oY���,�p��d�*�[
9B�� ��'>u	���(�1�h3�3Sj�ZD�%�O@M@-��έ��Йs�(���G�g����6�T�Ofv�r��{lۈj��/
�U���'�P�p84J�a#w8��%R���]�-��eq쾆�[2c��i�+z��e������3��£��d�y���gHfsY��ʷZ��h�V�v{	�����3i��)ҳ�t7GV�v%����-@^E�7X������t�$R���7������m'R��rᙙ�|�#��R9^v^~�v�1�>l��� �S)�;]ܭ�{5�钬�*DZ��+�y����N���I`�b}cD�k�6�Q5�;3h��^�nobY&� ;��C/:����p0KκOb����H��r�ñ������]/<�N��RL�nn8fPŲvc�C7>��f�P?-�Ŵ���"w`�~�|��7���v�g�C=�y�lO�����	J��ǹ��,���*6�=��h{l�i�o(fA���]r�E�c��ҷ��V�34��++@�Rf&�׵�M��ù�s���^b67_؞h������Oja�0���rJ�N�7�}��l�A�N�T�`A�@fT�&E\��{6�i$9��܄��Z};� #��6�;ǝ�6�v���H��ߪ���kUcm���A�4V=f�.;�D�[ב^��lB�N)E[0�/`�ԥ�6�B�2/�&C��V��T7LA�1��CY�W�O��`m����g�r���?圢[����yg�?����q�,�!�Û�j��g��mO����h���PO�����l*�4�f�a8��j��^tP�����yτwHt�πKո��>�c�,�1�����eV�
m�jm��[$�b&fjkB��Y܂�������_����Uj�¥��i�R���P�]1]Ag�"d�ZcLf-�-��FLL^m���ן��!���5SGa*Ϳ��>~�`*���1�Y�U��Y
P�v�r�q�5����M��������TܘыnP�=��n��z}���\_��i��T��с|W����rT�Ř����:�%>S��ؽu�r9T\�5��nq�i�g^�����7r��� ��]�/���{$(gqW������W=��8���݃)�H�r���؋�o��� 3�Z�L~�e��r����A=����
�<Xz�!@���ֈ.=�W�$��*���{�wKjVx!3��Zb	�љ���)���;��=�X#	PK�2U��t{5Ů�]-���;���Y-^\>�g|4�ه�)�hE6�'k݄,��o��
�v�P��egNx5S�%�]�z�m�I`��I[�M�hdȂ�\X��	"+����]Кtc��DonxA����c^�{qSŲ�*Q��n��W���u'��sm�#�d��\�daN�/(%��JZ��-&�:��Y�:�1%����E�����U���@'V��N�+�.u�L����D_Lx�fѹvr��wMv��fo��ыi�Dy}ُoo
�|z���f����5�Z7.�Ke�2��.��RLɶ�p�x�S� �[��m�����0N(��+�࠴WB�k�����i���@;.��&K�N�����G�5h�%]I֙dm9�\���A�(UCX΢F��	�X�	fWi_?�C�b���9�_;pd��re1��Jzv�!�Xf���.e�ƺ��<�ٺ�Ǚu�Ga�6+w4Y�`����	�$V�wXY3.�Bj�w+�+���Ԇh��#۷!�a��m�k�m��rHW�N���8;��L���r��e�}�oo��B�~�e��r�W�����/m'8�	��ĬEݐ�l��o����L�:+	��	TZ�Mtp�v�Q����KؓS�4�9U�xLsD�q��-��\�}C^���!��â���m�1W��w����ҰK
>�yG��ܩƵs5�\�fo�6wS8C�������<�2 �K�.;/f�V��E���.C"���
V���IڏMM���U����!��ݳT,.�c[5��Sͨ��-yɛ��K�\���If�P�<��<��mT�4;!k��uEҷByt�at���{)���E�&p�N�V;��O@.�����n@"��,���q�2�|�7���N/X��<7�݅86Pg%d�x��\�ae�2!Jڛ��͜���m=�1{G4A���y<����މ�l�gT�=Zy��D,�x�l�]Y|�棢����z��r^��Đz�i�{�hM���'JX��	��u��1uogvVvL��fr��� HIEWk�ˬ��ν�BwH[�,-�ͳr��/�����OsvmY����q�B�`R�4Rڹ���p�#/��5��ʴ]ϓ������k.>%�2���g:U˹
����"]�n���p�8_Q�Gq"C|��x���%�������mL��6U��G���{k��9�r@����4�'8l�k��nH��������2�rG��2L�)h���-MQC�d1Qe��EUE,ZΝ8��������q'	2B�HrH�)I���
�<����I���q�������/r�"))R!"(�<�S�2�	�d	E'v@�Zq�oO��]���4�SAE	K�fY�A���P_3 "R'�,�
H���ju:g>=�x�����^��RV@eQ%PT�y&Bn^GP�$M6�)���*h]�8���׎����2i�r�ueB�9U	E	�E��t���o~%%!P��U<�����Z����zx��������'��w4.��!��.MRJPud�'N�t��������2
(����
+S�TPjC ��

F�>G�G�(���`)H�C�@Y��T�2SAfHR@�D���V}��泆~�o�Ŷ��o�����)�iгu��s&gm(��3[W��K�y�q��鱠I�M�ַ�~��󭿀�}��L�
ȇ%Le �&�� a�=U�h�5�ߟ?7|���7�t�����/��
0[��sR�li>��©X��&�����%�ժ\����"���(���6���s�+،��ɞ0(�������R7z׳
�^f�,�'�aCg��-Z���}n��5�w؏4y�~�T{ F�P���v*��2���]3���x���,%%��v�֐9�GB+��%��|�]�^S��>��Y��MV�����L0��hm���P� =HhkI1L��`��6$@����}�[��]�i�5��\6�����,�F4��I�{zY1ͳ�j@D�,��`��_0O~1�����'�����y��}������L��,��s�� Ĕ1V��4�����@�^���e�`n�tE�*��3�� ��k0rϐ�o����!v��_t
_����*�������ڡ{��B���gǯ֨� d �|D�_}����c�C��a J�������g�J���w>��6�1Adߛ(�w>9t�6���x��߅U���~f�[6=������)��ڳ�N;ѩ��9�fVF�?�f\<uwo�ޤ�3+�7t1㩨n�
���c��Z �B�ZR� ��Y!��~>U̛���nH�>�k���3JߵcS��u0]x��X��ɏ��﮲��l:��7_� ~�*�ȁ2�L
̊�%P��.�6�]cPo7�8'5���[L�&}[�0��YWHx�L_ǿ\��X
�ճ��c����kc^77�����ۊ��dX��k���c��n��
��Fĥ�uo߸��w�_�S�	Q^���ȿ���E?o�l'�0�q��[�U2�fe� J�QQ�0�=����3wY�ܰ�'&���f܊��e�X����{I�z����t�nT�[qf�Z4K��M���D�;|5kZ�)��z	ŵO���xϛ����:p�Bi���3����.Y�TlF0T�C{��~*����Rb,R���\D	߾c���F�-/�Ֆ��iOW���Oi%^���r����B�Q�(�:�e��:v�ŷ1nw�Fǆ�gZ���}��6���׏R��{T6%�%�Vl���~c*s^r��z G�4���٬�C2kݻ7�J�����8~���)� "�Ⳝ7ᘩ���6�F�#��i�ge�.D�lm�{�����ZZ��m��6L�gB�Ʉ�<�@x�����X��ֆX�����i��}3�y�d�q�r��n3Te�+j!�6�r�RXKH8��c�=[,kW0X��r4�e�:@=h8�� ������M�µ��lD^�Nt��8���(�<�kL;�RP��־G�)�&��:�p�̩b�����i���{ν���w���Tg����0�Sz�\`H8��M@8ɨW@>���c�GO4oϟ^�s8�%2���ZR2*@'&|HZ�[�~ܻ31�6�o	��`T�_�F�qm���^�y�W+�ř��y��j���97Z�ރC؇l5�`0�!\�W��*+�P톲|՚w 3!�������[��P�o�&ل��K�
����Ӊ3�|����SVy?���*vv��e���b��¬0`�Яs�И.Ú@)��<#u0�s�j��:��������g8զ��c�����f�r=I�=Z�͏���j�vM�Y�0[ռ6�uV�������H�����v"�<�c��A�M�M�ne�+�%t�s�ե�}y��9�7gt�(SМ7f��ÿ��Р��4�� �l�����+��.z���j���E��o�o�2�y���}Gf��B:�+۱�gcť��������Gs���S��!��O�]~9���a���D�z�R�,���%t��ɥ��f���;�g�0��,���1������)�j���}�!�	��9%�\c�����O����A��X��=�2j1��\�<�����1�X�{(�&����_<I���T��+�^��͑Y��H��L�%'#:�ӧ�ԯcYݩ�\L��,;�Y[����, ;�t�ž�pM�}�@��Q+�.���5�� :v�󡩦�����Ջ;�慌P�Ya�"l�2��%\d' y�� �o{��UV*瓉G!a����|+�L3���oLs��y.�1��G��ֆ�y�>0���'�~�X��qwov!�Y�������%��`KO�cy���2kH�dp��Ɖl�w�:9�i�-�YX��!CEC<cA�<�'M���}h�̵8�<�/�ѭ	�Y���.A��6o/7W�
֩O�8�$L/�wˍh�A��Ϫ�ϩ!<(�����P���{"�P�C�`=ʪ�%�ߘ���vl�}.���V�^�v	,ݧt���I[��zK�k8s�B�L�{�����U:�Z��@�����D�S�~��m%����X	`�ff���sG;1kW�������1������9�gO\��z�G5��1<m���KUv�R�<�DL[~�c�Jo!>��$������J*�U��B����؎���OY����
r?���ə�Q��0�������<�7ί�d?�c6灝���+��u�=��r.w�j#���Uf♥��E=0I��8�C)~��٥Mcs��"Nej_�Yv3y|���]on�'n�+e�A��\$E�!9g�4B���8�����,]� �a��4�����S��%;;����Zʔ޾�]X�1�N�NU��A��>�/�-C�� �+�E�	��F�����(�)��2	2a����xyUP/��h��M��i�ڦ�C?e��Mr=�0>B�A_�ߖ�ve<,����E
겵Y=b�r���Ϧ9�=�� ��~[�6�T�8�Y(V�D~�AA�֠�G��V��ư&�A��[��N�Z�R�ZGC����O��|z��]b����+�X��|��-pع�'��a�(�7���d!��W�G��qA��~N ��\��)�H�r�٩̈����]ʃ�_O6�Cuם�n<1u�4d�y�)���q|�Jm�S��a�Y�ge��{^�s��3|��*/^��2��6��c�z�e�>�mO0���Qއ��R!sv�XH���Ϯ�!�3C%��:j$�������դ�y�9�l.u�]�Klz���7`�����B�Z�z����X3G�#K��jv�����GYp��u�hB������cp c��}�S�����tWʀ�w�<�����oWm����	�e^l�MWS����<�j��-lU@m�Mt4�Zu�j�;$;9s��N·�Wr�)M=��|HWPU���ެ��h�2��w��|�<����M�rW��;�!՞�����~5���lײ�*�3�y�^�/5� ��gz]��z����{us�M(�e.�!��!*�ih������dח�7�'��?� B� �0�1�I�dp׿�]������t}�R�5�{>w�ioe^K�/8��m���qL�MQe��t?L�c��x���<B���t!���e���3�)̟~[d%�������XN�1T����A-��]��m���f%��8u< ��Ҋ�WmF�Uo�D��Oe��cu��>ٞ,M�na"O��7W&���Sn���a#fϨ'Oɪ�w�/4�-?��WL��}խk˦7���y�&Bm����,W��(�����L�J�'�'mZ����m�7'6��`;\QW����W���Sn�b��bU�ң�e^]5�وz��6���T��ET1U��N;6��ۏE@-��<�X`ޙL�)�Z�nM��Kv݇?.N'z�]�.��c[0;�B؁%�]�Y�M�j��،�����]0ЕJn�;0�qخ]��R���Ԣ�c<\[H�l0�f���A�m8L��C��0�|�܃'YWZ�����;�HQ�]>�'Ʊ���^J��R�>��Z��z�?�#Ɋ)��G�CІ0�<��V���M��E�Z��a��F����t�u�5 WA7L��6V�n�!��흱��i���+��O�R�ĳr��T{�i�� �1���{�3k|q����H��!���h�p�8�=��s*��l��=MM�e��a�8�$�,�30r�	�F�}x�Q������N��96"DFPm� (�MI�P��M0
o�7��hE�Wd��u����v?Q�]�˒o[?�������c#I�Z﹗��u���e7�%��vy���u�n[
hdell�x hg-S��ۘ���+o�삿Gp�����CD���%��M�,γ�+��	�N���r"11�M��=�b��ؘ1jv�^ld�d<������=c�y��� >B/w�=Fװ\/��ٔ�������w˿{:2�z���'�ZS�d��o�BB�/��w���c��L�!���Z���V��<{���jp�dE���흏 3dP��5.Q^�f�<[��^�Y����-;C-�s"���������KL�L�7ɔ,	�~<Z�����m��*'��5�p�[�V�yk�����:�!�a�am%[Hy�:~fmZ��{���,�+ݯXZ�O؇�w�)��A.K�e�l)��x�	;s�xl�R�zxA�k��ΰ�z�m]�+�ٵן��{�-W適�\%���n��VbY6y�U0�s�+�jo�����O��j�.�Ƹ���{|�ո.�T�5��e�%kk�+���{˨;������<1)�Q}��T�Sk��ȃ� r��u�U�M�K�)ufcg�#Nɣ7��6�U�)�+�w(���O�<+��xN�|�\3>�퉙�q�3�j��>����؇�bS���8s�.��,��G��\U(	�ԶGW<,zބ˙�pQl���}�Vd޲���o�6'��k��CWw���h\�x�_��>L@����A�#Q��$d��Ml3]Zq�w�;��:���Z�m�н��l3���'e�6=S�{a�T�Hs�k�TGD�{���k�ږb9Hf�ݘl���b�����Ui�n��5�ۆ:�_SF7�gc���H�ƾ�=�򷞥�1kgle�4�E@ޘZ���>K�!��.�˻�f�j���\�����n��e}�"��c�"Ԋn`7��)�X$�dKǫ��X��|�����������o>�U���>V����Z�DO?��E?/�(x���l�9�.F3��M[q����~���M�6�{?{��3�5K�v/�[1�W����a���ĸ�b�='��>[.��zTf<��qq]�"���u�5X��b����~[�D�>O�Fyg�'�_�u��㌵���1
+��^�Ae�{��� �,2�l����1OY���pk����������#�U4h?�
��Q�款h�]H�P,jr�&Z���Wm�t�Px����l��&������T��#!�W�E�w�>������z����n��}��2�Vr��2��XB��d���]�p<톌��s�����7�����0��7��s�^���ać��/}�m�����L �����<���v�MN���ڊ�|s��3^@�*KxH��c�~�����}�Z��~1c��f�J�rZ+2��=����F��r�G�tH��w�	�)���+f!f��/��?5��e��dX��vD<���ԡ���ۥ>�Չ�7�)�c ��xU��b��R��BP���i��J�v6^�R����D4ӤZm�+5M��з%��uC�{Y��޶��a� s�T�=1�ܜ+s�Z�����qCZO��-An���8�c�Sx��bnnf����E��{h``Ӎ.k_�0���#2�wa�ڦ�!�Y�N�6���;ҩ6�^El��}�g�J�]C��M����А���ٴk�0���S��[{rB��(:���'��m�s�G����+7���j���W�e'O.��D�c��.{d�z���S	���]��Ǯ���R��^\�9�q���j��l(l^���(�78�]b���OT!��e���@����_�]�Y�C����}ړ^�Oϵ,�����Zip˄~����㨘�oG�=L�B ��6�r�(u�/j��K�Fμה�lL����"{��G4�[f�n��.�ά�R�ފ��SO+��5��F�y8��/6[�}Af�w�߇}�{��a�o ��|��H��}�l>	�G<by���)����>���kuLGL�)��Q�Lã�7���Y�wGYi5�҆�35/h���X��nq����F�vm�q������:�#�-�;�� ��w�%�RW����@�<ޜ��8�=�{� =H�CZA1V<:���ܱN����?u�d���3 Aƾ�� $G6��[�Q� >����-z	�ѯS�#�����s�C�gd��s�֭b�ND;kǝ)
3���>0����EK���+�����)?9s���Ct.������w���@��u��o����|�	��ʆ#�9d[��-��k^���N�s��O^�yR�u��M�3��PO��L������<$,vww�nJ���$��_+jCQ�\I]v��M�fC��C��kĴ���p����FE/����P���0��ܵ��;o�6v�������nק�D&��y�A=���j:x{��{��(ߋ&4���ۄ����WB����(q-R`n���i�%�ۊX�zf�v6��*͋�YS������0/dﭣ�����Y�rb㹺Ї��F��Q��w��H��r ���>���8���Wlgs�),U��l�펯��-�:���(ꤝ��]�;�L،�9�w����v��a
X�n%52�,M�OB���R�����蕑ƲGD�uيn?�eVpJ�;e]Ʉau���qՓ_I]�9�4j�/�v�7űZ XW蒛N9*g^R��K�X`�.U���i]kneΗx��;0�mdk��X"��ջ��Of��V�7�b�E�yV��j>�Ɗ��r$sޏqv�+�}�U����t��\��\�^��X*+��-q,�KhP�(���R�חi��WS����V�F�v��[��X���-G�g���vH������WiA���ɣL=��4��F�}R�,�iSy1k7.T�6�-
��\�]��j���s����ˮ�r��x'�i��*��S������(�a/M.fR#p�[o_f<�il�{l8�
í�����Ʌ���Y2ݳ"{���75Xz���A��^�
D%��u+�c���뼚SzmI4Vf��U���ۨ��^�P���1)\�w�f}���oc�]Hg����9���P�Z��Ԝ�v$|��U�4'VG�zV
ޝC�vrl����=���ӹ�:���2���`�,)D�J�K{Bl=�v]hJY���^m�P��ZK��Z	Z�h(࠸ZH=�o�����Խ�x��״�ud��c�"�B����/���n���T'��ڑ��^ي��R��KǕb�ই�ؑ�Ë��o�},�a�ٕ~��T	�2��F̮<�ݗ�vñf�~�z���E��ɒv�2F���(�^Ե�B^�68rw����q1��^iN�ja��3��W�+�樌z�3G�b&C/���u�z�P׬��8�2�^7(
{�)���ۡz�U���*�g9�:
�y�z�QXq�z����&^�ZWe�f��BTj�kpnj�Vq�o3]7���m"Ļg�o3g5�mX��r;�)[�f`jk�8$�3(u�8�V��V�r=��e��R�#�H=�D�ZbS
KS���p�5��v���ZR��M|�2���k��1n��1�c.�;�S�%�oN�Ե�)M�<�_*3&:�`����GU�u�ڍU�b�F��}�N�+Lo+8���������̤���Y)*�`܃Kݨ3Fac7���v��}Ϫ�p\�9���@)<Ҕ��o��\���+�.�❉ƆX�m/2��ra��E�*�S�e����l�-�Fsz�Q�R�iۍ��+����r�Ê������+��^oYz�
��"�,WP����ݶ���U4�ऻT���d�0���Krt7�F�uڰͪXyw�]]���w~�A�)��)��7��U4d��K�}a��d�uPS@j3���ǧ������U��	�"�F��lօ2bi�Y�Ʈf:���Z�,�/��t��}~?�(*����s ��	�����R��dȠ�N��ImӧOn��s�3 �(=,�(r$�d����r����n�]���sB�"y9)GP�U]:qӷ�nݾ	�4���4	��>��}i^��QZ�r4��Oonݻ|{��ƥ��C#R���Z�2��|q�N�_�ߏ~/w%�Q����p�B�t���Ǐ>�B�>K�k��i�59 r�R@( �^G��|�{�M�H�7H2O�I¤��@1r7 $�r�$��(���l�e������׍l��M��^��yM޼�4wb�o�$vP�p���>�4+tF#��
:������$ʊP�	��B�`��f$�e6��(��"�FB�!�� ��Q@S%2l�\e&-0�$��5�&�D�m$�1��߼�K��K�`^RŐ�
�:����ǆ/"�h�C-��D6cݥ�&j��*6c]�������ze2X�S.{l50}��^X��0t�;OGZ��@�̘y�ީB Z�u� ��]"�οy��#$>cjhg�����U�v��,�6��Z�Ob5<53�S��mz��5�@yA9�ڛ۵��p�a'b}�|
�ǔ+~nU����0&!>�s��*��R�<F�[��C��-��SM^�⧓�}k:9�n��ۚ��;�l�(mpf�����2��fqӰ@DW��2�[��D���-B�u $�ܲS4���!�bu�c�AKt5��L���t�'��π��'�6�t��޼l������9~v�&q�hFj��8�^m�=� ��1c#&C�	ךxO�nl/m)���"9E�G��mƦ�s`�3T�ܴ��g`�*P��g���Z�h�i���F���1�g�q��3�F��Fk���~��{H�@�s�>ƗD���/F"�Cw��a�ϦßK�&�~Ţ��[�˞��3�D��>��:I�%���=����x�Y1X�.�����0��)��c���dvE��ۅ��ht���\y�i�IhB�#���e�e���8(�ըQF8b-�]Tx�e_<3����!}ܸ��j
͊��i�6U_���]}|>���m�)Kbf�;>�ml�e � ��u�x�����!A}q~\ZZq&r��l������]�|�O=�e���+��n�^��M��Y�am>*�F�^�t噻���(wV�S��Nh;=҄�O�)�:�K��4��=�ϟ���b�[ʓ7=�^�k�r� �X�M�O}ˆI��A=;�z���H���4�h'V�n� Z��&��9R)6�b�޶���f��7/r�Xf԰�j�#��\�c&�_�&�j�u��2��yZC��W���}�Ȧ�*�p1�;��ò�q�)��AS�lnD���*�b�Ƹ���-��l�wfT�%ra�xɕ�`�LM�mՓL5�ܮr^�ǪY�*G��tF�������7K-�Mo��f�S}a�i�����s�w*�jjF�7"�Gl̨/�F��_.�%�����w��c�&�a�=g�O��W9��<�E����G(m�؅G��z�˻:g���3*m��hoc�Y!P��������\��Cmtw=�Bd�2yШ�*�MSK���|���7Ѥ�݉w�/��=���=�C�Yi���ƺ��T����yV&od�
��N���@�x��b�I�9bYt�T+��#G�����Ň3��:��{(Vx���Z�-ӛ�Yw4���s�,�<12��||�����W�����~Yh�O�68f�̞�`��9��S���Cƴ�xB��qSM�z�Fܛ�ʫ�����u:+���9�����/C��p�ε�T*��{פ�NS=�C���m�(�T��_��W��M>3,}uf{�����������n�6�t��혥�u�[g3v{%��y�����>���4�1�2��༈|��;�@����c�xY���ۧ�__�|�lj|i��6�������Ăd�{ ���L�1l��T�5R�1:�b��]\���1��������g�W���:�DL�D^�wB�Ι���ћ��6�e2f�@�1V���fp

_X?w��q�[K�~/�,}��K�u=x$1co��^���1s��p�7�y��Z�ڑ�-���`���$ͻ���xsB��?~�)�>����* �b��W	���ě���v��<ι��&ҮKVkU�(��Mg��#�
�B�����\��N�ݗ.n�yV�k�Ӌ��N/i�Z�Y1ע򟵲�b)�qv#�0���S[8>�y�v<�.g���4K���F�����������z��0���R�Į�i��(�UU�&!z�K.��ꡯZHzd-H��|H[ñ��=�U���af�)�+=f�I��,�10�+Ip���<�2���iS^�)�Ҧ裸-N2����x�K��f��w�Y�4�2�����nf�ɷ�rèoD��T�q��`�{Y"y\��WHZ2�3slI�l�X��Op f��xnNP�4Yxϊ���j�=��e���s�َ�	�lm[�\+�����9�������5Vj�7\�=n�=},w�0���^n��4��Z�ޮ����[�)X�C�;`���vo7C:mـ�y�c�y��"�P�u�[ǲ��k�8٢��	������C��_��MD^���~Kߗk2OEoS���h�F�K^γ"T�%��8�a��s�&rÆ!s��ͽ��A!<WM�_~O�
z8i�.�o��QU�%��rz����FO7�؊��9���X.`CA1l��]�k{�6��S.Ɋe�ϙ�!����Њ�v�a0�йG�*����X���ϗKg�1s��ieө��ݛ�����
���d3zh�k��-Y�"?�,+=�HQ�r���!����;����(c�:��W%(52�������@��3��@L}�V#�o�cEx	Xm�M�~��i�vi��3;���F��q�+w��>�N�ǰ���5&���V��^��nm�Y(��
4I)�:&�k'v�����c���J�{�n�e(6���H�r��4�n��Z��0r9gGIR��|��뿪�~Dx��D���BQ=�?}����&���G�"D0a2"_ʋ�|�e{��a~taV>�Y_�tk� #��o��~��*,�6R��^y��A��� 
Kd<;[�t>��A-#5E;��\]C�؞�m�Θ��V�F���T�%n��G�K�jqB%���դBh�6+.�ׯ�'�Vݔo�IA�yv%�����~Y����PZq-S���3zu4���,^���[eV7��W��g�i/|q��/6��̧Q~D�&�RB� �A�|��Ҹ�����64-��?Ҭr� _�~]ٖ_7����[;*m��Q���W�梃��QA�&Z�1�4["�A��i�arNK�<�:6He����H��m�4�VgP'�Z�Oe�5H��X�{���WɧNc1���6Fc��݊�L�����w�s���^Sy���T+~n5�<zmy��=)~:^��{����m�F�/%s�<_��Y��W�Q ���L�����Pu�*�쟙ax��!L[s�w�M�r9�0t-��@�-����kwM��n��qH�����p�D��[N��db��.�I����%T���hl��x�����nV�+6�!fU5���<Q��u5wU�j�[h��`w\?��P�~~��Z9�c�J��=ޅV^=
��<{ڃ}��R�LJP���Kq�,mG���I�vԙi>6Zwa�>�朚C3���~��7�zWά=��_����xh�M���ϝ��Ĩm��lU���מ01��i�Fc����O �����������ɞ9�ъ��{��=��U��t�gm�'�<b��D}�@��=`oT-q���L����'���S4��1c\e��X�����c�5;�����5��s��@��z�?7��"x2ʈT�K�}�X�UT5Z�;}u\ �%5�c�:�`�	�pb��K��5�`�t�3ءS����t�]�n����:�\���ɰÛ1ݬg�E�e^&]���⵬=�G������)�¯>��~��A���?o�&'��(�]��邝�|��̗��)�^��%�cW6�s����r�f����*-�&�[�k�3X��.}p)�;�8�e�Y�m�۱a�L������f^�n���MMkI۶�r��b����p��O0��,nC5G@�Py��H�Z�#�1<��{W'[p��K��{���kdSm7�eF46���V���v�)ç�{����W�ü�{h�T�v�\�-�GN²�h���:�㨤0��[s+���5uĉ5} V�P��;���c��x�x���[:�%0�5c3��X�co�I:��4g]=�Z>�]\�17����BZ��Vl�����������p��U�,5���wA.(%5��}*1�ߖн��l5���fŃd0c^��=0בz���S�к���"*�y ��fO�q��`3PħO���J��}�P�R7Cl�e�ݦ�Іz־��!��!(Gs��f��(�%�Y0��"w�W9��<�G)�m�YM���D��7r��k���?/8MO#�^8ɸ���"�	iѼ�}r�6�^[)��r�/Eg��d^��z˫"��Q$�`΍y��ǝcD��ߺ[�� zCC�����z�����@ьdR�,!;�*J��֭�geU?�0tL�G=[>�1ͿcT�=�Z��I�������O�=�ѕ
m�=�q��BI@��.�f���d�}U��vWʾD$�N���=q�gZu�n�|�r�P��B��da��/�(PރoD�0ʃ6\�|cAvn� �LZ���]ح�6$1Ο`;D(��!��vk.k#�3�hn/�W��ܖ�R�����@�!Π����w�Ɩt����l���xŴBgy������_���Fy��דJlD:iߘ�(����+�Z��j�!�:�I��f���b��&K}I*>cS5^�)���tw+n�y`���x2��F�KzM�9ʍ�Rk�2-u���4��Kj��0��uz�q��2�������B���K+'*|�m�^����o ������IH�N����{KK����p|�@�|�-�x@�g�����TE[u:Ș<`]�~���<&��wE����l�j�p��B{�X��߂����BW����u,���_����e�����a�	>��J�����)z�	��U�y�,U�(���@O���f����W� ��=}�n���|N��@ׂ��{	�=�1I�����DD;�x�Q��f�CxO�d;j�6R�.Y�K)���!sx����\Yr�J1�f�H�锟R�-�߅����7���K�~�6)Gt�T�L�Ĳ~�fl�m��:dk$ �-@f��&_=cjy �^YoGs%��g�b��������Ӗ9<N���C�w��tۯB_�.z�M�&
�X@E0�܁ZӰ����Y��5@Tu�m���I�Q�5V(��"�P�~;ʽ�|�}�~�T���f��k�~ͧ�#�c��j�`�����|���GMrԑL?���6���֍�L\ �w������_m�UQW�b�qq@�:y�댿#%����hg2WA�/���&��������W�l��..վ�ٻ�fKcr[|���k�P��5�Gyy;��.޷ۈ����!G�et�$Q�P@��Y¢²c�clմ�ܛ[\{Nv"��j=Y��x�r�Q�w�izF�=³tP��l�%������>o ���cK\C�@u�������L�2�)����h6�m�A��b��0��OB^@m|�oa*E�3ϑ@��&���3�$n��I�=�'�=�-�=2���1m��^�%�t��kWu�2iT_�~EVU�|Ez�� �ݎ�qت	%s��U�yL���s��8Șk���6������9��dX6{/��m # �C]��Q�}���M:=٥u&ff�nβY�y�]To��#��DB�N"�s�;7���o%�IGov]i�I����6�=�w�~� ��¿)ѬS[���C"�^��mD�2�=�Lsxj���ܱ��j��/=�m�<�t�'f��Ķm\G��(�n�TȜtZP����-U1M��=>�-��EH��n�c���^�	׹%�*p�teJ�x]���Rq�Y;�sO�s͵�)s�iP��p��1,�ʬ`ʹ��٘�7��������Ȯ%h'w�?��cH� {�7h�h�[�]�~ 1_��r ޑ2ܷ<̶rڢx�fB���ZغKoz�{�����l�@���t"�e��#  ��k�4�w�w��:a^�N��f������ΕU��S�n����ڎ5�:QQ�NOR�W���v�WG�s3xsu�Oe=Q�P(���Hx�@�=�'K4\���׌�P��䮼ӺV�r\(���@\�v��2��/�������nT�{����9x�3x��{,�]4�?�؉���]&�i�iM���dYW�>C���ߧ���a�x���ƥ�u��5}�������s�j<��lyOl�Q��
���~U��m��<g][�Ø��Ԟ����0]��륭���;�<ޟ_#B(qU��Σ�m���k�%�53s_���<r.��5[�?[t�A�C!x@m�	{�Q)�DAn˩p%�,Ȗ����x�b�	G7-����"��D��gl�.	����1�q��ǅ������_�OM�>�ɦ��e�k:n[�du�h�9����y۬�0H�H8wZށC���3�>[��(��?�e����=�&�XiUg���Ϩ�Xï��oFZ�|��G���B8���{TU��J}y�����s��-cj��-�l1�]'�zFP36^�Jff���m�Q=gXGQ�_�i�K;��;�~��YK�Ϣ��G�>��^�Y#[��� �#���6\S���'�}i��[l�CeI�d������	*D�&-��O��ٚ���]2��Y�����;��> x.fN�#ߚ�{�Z6��yٺ���i7gFE�ou�5:;��l���V�gB���m^��n
י�q��.$��[�a���~:3�5��R����V��Pnxf��qɍ��׹�+�X�S�H�V阻���)��+>6��S���J̺i�S@�F�Ǫ뀢���W���+��9m5�=Φ��戃u�X�Uw={6�[�-�<�A!���R�{U�g=D��n��@����A����U�}	7ȝh9�`y���=].�#�fnQ���s���ԃq���;\���W���2%��IM������Y`}c'�kEpyp�;���KJꭽ�rVu��S5_�����d��̈A(�v�K�t�ժ�����WN̉�U���m��ɚ|;{��(�'T+�(��Jz���[u�ܹZ�rA������m��~r*ݭ�u�ej��t��W0�}G!�4���__|Ta��Ğ��;��=�5ڔ� �/`���4۶/��	�/IkkMw#H+��OZ�i����X�y��껚�fJ�k�)>�� z:v����!��Kp���7Z�N��;e-�Fne�_k)u�]ԛV&S���j`+T��;��kZ���٥h��?5�Ն2J�A�s�X֮HV{f9�V�G>���V�I�=��!4C^~/0E����C*�e��K��V�J�LV���=4�%�Fʴ��vcx/j�Z4���:�p6��͞�L��Yxا+2�v��(�� �
(�-�Gb�A�=��c���t��A����F`��
�)v�]9A�>���oEA�6]5�&
@�8��Y'N[y,;T#X&��{i�W��o�H�(�癤��X�$� M�J�wFM.�7B��J��D�;�-]-X������qA_��I3e��4���ʎP�����#�}�n��Hu�r�Y�CR��iȭ�X����/���y8�Ou����՜���_-��[��߻npi���0�(���{�wMtDs)��*=���{vV���ն����ԡ�urb�*�ngh�ռ*����N�%:h���9�2�w�8}�]�j㏐}C�h�}��� �ʰ���.�l��׈-5ES��W��3sys�7��@�k�$q���S"�li�3�e.I���{d�L�����5����P3�/Zdʳ�E��7R��ӷ�ɱV5ʌ�4 �,ɱ|k���+�<���.bΗ!�n<ާݡ�o\����;p����B�
�/��o/0s9�y!���fA2�'�h�Y�N��Y�D� �'�JǸ��Gows�¶��U�|"N�5.�=�-�kْ0B]M��t�wKv���T�%X�[y�'�.��2M��Ǿ4�E�'�#��#.��K�ԙ���ǧ��o����Gi���ݐ�J9ORj\{q��۷n��1�CP9���@�RRdd�d�ӎ��ݻv��G�e�{?X=A�vHv@eKT�9!�S#�rG�9��+��枝=�><}v��Ҵ����'������˨��z�b�58㧷�nݾ"u������1���fM)��}b���=����۷o�E4�u.���rZB�/pL�!�_�<zq��㷏})<�u� ��5�R���:��ێ:z{v�����=�@n@�(u���M]K�>By:�O%�7&OQ쎡uUx�S�{E�S�%uU��Z7<����<�Sc��ܖ�l=�6��o0hp��Z���:��ۻ�w�9�s���}/�f���g����}|)-_/��Bbj�����o��)����~:�O��#�}��'S�/aRK;Zk����P�^�vz-�'��={hr�U��@L	���W"S�v-��%�j跢�W�jeh���j!�BYB���xm)tHw��nD����(	��h���,��v�/���j�>�ΨL�����ʃu�n����Tk;E\;.�4y��)��`>fJy���׵�b,��Ȋ ��lz��������+����,D�V��ܥk��յ�9�yem=��3��@;g�u|�Ɗ��>nv�X.4�є�kZ���\��OU�P�F��T�,���D��鬋��|��(; ����a)�>K��.��ɍ�>�6g�:u�]��y}�|�S��(>qz*���(lۏp�e�� ����1����~=��j���M{�����$�KNnȼ[�jc��/�BƉl�5�A�����	!~[� 
|�}l��N���s��5J�S���E<�J�u�Wd�*��]wӏؔ^�pG��"^��\d垻�IՍX�o-�E�Ǜ��jhԘ�v���1�Ӡ/��P1��{ˡ�	^�?$f�׏�j�e�vu�M��Z�
�����xe����#��\&�L�k$��(����˳�t����{�Sk���������������L�o�3����}|���}�Z�I�O�P��)�Y\j �H��j��9z�6�;������[;��)?Ig�.�;�~}���Ӈ�jF7>�@oA���*�q@�	9���O~��o�ϱpU�HH)�_����?�C���0��6z_��鏠�:����UXb���ً���D]FT�f5�wX��o�������L�Bj�~V���@��q�SY�j)�c��u~�V�],vL��~�	m~�9��o�S�W�j��Q�X�
qm��������vi^,~�L��ȟCv�C358cf5H�-%=���'Ѭ_S~���"W�1��~��Ӵ{��ޡ���K�oB�81��0�J�޼�8��<��a��wo;����ڏDB���ih����_���K�t-k�g�=�Ly�1I�����f��ݗahSm�,��o�D�N���ؔ9�Qm"y��9foJ{ca��z�tO�'�	K0I�X�9�&�E4�Ŧoy�S9/B��4��\��8�Yud�^x���%AקٞOT�*���	��|�g[��TU.z��Y��r��v)���u6����}�>O2�n��|���".JjfT���ϲ|v���׵�FG�{�d�������=sU�G�e�:Ѳ��E!�V���]�b�"yl�P��qF-S�Չ�k�ۭw�l���1��e����Q��,9�~�p_�ݓ^�����R	�I��2E��0����m��b��,t=tG0�}�=�z]2��/��>6��5!�,����0�vnI�E��S����Jm���+W�T� �G��_`�n�33ߢZ��L�b8f�tj�}΀��qq\mP�����˿O��&~tt׹M!����������G#�}!����2~5��3�[cqW3`OIGs�����F� ��մ�}Ȫ:�fTRc��C!����9���&c��C+��oN"�|�~����7��Z2u�c����z�f����XC��"i�s@JC�l&Z��i�L(Ɛ���X�	�����oXۦ��If�E�0,�������؞}�~y�P����%۟XM�E��Q��$�:R5<��n�t�@�p	f^�TY��� ���˿����S��N�'�j�)����nm*���ڱ������Y;�Z#��)�(�o��)����)�9���*�M��2�uyg\��ȹ�
E\zE�-McpcG��C�\9���e"&eF_}����|7������&¡�k��T���nֹ/����/Ǽh�ߡpxkvw��v�(�.oE���Ri��{3��aև)��wo���j;�/^KLNT;]��A�)�_d�32l����c��أ�)l��{����o�)�t���sX��i�[��[��W)c�g�֘�:��4Dò;j�D&�0f�t+�Ս"����	7�"v٪��u3�Jj '�t���v�Jm�KT�����O��B�)����F%�H<�z:�e�43+�L���Ӭoj�7�.�vċ�#t�% #|d���I������arS�[&K#oQՍ[���^��QL��#�m֪q����`^;��a�@sƺ1�тւ�s���i�묅_����HIF��xN��@J�6�G�m��caF6E)�q��ؓG�R$ِ�����v�8�5�ezd;zF�q�c����Tsu�c�Z����6�	�y�~�w��Ww����ٝП6 A~h�b�o�)O7��ĸ�*t�p�G2���^J-�����h�ʲj�zұk�Ћ��|��?P!~+�@k���@!�?8-t�_8N��J9�gEV>�Y7�U��t���L�A@f�C@r�"�p,K�:j���|薿b��
�j��d�5�}f�ucE�>f�=8�	 ����@�g�����^~׶�{�uɣb�N?��cO���P�URɃv�q����ڭ�T��vR��205m��0�v���7A�H�.]@�����R`�݄W:*��I�m���b.��
�&�M�9g:�U+����Fs]�Z�[�{����׻9����i�k��p�`�of��k�C���^����[Wk
��1���R�W�M"u�����@{4a�K�1sf�1��g�wݯ�=�����GHn�m�A�	p	�b��"�CwvÂ���eN�\a��K����ֈ:���� ��W��#�vl98�f�H�k�Z{�
�o�W��\��ܴۘ1ڜ��uP�d����P�]��˞Ę,��ܳ�>�w�,��e\e�[�K�����͈������T��;O�H%���R�(�o�'�S�6�O���/7ҵ��d��ۛ��'�s��ֽ�&��J1o>�{.���*E=İ�`iy���z�Bj��s{\����<��4773�j�s-���
��?�y?\�%f��ń��R��SP����щ�ɭ�#P�:�(a=���9ΊO���^*o{�C����Ph���	���*z�k4��B�>~tb�H�S��B�I�w/-�{K*�krS\��w���*�{7,�X�>��|\ iO��6>��}��%:�`r0Z�ޤ�%H�`<(Eڨ��Bnع9��SwΤ�b�Wj��pu��G����8	��;-�{m�/�7��3�XI C��/v��r��J�cx%�e�f��}|�9��*���j����Y��N]:��%t�P<#Q��1�U��\ڂq#���x9��:�{�����}���0�I��c1�d:�y��|�x3�9A�O�/�����fo3�z)����Ss&��h�R0oT����%R�0�Π��k</ot~l\�X�46�������d'��^��H�y���Y�Z�v���\r�H��q�àU�d�Q��g�y���(kăkk��#���G��A�a���Q�~�U4���R*�m��e���o©Q�ߏ���@��ŀV������u������������X�L_�='��4+\��d[ogO�a��%�ܷc�`�xRTvCj�tӶ"$j���_����1l#���o�}����t������@GO�Y2`�c�:���9�vc���8�|{�!�)���Y���z
�A�2P:�|��rgԺt�S@4�N��!���\�2zg���w�[@�|Ğ��V@��>���v�y������ai�7!*��̻�����-� ���M�����9�Ԣa�^^��f�~U�гj�V�g3\�5��N���|ւ�v�S��~.�w8Mdj�wyFm�y��<:�ϣH��/����f��n�ޤ�^B��,��{��Ŏ[\��쮭�Qe��R�%��u,v�D��,d��H"	�V�f��t�nR�h������G�e�ۭ��l�j��zFA�Uf�KqlP��׼�w��7�:�=�}��L������GN�H*D�mx�"�7�׏�V_!$�,�"DI"\^M �)��8�Kĥ�ӹ�n ?���s�*��.��?�{�^{VF��Ț�P��r��:8��gK#ZeSr�9/�|�%�}�^SU�{�I��=�)?Xr���Sx���m��vz�b�5T�`�÷��������r̪5���#z!'�*|����Gi�fN��r7b���7k=k�����
?��܃�]��/ؠ��A���.�)���5e�J)��bS�H卿I�Ɋ�O!��C�4��:���*J	��>q������yl�	�R[��jSm�TX�P�Ā�9��FEs�w,鴧0�&������-��}h/\`Q}�qXޮaaR4YO����tp֮I��_NY*�������B�|}Ύ;�vS\H��.o���
�\Q�t�(�q����ֱr�sk� ~�����ە�,jR&�H���bC��Ϭ��.z��/R���9�c��f{���(�Q�jjsf�Q�Y���q�&o�����vp�|x�-X}�
�@ߵ�d� Y��69N3)GC��p�ZD�!��؛cL��io�zQ���s�lY���k�ڥE�oS��"����R�{j�{�ӊ�~^ȊX<=������|��@y<���p���NVb���+���ё7sgƛ��̹�4:��P�)��k�����r�����������>o0o0a�o8�=2���h�M����I��`��@�P/ߠ��|����X{dL��Y=�3/�s�t��O�5��y�����&>���A}p�����0"�*p��j��V��yU��OGY�]k�qv���^�C�&5�"E���5��`�������\���}%C׏�x~>����"^�,�`��C�[�v�Q��{ ���c�Y�w8n���p��;�h��m��ı�Κ���< ÚtTSrQ�/��\d&�n�c�^�Q����h���A���(�X�D��|fڄ8����4(SM^�R��*cKhW��K�}�؉;G�uy�_�T�,o��̟T��i�7�"B�">�)@M�A͛���/�V�r޺E�L�7nj�s�ylЕ�0��2b��pV��֡4k�;��߀�+�.$��7(u��a���� t�s�tU)��%V�B��i1p�Ņ4o�퉍���!y�{�*3?=�Nw��G`��C\wH~P��>z<Y��w��徶'��*N>��R��0�gщ�0���mfչSS���f;��g�۞1P>?;
�������!��!e�.��t�}�s��(�ZY̫6�=�`�Uv&��P6�����T�l=�w2	�3�o"D��n[�5ݷ�t;��ܢ��:�sa���O�N���^y�[��׿^���C��1���6���)�M�-l
P"AJ���5��S2�$w?Yt����p�F�c"K,kd9˾ȓ#��s��K�0wpoeL��Z�L�5��;aI��b���rĿf�5v�a�Cvl%04@����u}����Na��?&_)�4���辐)��<pi�@�&��t����ƿ|�����ʞ�g|.	ȃ�R��{ʎ��~.���C-��L�O�}��c��m�!���~z���8�7�:��U/q���� Z�}Dl����s�S����4M-���k��Xz�6 u�8h-}�}����&"�C	؇l-�w�t�Y�5T�գxb��;>t$c�;6Q����R2�`����ګ!�K6�"��MqD3'.��%�~�
��U���g�^Oqwq��+�������r� ؀�	��LÙ�����띛T��:�F*b�Eߋ��v�� H0
��_��)u��6���j��^f�Hg���S1�װ9D��+�a(żG4��|1�>t�[�U�)������h�C��x��3�&r���1Z���J�8���+A��p繗Z��N��0�1��[B�zf,z�j�Nو~�P���y�²��l{��(v�����;�ڗ	��B+rS\�Hb��1=��trq\.��G��C4�����Qp-P��_]���;{q��=5e��I�u�G[�dŨ1,�ϖ	R���pܪh�7#�10�mv��k἗-�i�k.�m��T�P�	��<6u�[�l&<���6��`Kl�����\>����9ъx������7�;9�CH/�$����,h�Ju��>�����1��:%R���S�dVϕ��+���^�W��7�|�y���k�n1�N��n9��6'�lm}�ȯN'�}���W0zNh#�si��-�����Ӱ�`Y��aL.z�70o�k�_|��^Ti�9n�z.p$��܅v�[���X��w�����(��x[5����R��H�u3ع�����F��d�S!����ʂɩ.�b�u�堠��kQ�
�}������g���Ay�4.͈�Q�e�V�	Zg�evN�'�;=u�N3�j������j<~�.6�J��6�k����	p�Ec�y�H� Э�I��n�u�k �Ȍ�j����r�k4�Gk| ���}�ś��X7s�Ͱ���[�9���3���Ћ2'z9.X^o� E������q�uo�/��Lq�A�8-'^��קC�XK/o�;�g*�)�%ÑT��&a9
В���I�@f��g��J�|���2�U��8�]8GnV�ǰ�_@��u�N�rX�;��qy�W�:�y�=�um�I�xkM�|պ�<&Z�L��gm��qY7ent��_K�K��i@8k�Sź�ɯ0�`f�=h+KKf��
K�W�_s�r=��
��������^4�TU���5��[�7+$��*�Z�,(�\g+�=�oT�	3�b�ɔ��쩑�Ւz�����b�KSF_IWP����0�,�v�X��(�ˎ�ە���v:�l��P�ӆ��N	s7B�<�o(Ό* 7v6�u��Nb�{�mG3Q��6�u�v���	�F�s�GQG�ݽ���'\���0u`�̒�=
��T�oL�F�F.z�A	)k{gm���ʽgG6�w;��wshq����5��ۉ�.9��;0�#�K8v���[9S���3Ή��f˭a[����Z��n�씹qp�8��TC8�Q��2D_R���w�E�*��dm��n��Ȇ�׆�dWj�2�u�����[Wڵ���fN�QE�ݣ;�t��n����]Q��3�w�E�/T$ڼ2b�;׬ۜo;��҇UѮ�En���ƦN�Oq�n�J�����&�yNVݲ�%��=x��<嗙s���{��6
����|'Vu�Z^���&'r�l������~m�0��z�<��ny��#=}�XOV��ƶˣ�F����I��/�gi��5/���w��]/���M��Y'5ΫǗ}�/�Tn�ҦK�Q��F�(�Q`�݉�N����Fi�V���nh�Ɏ�2`����"�#i6�=�u�cR��hE5�"�V7�}��)��o�1���R��  xJ�-�Ի)��͈n8L��遉]�.�����n���7����0�\!N��[��!mK�pB^n�vt�/f8s_5���G�F�wZ�Y��M��ЧI���}�&�;.�ՠ(�[%��wnb`�ء�;ٖ�.u`�7խJR������8
�J�;��m�
Tko��r�+����6��X[g7�R:8z���ta�S����Љ;e��\�.�S�sҠ�X�p�6�<ȷ�e��at�A�dLr�
TJ������dB6���gE]'���IQ�E�����`(�+�"(aW*�YK'7���;��xHe�|���=�F[�5��2� ���s�����8d��1�A�~2��Y�4��y��{FJ ��ݾ@�lř��˦D6峝�0F-��5�!�����O����B��NUt���v������m���U;L3�*Kѝ�����;vW�,�΋֪=>FZ�����5a��ޗ'#ؙ�u���N��:�P�zq�������ɺ�k� nd�R��:�P�s0z��
�z{{v��簞�9�:�	\�� 5 �r��ӎ�><x���+��'P��uTSԆK�j�\��b�#��+�d7:z}{|x��=�=��L��� RД�@��M�qӷ�nݾ+ԯr�.�)2S�z�����:��r�ێ:|{v����q �@�`Е@+��N�2<�P�m�ǧǷo��� $�.���j"�
\�����=������������2R�oFb�� ���.㾱%;� �ԩ�2˨�
�JJ]@ω6P�,�)��Q5LH�i��i""2�BB�!6�a��� �4BQ2lI�TޒI��&�}��]�s�5��ǰ,�sR�G�Vڳa;�:�Lm�M��u(������U؉�TЯV�|�xeR �m�7$m2�H��4�m6R�&,$����H#$��J�DÉA�a2�"&���Qa�=���Q��%�I1؈�fTA�c�{���%��SM�����UkPЪBbIP>M��r"�cix��$?(����N�)x�G���|�?���M��Z�Fa���4��K D���'JM�-�Uۭ�1��ų��}L�����O�"y�g�+��~�Me@���.���.�'�&d帾~f���5tI�wT:<ڢD<�Ϟ̎�l�V��oC柡����~�Us�Z* ��0�
�W��-���{1�w�|}��dV�*��,=��5\I-�^9xJ	["���vD������ft����	��SRӵ�KZi��Eh�&�s�q�3�w�i{�Rߊ���<��Ex熪����7U@[o�+._n�fYq��ֻ�6���DU,9�~�k�ry��F��wDw5�¦��5�u��9���sۍ��Nʈ�,��-m��(��{�?g��M�l[��l�c~m�����4��X�����7q����$>Ϙ�aY���-Vlvf�v���5��};��}�dֆ�YXwg�w�+<�{/O�g�'.��c��po����a�&��Uz����5��;���"��j�-㗆Z����V��.��}�cBYN̎f�
=a:�OU�
3۽�}R�2,�:m��iIfi�)vR��1�kV-w��h�:��$��� a�9_}�k﩮��F�A��Q�#z���$J0c����v43@�w�}�.%M���e���#-��k�;PP�V%txZS#{���R	�5bQ�[��s��4O�|�㽮*Ύ���o8!3��ThN��&_j��,�,";�V@�=x���i��K�j��{�I�6>6�Eߨ�u�O�L� �QOu*�o�˻��zr������dS��
�Uˑ܉�5�)WD^�������\�%~���H2���@d^^$T�Y��#tk�@��vf�T��-@�^xĶCg%\�v%+���]��6Ԉ�v�0�Im���Rt��w�v���bl�Z��S�S?uy��,�~Gj�a�m6��m�s��vHt�ykFXe��� �ʑU�E��w��ږU�B�CvR�Ο�g�=m3���o���w�4���&�|T
��]Z�w{P(�ک�"*hF6����۫�����r)N��vnP�t5��6b�K�8a������XSm(]K�b��!�H �}��
��-�ҥ�'q��S���T�:�Ax4������T���^]��w�c�=�7o3/~8�������؝O�����Å|G]oZ�)n����E���]]����g�.ޝ��}�Zݷ}������Y9$ՅA&�dM�y��ff�ME
� ��}\��� �s#��dk�%`%K{�������q��Y�2�]S�y�����CrE*�n�ƥӮO��*��R����t�m��$���i��d;��5\-\�롵L`�]>�E��A��ޙ7\Y��0͎��1N�������K3��0}+����WV�u�Y�9�s>:o�����"JYj[E������k.-���몒��ѥÊ{*���5ū)�7.���;�֞���* �^C�G�y��k�+N���7	(U�-��ْ7=D+u�VnQ��;�C�^�8�',81�Q���DGO?8J;vD�a����V��^�� ��zb�O;�RZ�p���"xŰn�؏N��f�E�sW��et��5���Ȱ� �V:ƨ_Jh��`�.��s��CIs�gs��9K;�l7O{�5���Wз�=]�����G��R�;��ٜ����rz����F�=�>�C��/ݩ�%b�m��㝵��W�w�J�mU�S�Y~nD��g�GTQM{�9�in���;�'��qߜp��E'~���de���ْe�n�.��6r*i�7��V͈�Sd5>Ϛ�ɜI� �D�²w����c79����ԍ���/	��T�Q�x����=�e�>z걯X�ڢeM5J1=�x���}ї�dr�
��Vߊ�ܞ���c��}I���sb���� �9�v�����:���tڕ��U�^�Qoi����};�����g�˺�ߺpB��]�9�,If����2��ć��8Uv�֣Hi���N�k���qZZX3���P�����E`�NLB�վ���YC���ݒ!-r4�_��:�{/����[Q;j<�?t�����7o�G��{����fȹ�(Α^��{IB�MF]�Mz�a���4�S��MA:�X�Eu�+�cC���u���T�ȼ}t�X�Q!i�8g��Xeqk��^Pӷ�Op��`Υ��Vm��N��ŻsQްr�+������bV-Z�y!���vl^�M�Iޟ:��5���F��X���'�~H{����$���gᛚ\�$��e�$���&��"Jp��@,��~��tWRU仴�:cC�,h�i���U>4�s�GVi�U�Diꞿ^tޞYgYW��{i��A�uS�O2X��y���i���F܀����|/����#��8皴��9��^���
D�A�TӞ�nÚ�;�Ê<ɱ@q>ֺ�mgy�<sx�xmb]E⍸��a=V��h�E����Z
��P��x�� �|�f���c�uz9[��E�j�v����zە��mZ��d�Vg�7�^�3��GR/c8.�^f8�».Gi
@'G�ĕb4۩�h�a;-���s�R�������O�Gf����Y^�P/�Ŕ��H/"b/?t!W�1�OM��wr_���~�b� |����y�r�o��WUmx�̢��3���j:�7F���^��c�� qT�nIQGEaGc�0�ӱ��
�w�P�̿pٓ��TJ��ô�n��껙q�/g\|!k�,�qӺ���p_c�d����C�<꿟b㤚e�����s�6�Xfm��AU�H��v.��4oUǪ8�eDbr�ם�m�eشÕ�͸�jw���_R��ɛ����qw��j��u"�Hk���>�����!�gn?N���Y��j��wCO^�!�jאJ
+d���lh]g,�Kg�@�̸T�z�vD�=��L�c�Pׂ���݀���#{�n�z��wf�&��_7��7'�7���؊"���h�*F�6���#��)fR�h�Q0�R,��j�T�i����0���2R ���w�j��(َ��[}|�e�G^{%�c�5	�6�$CNƝ����z�qqoU�{%�k���Ԟ�+��*���g,׺!�C4�p����5�̌���jic�DF��R�݈��Nh���ZVv��mƢ	i;�ܬ�`ݺ��=ũ����.J�z���m�3bK��7f���Gn)�>WC�>L�gKaa���?bѡ;T�l�lV6��� n%�*������z��Cz,O* �jۇs'!�Y���ga��L������_���L�9��	�:�­�v�\I��Y*F"��h���B�΅�����"ʞy�Y�}t-��IGf���J�s�Ր9��ۡ�'veowU�$�w�I��r�g&On$�&�,k%R �pXk�p�=8x��+�I[�?,s��
�@�g��ex6�<E��o���3L��ػ&�����vu��m,��7Hk�"
׋5w�MZ_<1p3�����dGTGv�[�(��q����*�s>�g�渳P#��Wz�-��pO�����������)�j5.�����j2��HsS��XWm�z롇LNm.���Y���������|n��1�M,ҳ+��I��.�8�L�/1*��ߘ[?�����ޡ�)m�+id�nY���
����:�c���>7<�wE�s�ɽ�y�=�Ϥ�7����u�3;�OT�-\�\ѝ]uWƍ��(A�o����r�%���k���?RGr
P�#e� C�:D�tyd�l��j��%�W�H��K�=h����E���."��篚s��l��W��x��*��Lۓ�Zg��R"�	�T�&��5K�}���U��j~�9��[���P`��`��ucyʵ{Ԟ^�'k�xֹ���&��,���iMU��r��l.7���ç��F	��ٷ��D�:�Zr�_'��X�9��' ����"'�1;�ٮL÷�;�=�)6���?W�||G��n�+.�o��\׵"V�+�<��5��k.&#R��w�j��=��2}:c1����.�zU���ʉ'`*g�zݴ��*����k�y���x��^��E%`ڼ�/2��� B������|��VV�\��{�t�{z������3�'���zH��ox6�`�>��n��n���;I�qސb���)�"��{e�7q�}pꝷXL��t��`���ջf�Nip�l�܁Ru�J������^��vV/�N*���\�a�n�ѕtS敛�k�=��
ʦbe�p�� �S�������'޼��*	/��O(� Ď(d�KN*e(�;zW����**|fu���B�>p��߻EI������Pᅸ�==�d��N���ښٷJ�1�,/�z�B�����U��P~�S�cݴa;V��m��Ҫ�)ZeU1ܟ�M��!�z��\�K�3�&��Q�;mUox�����>�����?�r!����A-g��}���sϗ�B\*xL�ǡ1Y%�bצ�a�u��R�����M��ٲ,#Mq��F�u�o3���(�����M��;?����^�M���������γ3:���`g3�n��A�Q��~����y��$�1 ��Q'D2���D�X)?�m��|�jإ�"&��/���C�-�R<4�e����'+��{�}K�%o��vd5�������(���\ %��Y�%�.�i�;S����]݇���b������La�sȸD0N�ɯ5����c����Ξΰڒ��F�l��F�>M�k��}ϐ��r�l��烗�b����ʁ��)wWs�row��{��a����]��F���O�TF���a�K�A�9e�c�����t�;i�Ύ�Cq��{O^{h��h^=��x�}1������s�!�C.`<�1`�_.n��r�+��e�g�Y���*��ţM�]�I�9�}�5��a�̷L��D@���&�W�"��Q���gd@w��T
�n�l�h���r�9��.�kM��,��[O+u/�7��a�X1 +5�ާ����#��P�;�la��+��o���R�킥twX��ϊ�cT��������.�����j=�������q�ߌ��'R(����ͧ�E��c8r�����70�_&��}�u[(V���M W���<Hi�ّS����Ed��UU���ܭ!H%��
�f锍�'tϨXۛU�p!皋.�c��wLM+���Zk%�B@�(�=�n��8�-أْ�c�m��%�{�m����C"�6��&ga*��_+��+yen==��h~����8��*ަ~�BeK��j|����Se!�;&���5��{���:n��Y �w���Q��dj��ʶo[�C�����I��S��?m�����{���+6qT�򫉫cO�{ο,d�D<US�'��Zo+]^�X
;^>��h�NJ�%oz�ͯA����[�5꧗F��U��~���Ǜ,�=��������f� �f���H<m(��D�s'��/3����^�aֽ���.���=�ҵ%݉;��D�����qkU��[/]�Y�z�S*��/��r�����gW��8Ȁ+� 	�~�j��f����|����y�s��{P�t�+tvH�u�XJ��;�Eu����p	�k�1Mk������;�J��5v���[��^���f>aM��XvQ�ĔWM�tf��,�EoX�h�bt";OjPg^t�B��oig\=V�����;חM87K����7U���[�I��E5�xdRp^G+���`�yL��[��+��]cc�p��z暊W �U�Y����S�����u�9�d���[���:d7ܹ��4�J�HP��Ѫˏͦj떝��_.QU��=V9��d�4���n�.��fM�M��2)-&f7yլ#	�,b{��pEJ̢hbY`��h�E��\�\��mv"+*oe�#�v���{@��6^��gNZ�h50^�t���osY�u�0������	�,�j�Pu2�?fЫ�zN�'m��+Y��M�h,C�����l\�M�`�K�z����n;����h&b����m67I1�7Qy�k��i�J��voQ8���z��o$ƸV���WD�p�I�nZ<"E�b���{&LT�3$yA�Ys��K�m^F����p�۩z76�qv��}�O��zua�|�wk�mخ��ǔ{��y7S�=8�j\�U(>�����݂b[�! �q>eւ� ��7�{H���5���B�]>�n'����[�fe�R{��r�[Te�� X�n$녉Y�ZM�p�Hg��Lѳ��<A�)�V��I������_Y +gZrKH����Gf���5���F�O{�eq���	�hrXz��3��L�}�Y#��tf��#6��E4�
���9
J�+�9�GyN`���w-��#�V0TZ&�򴺕o�1U���N�M��(���9���Jc�u�����]el��i'���jŋ<��d:�*��:�h�K��t�lD͌Mu�q�1dA��}β\���miҳ^K���c���nq(�E�k���IrвH����`S�׋;��Sy��P
�4�
����:8��aV�1�`Ff���B-N�o��S%\�w)�oFH�,wlQӼ"n�e�<3'�:�}>R�x��̫��}��һ�ƹ��a�U�����F�����S^p\D�3(�v��S��}N�U��,c�0mjrYdSU��Ԛ�$G��+tc��6����fE���\�˓it2.�<&�(�9+��\��,v��:���K�%��Y<��ML��w}s��&Ϧ���]�u�Ⓛ(^6��ݺ�nm-5����#��)+bP8w�"d��l(>C�S���k!�D���f;ҷC]:��jk�EG�S5Ek*��������[G{�CJ�U�_7����(�LJ�U�$��X4�Q-fd�������IBN�f�!]�;��U�Թ�[��gI�t](ksr��s����Hd�s�@�`�WR�)^Ha.@d�ێ:x������ݸJ/y�ԥPP�	A�n9�L�E��6���o����}W�e3X!�K�j���`���h)�8��������&EE	CT$f'���C�I�n=�z}|x����}�*(
�()C��]h˩6������뷴5>FH7��Z�<q�ǎ�^=�/��P��G�J�����&���?:}}~?�h�C��-�CKJ^�QA�1��2co�>>�;x�i���FC�p����R��<��PSI�y�d��R:��{�
)�ސ�䡓�{�=�G\�����Y|rs�뽔�M�Umq8C0J�W\�՛�}�36f�(&�V�(�WJ�b
e{���������)?D<>�~�d :��5�Iv@<��/	s�M}�{b!�#onº��u�Z�wUvMm_~��R
z'����9�Pb��[Q��ə�ۘ���O7[�\,����-{�yN��kL�[�Ȕ)R~��uGk��L�ktQ�����Ye^Pm��ќ��z'��z���x��E���m�L�ha���<�A���W�6.;��9!��"B2�+�xĉF��5I��n�u���T�&��,g8�g�/��E,�j�h�4w;aSi��vs,�e�5z2��}���ҵ �0�7��~s��8t�C�&��F������x��2�pܩ�&���52{۾�Sb�ooj>�*�5�t��,����VeV,w�r��q�s�9�o�~�'���I���;�mo�@�IRR��rm���+2Z�տ�/��eR���]q���:l�1�\V�x�P�U�������w58$�����hT}��R��,���s-Q&���"�j5��Ə%�᧔�bj�q�u��i�:d��J�\ޞb�y�]`��Ųm���vp���CŽ,=�z�މ�-9�/�z��"���#��ԕ-I7�4R���֬k�����\o�������\����]��Iu1�
�\���6a{�N�Szn�w���F��o�����ȷ�~��U.�L�Q W^��eaS�X6����ϓ<[�eq��Wk|�i�fd�!��g�q��%?8�\�'��_L�gۮ5Ⱥ�%ܱ:V�s����m��7}7�¢(pr���;mf�ܨ�Nñ���Y]���yE��_�
c�x�duG�i}Pe�k�yܟ����'�Yr��=Aߓ����s^��n���Г�ϧ��0q͊�(����v)�!Y�9kWw�s�O\sE]��/4�t�`�oO��:��Cי�3��b+�fG��r2�{#e���Λ��-�����Hn�Z�0_;��ʬ�)����`]�(��1�N�p�[f��◄���>؆�p�C1 �M�Ǻ��M�g�M)ݽO9G5G�N�y5�ܡoZ�:�KpÛ^���+ña|��:��Y/�S&��̦��8=PSD;�[��m�:oI���G*l+&���Z�^�Rg�� �7����Y�?��"�]ܓ��y������}Q�,�"m"p�O�������������?[4x�e>1@x��Q��_'.�D6F)���&�ɝ�}�_��AD�(d�T�|����k2�$���##v���ф���U]zo��x�\38�
�����Ue5\��w�E�졑Nuk��l��̀������7CQS|�ݑ�X��)$✂�7>"���.nF;	*O!�n=������߰��f���pë�:%,����s�6+.66��U�9�cr��ûB�aW.Bپ�����݊�vZ��e����͋y[[�V��՝����W�R�#Iq�s4�V��g�^���{Ef�͓�m�j�}�a�@���z��(���!�*�#}�S ${rq2�E7}�޹JR��Ε�X�ѯ�UC�J��.;ws�����I��Xf@����Rs(���!�*�3;a�f�U�R)�p����͋"�ӻ�S7�J��J��m��su�>���
���wV��P�X��:�\��p�}k���}3��j�y�鉂b��ƍ&J@�XQ��\�X�d�+CHR]�Z�8�	�F��ѣ�e�ȯ�}�X�f��Dq�\�ֳ���8�/q7���P�c0���9�AH������fu���83�K���C�v��~�>ה�Xf�i�]|Y�dO�WY~9��d_��:�D%�1!��X�Ÿd^!P`۞�[_���χ~X2�ݲ��Wu���(٤j˭�d���Oup���_E��י>�[�
3<[y���B^��9�骀M�;��sP������V�t��R#���O���������~]��+�P��e1�yE��D�Vc+	H�͡�ۗB�Wܾϸm���+-�B�H@�
g��G����R#��ĥw���C:��w�*������q�Փ�1K�:��xg�L�zx�В���J1�g�a��6�M;�'x\#X��Ԗ��SSF�`��t��=�6���HP�C�QC�i�|�}Y�N�Ը�����ܮ�Cշx�n�Bv�ˡG^��:3�ݘHj��i�(H��;Fas,�C�Z��-����z�h��9�H��O�o^�++��=�{Pf�&���}.�;ؗ���Dv���P��JK/7
�.:@���ܚzk%���^�#8��q��I���x�'��}��2��G�5}q���+?�{u����X���G6���&T�xf�˪�(Mޓ=��~���-���<m���b>f��)SL�3�����YZ���܃Ը�U���J��"yY9!�.�lQ���_5�!�FP�l���ܮ�OlFdj�ӡ�F=7���
�N3e�DKS��	���i�N���;o42e��� L�ۭ�l;����\��wm��y���t;���0��>�ņ"z�nfb_wZWe-�jH�0�{2��S�nA'=Rs�fC��Kaa�ј��x�;~��P��*��?��"�����ͺʉi�����H,_Ew5��o[�C)��ۯ���b�]��Y2����&*6E����t>ŦAm����-Dt�*blݯ�g�O/X:WH��گ�yVu�䙄��RR�\�#�� �f ����{"b�]N-�&.�,���7'�J�=stnsVRLB�Ï�[g�,����q�*��p@A"��jp�g_]b7>��M���l�� �Y4CȘ���TB8�wX���j��bXy�y���{�=�m�$�=!���:]���#���%��T׉ɉ������Z�v���v��c��MɭVв��e����r�{��<#Aٛ*o�7]8��ٙ���4/�4]^�6�������y�]Ӆ����]$�5>�.�'ܹ\��gr8�B[IH	PY9$ժ�Y�=�5�Sex�?6�o7qf�ʉ�ɽ+ �������o%8wk	��ǘiܳ����e����H*�]z8Ǜ����hԳ��w��f�t>U��-n㹉��;�(,{+�̲ێl0iy��n��&�˧u��>q�1S�{���_UQ���k��`�R�2"�1�D^�H�iC���_ou��:�GdG��6ҵ�g��ړv[E��l�+��ۡ�cq	[r��u�m-�/U	�O�6�N�,���uGI��f��h��Ͻ���I:��)ٓk}�<���gީ�$4�|�U�Q�xU�r<ĳhl����vV�/N!N�;����]6�A��ވ��<���}^��r�5�d�i6��f��Ss�҆g$������X5,4k[o4��4;�l΋����R~��<H�)��$Q5���aB6.�g���a�?(R�KH1�x�~$���4�^�Ob���μ����׹96S��)fp���7Լ������me~SK�{J�1��P���Ű������a���Ǣ�Az��Y��3�~���9j��;�FdZ|�S�O=�h�]��܌���ƻ<�Ld��g�k�r��"o�d]�5<=�CN��v������ġ���V��(�gy�h�g�vO3��:��2%D�^Ku��ZUT��n@�!D�����S)g���m�H�e/�'Ov�v�N�7l�B���}�d�S޼�U�Y@%s����f��d��d��3���t���r
n3Oo���`2aگ{�稌<z�+eu*3����]Fd��Y���3�����M�y�6X��ߠ����K����fr�N��έ��^�ni'y���n� nԆ��$�$-�|? ]~��� ����#��t\`C��dS�o�=���C&�j۶�N[�������ԆCQf�����9`�Qh u���c0�ŷ\�T����N0N��"������SWQ�I�|=�v�w��m323E�5������L_�΀9M�^��(�[��gb��/F!m��<%����lؚk����֝&��BF
��	�w��q�8���+���臛��]۰��J��`��x}��>��
*k���$�w//?�~7��N���V��?<f�t>�Ճݞ=9= D$jy�a�Z�E���QݾM�q���b��m�X����R��M�Cf�X�0y������<f�z�y�+"� ����Iǳ�4����K�G�*鮎I�q56�*`7e�V�m�d�G1�!�6L��{?}E������n���d\0m�2���@ݹ:y��<�d��k�g���Ra�_OҦ��|��O��m-�Tǧvdmݑ��Ժ:��jx����M[�gc�� �,�鋎�-w��4��M؃�	ffe�򔈚��-�K�� IQ�����l��l��ѝ[ekXG������Cӵ�1�����y�V7��v<q��A���c���b8e]�7�
����s�ە�M��3)���ӥ�z7��6����E2�]�t�.��ľ�ֿ}��@`<�<�rN�*�u��M4 a�$:�djC���zzc�5
�����jٸ����#���;JN[?t���n]!�|��e��35<�s�Sk�����]��.7`a�ՋshYN//7w�dd5�m\�yRͩ�c�SYɬ�[�״ZG#v;Y+���Қ��+x�c���|3&ᵭ�ou<�Xyǯ��uޯ6�M(�k�*6��x%�u�7��ͅ�VvG.�Q�g��C�F���}�F��G0\����n��,�h4�c\�t+��i�1%)���my��ľ��!oh��hH�/<�t��Ǻ��=E��w�j�W���k�uC��ܣ��n{j�&��^u�g���>�n&3����6���Ja�Q�lWB;�4uA���н��^Vi;Ĵ��ݾ���Ǝ�_:|HTW�ԐI��T���Xv��4�w�WY�{]�(�_ZR�����P|�g�<��fM�fdFQOS&ɵ���e��S�`��~�76�3U�x�ٖ�`m�'R^�::6�NV��Tս�R*�ӝ����+jvz��y�{�0�7��Cw��)�?@��w�`6#U�l�qL2�����.<j(��q��_�'��^��<��ʏ�֍f8k��6oOv�RƷ�6����M��ֽhg`��لt'���8s�ef�l����� ���f{5";dX�]���G��Y�r���>CVp�S�k^s����4�8����k�M��Qu��FΦ�i�;���ag��禧~J��ösXo�m���������x~���t�Z]E,��YL��g���o*�@/�h@�����}�gyN��{�^�tV>[��JV�-�mM66��k�m�[.��<&h�9.v��a�7�-\��ތ>�\��Z!�CӲ����֥Y��D���W.|�&���^$�0dp�D���ci�������=�Z��W2�
��Ej�}���\�~ x _�
�-��}93"h�!�}�^�z�sR�MLS�V���T���=����`�)�w\������7r�G�M��⬊7P��-R�,��xk��)��]2r��_l��KDZ�k�w-�[��(
Z~@Keh"Af�]�J��w]��o�P�[�E��m��w�V0i��e(r���������Vk�٨z����J~�i�=�(���Z��qۘԽM�
�r�}�c��gX�*7ӄU��_q��p�S0o����R�����q��@�z��
j+땗�z-��8!Xu�z�E��u1�z�v���'qZU�޸noP�ܢ�΀�|�B��d�uq޹������2�k��M�܆Ժ �̍��6��$�6�oϟ�f�,f*�d��F�إ!�R���@Izu� V���w��ʃgS˖CT�M:j����-����D`/�gJ��Ձe,4�.H�ЛĹwv��( ��,��7+�X��}�����N�����3L���̋[��fij�2寕��+8�o��f����\�-�}lP�4M1�<v�n傮؍����5/[�8w�v�u�unYa���[OYi��Lԫ2;S���psUfj�d��+]��Zե�;�O���ʃ�kI�W�B��x��.��s0���3;v�|�J�R�('�$P� iӨ���bÕ�� z*0��ό��pu���8�\EBB��#��B�DӳQ�ah��ƻ�j����oɋ9�t��j��m��TT�!��2�)2��]y��k����іJ'rn��-�hu��Sl�٫+����.�53_}�o:'���U��n1r(!l���WcJ�h�G��5�F+���\{Ħ��9�\!�����@p*+�����7�/E_HS��eVca<֫!Χ��#�X/u�h��Ǒc�j����$X8.-r�I	��ۺ]�uu����G�%��x�9��o_��F�[����pw�-�|���/Z��u��\���т��Eرr(Vp�{R�\�`u�`��݁;w)=���1�濋/o�������XQv�1�sk-_
k.X��h�_[Ǚ+W_6m��6�{��nC�t:�A�'9j� ���CcRd��)r��s6��3��otF���i�"Xn��z�҉p�X�cڔE���6i�N��k�P�Bc����޴�್-��sz�ޗze��y������z�u��e�$����GWc�v �/��.�����CGF��1C�%&]�[��Z ���Ҧd�t�Ӎ��Z����H2̄�_�r���㛑�v�N�LCyWF�%N��9k���P�Xx��h�(�pz֝���=5�����8��W00_l8��D)r)ܪ%�A��dxvH=���dPR4�߷�OO�_��%���$j�I�S�u�:�hh
SR��ӧn�]��N�ȡo3!� ݒj�&
(>NAAE��N��>�x���HR�y�!�%��4�I�#��ӧ���������(����܍�{9EP��QՅE|�;x�Ǐ�>QI1PNA��VATѐoXRTCu�����U	c�=�}v���(�j/$�X�ʆ��#�5,]]y�ST��\���*���N�_^;x�T����+�2bik$��Z�!*��Y���b30(��������~;~=����DECA��VA�'&�Qfq�j��:&����ՃT6Vd5��"���,��Z�"�J
58T�Nb�w�fٛ�k��,F$�72$� @�`��lP�h6��%��D'0;�z���ƣW����� >Rv��0ࢇB��L]%n�^\��aں���}%�;Yq�]�����$��m�^2�na�L�Q	�Pl�Jj4IE!�G"h"j&��K���)�m��E$�D��B4�(�"8�"'H#�7j"�S�x> ��%�l~f4�w`�A6�*	%@BFx���R	%���e7�����Ia���`K�~t�j闌���jhX:Z��$�O@�R/jVcvJ��<�3�?h�cbz��H���;�cb�j���e�m��NȭE�%ܱ>z[=ױ3{#t�7,����*�s;ng�/�dC�4�;}3�J�ո�z���D���Y�:���s�$:��|�"��0����lF�q���6tԵ
�����u��~Kz�y��,	> F����6�VƪW�D�������A���=��^�Q��k�Lʵ�*��q-��sq�5[-��o7k���yf\�_N�>� �2ƙs�-����BOQb���D>�Jʞ�������e�fa�6�q��me_����'�t
�h&�Ic����Ǟh
��4�v�(B/4+��~z
����o�j��~��g��2=�TAZ ,4:'s?(fV��O�]�L�����E1Z:�/�ߑ�.ܮ�e'�'֊2c�VX�^ێ�,by�{�b�6}�!�Ձ�_\  ֹ1v�����{���	m�2�}�rb�T�_]��3��Uխ����ςz�WWv5��v=t�^���=<י�AĲq������}3�R�ҁr�%�/rm>�%�og��S�Y�� �w���ʆ{�kʔ]��.M߸�_Ny����}�Oa8xn����>�����̷O�^���K}>�K;��h���U�唏TWhk�'��9Y,m�-�Y� �R��4��B��	�T�A�y�Y��׶��e�W�r4�Sb��ueڶT7���N<K3�>E,l4���4���q�+�y���AO�ivXn)w(��h��V/���d{��o�FU�t/ףּ0gf+��lV�\a�%3]�~�_ZYi]c�h�#qT�:vߔ�j������C" �Q�!�`�`U��Xr����cM'�J.�%��o7��뭬.9��cր����!�>9E�%������(S�ؖ�ٳ]�C�������kѴjRƏ��q�Al
��뚫,3�n�.���wJR�^���{���סu�`!�ֺ�; ����k{g�f�"PLs�%�N�5�$s�mƨ�+,u��U��\���^=���^�֛��x$U~2���U��tȻ(��*.*�
�]Y�KɆ�Pt�ݥƔ,A�qj+f��4h����j�w��$٭Af���2;����p�Z,�}�^�"�X���wyMft7P{&���l�W�{ƌ�Q�ʡ'l[ԏ�+�����Z�q�F�6��o��bl���"EoXkx�#nW#��v�����Ѱ���S�e4������uX�ز�d�Hh��-��F	q��}����R��M�K�DR��~�>}NȚh0֧�r�j��~��ԧխ�r�B����!�c��#z��6�m��Kl^��3���T�e�:2�"Lf�s��y��Q&*��=fWVAUuB�:�^2�k� n���lR�U�6V[ڮ�ΙHa�;�#_�ٰ���;[B)r��m&vS�G��UZ�\��[>s���/�K@�v}����Ͳ@]*�n��.�x�u�ڸ���6K�?���]K[ū��v���V[9,h� 9 	Y;0@����錥\����t��'z �R��͛F^�]�N�#v�ǘz.=DPk�:B���P`�$ ��Z�^x^x�9k�{�UcYC~��W.X^�H����=FN�lUU��
e���ݹ}8Z�4��q�����5c7n�MZ���|�+�GCl��x�<d��� �7Vk�c�`��50�]���脀]ȫQ�摊�}����gO�� w+�{^�B�2M��n�uYq�l�M��l^�%{���01
���|��h��T�7l�J���g�U^��,����ǚ�i��>%�gs�pR��3ra�<��������b۩�Y˓up�O/G���𠽝K'n�f5Џu��{Su0��;8w�ѓp���ff|�����T��I��~�۫8}ަ�����!��k,�Yl���qeH�������8a%hg1�d����0&j7���}�#���Q�Q�.���j�Ig�s<ov:t�_K7�Q��D\#��_�a��%��׮A6�GKb���釮[Raq,�ƍT�vg�2v3��<��Ւ:��3|J�np
�l� 6�TK��m�Ӗpklm�#ӥ�Wz�ւ֘�`7�u����GE=���KN�z�̠��go�K��5����J��/��ݩ^9�7P����q�
)�u��XKNݚ�����Y���k���G���R�0��"ip�]l]=�):l���|A�4W���D��7aj�|{G݂�PhF�8�1�x���������3�'S�꾴�^�dQ���nu���V�\k[$l``�	u�i��p��\�6���D�3�^�Zf��P��N�lf�h!�^L�j�b{��/y����R8��zN�H�k�$�l�x��Yî�F�Ցƶ}]y=�p�^/~����*<�֪�c���9�'�3f�*�Ý�4�n�j�]�*�RZV�=��p�n���Mo]��w�,�"����\]k�|q��XP���A��Ek���gqi�F�<H��xw���)�%ܲ�=!8��k՚�]]��rm�gڑ�r/'������羉obG�A���x��+4�IX)��n��;/���}�y��thU�>�nI�B�����7��k��{.�"	���2w�3�i~ t�;A����p������{=nA���1h�ˡ8C��^���Q�F�`�x��e-N�,N����e��錚��]����<�).�k����}϶�~R�P��2�/c�����ȗ�����N��.��=���S�}V��B��0󺱜z�9�Xpt��)y��zCy�����Ƹ��/����	�Y����z6�P0|���@�EY{~eliƸ�l�����g�sP��0�>������G��䚞�]��ݯ��� ����iG��Ť���o�V�[��u^#Pۺ��3x���/űT��"nj[Ǎ�3�� ��d���,���C���7\�`�3I�dd�;�h����o�U�0-�u������z~�	��[S~�������~R�M���ɾ�x����5A�&W*f�܃��z�Q�[y�����m��`J�y�js�\����l�CM[~��� pk|p��?e�C���m�ߒ��xn��'�5�+F`\���r���M,�����է���Rڏ�M��+Ut�ħwwf{^��m��e��x��j�Gg��ϢDӆwgu���+�ףZ3eoXn)u����@��C���3�1�����E�ƕ�dǮ�%t�7�^�y}���D�;ێ��-�q���t��tC�n�B��h�nS�o�k-fh�m�TvI:�%7� w,��4M�`��-���.��-��9�y	O`�f��%�`Tx���NڡNI��j2�׀�����&����g��@Nzaq�q�))�w��.V�R]�z�1B½��s.�s�O�aiS��ygdV�������T��4�&J�o�Ս��l�����Y2q�/p����֍��	��vb&����+SU��ϗ�'�l��vwz6�'��u��-���l ٺ�2j���u4��;e�0����ú	X�׉�l{|��Mvi��`���3�v�T����æ�wZ�~��Tv���a�+�����Co�4 r�e��{t+���&��q�m��49�1B+��;X2����Y���_P�^���Zz���L�ة���(<�OCf��.�����-B�t���/����	��=}�Pj�J��l�G��901T��G��N�j�/=�A�i�~��'�Gb�;Oy����u�]cU��+�������c�{�9�s���-堗t��9�]�WԐ��b�F����,��f�F�@y�Tf���|G �y+��Y���G�9�us}x��*������6\Ѷ���Ҫ�&rbx���<�o+f��F������6�25������[bEbG�����M/Vb���j��]܆�Vm�aC!λ�M�n~v�H'�~�t|�R����ȥWʪd�f�m������l�R�;u�Se��d�Y+�l��)z�ݍ$&�t�g���W������sJ�]&�$uL��rC�[! �Q-�W���03��}���ne�mh�^��^H�є͹4��d�ս�wԎ��_.u�7rk ��h�=Y33T���"a�n�;}�ق|�:}��v��F��*"���Õ�M�ň���4q��]���F5
�gC烶�wN�dO8�
T�c��겠��3��H�PǨ;h���o����s���w2ƻ�1y���E����#��P8��if�y���ku�"l��91�q�ȶ�p�Ƌ�1lz�m�1���捾W6g:�ӌuRt
b�2?(�L�Obn�g��8�n��SY�����c/�H��~=%�r�����p�o�t�i�Pc1W
�*	,��6�2�d���g��e�1��2��3N�¾X9�C^uM=�1��RN�]�@��G���'?����
�H����"�P���Oÿf�;�(��4JBF�S�D�kѶ�D�|�Q$�����A򠟾F��~�%�B��V�wN�Z�؄���w9��̯��wI�B	��o92˝�Av���	l�f�u�\֍����O.����93o��Z��|���� �9�Ͻ?���:���jCz�����>�ՖaeMQ���!=qM�2���ܳ�
Z��ˊyw�o=+rvuL�ݔ�h�5�]T���W�+�c킷jf^L���u1I�=S��C�wf�G=5\y�[r����ǝ,ҥ.];�Tf-�o[]3�M^in|�/�����<�t3i����-�^��U�~:���t*0U�a��O�Jk۴N�o����&�pmL�����՞.U�.f�cV]�v��>y��\<ALF�NA!-������^�`s�:��cӢ���~�ql��kq[�g.�}���e�.���
���i �n:7�����O���K+���+�E�ʉ�v15�]�� �6���ߍ�-Jnfgtv�m�맥VC�*������]t���Gw�R�u��u��L���78�\)<���gŏ(Sӻ�Ƶ��ʼM���a깸[3F_F�N�j�?)����*:�CI��M�\9.帡�h�����ϼ�o7�5/�����'{՞��|�6t7�H6��[{U��4;m�Me��=+۸'��j��>��R}�w)�X��V="W0�w�Uݜz��[y#�rf��?qa��d��7L��S���9R���זּ��n&G.�e=�z6c��q���5�|�8b��4�Mn��q��+��������٪Gp����;�o���y�4�)��UF�A�n�v��]�5���G*ҏ]������8+���ɦPn_[E�ᝲ�o1�;�Ch���<��]���`�a�/d�rC$q�Gp�L����^h��dBV� ���5�j3/]W^�5	)�]�9��䊍��2�]5*�Z_���Sz;�I����m鞺�&g��==w�/�oW����?ԦkDx.1uO���<n��kY�Cwwv�w�b� �|�4���eٛN9G"�ʶ�Jyj�Umڼ���r�"X�8T+�P�n�S���5�낵�d���I�_w���!�4�B��9��q/�K׎�����ؑ�j(Ev��*�w O>ks
��:+2<�A��U�u��6��I̼ݻ:����Բ9;3v#�lÑ
w���M���3ö��g%{h��7#{
�v�<�>5��Ѳ�⩗O{]�:.L������M���,w\�.}yԐ���N�n^�}q���b:�dbgl�a���hoe\���l��3����R|[U�sy�^v�uCt%��d���`��4X	�^��a1����é�b�sI̓�X��f�t�KR\ʵ,��/jl#�na�	��k�C�D�c�qN�5��P�<�7�K]ڰE��2���sq���&N�Q�N�*�/�s̝\q���%�g�`���Ʋ�6����!���� 
����
W!)a��c��@���j8�ړ�f�!R��:��ˈ����7�mJ�J�*�Ŕ��ʵ3�B�6�E^�A��:2�(-ChX�`T2���^I�O���R�R��Ii�F1Z���s2:�-���;�$�(��J=RD%_<�پ�s,6N�sf[���=T�^L8n�T�2C�>J)�U2�ڦq�V ����l�3Tj^F����4(S�2�"m���ۨ�*�{6B!ve����k�2wn�x�30]g�=�\򞹐��wN7�����P��ܝLI����jmuh8�f��6�E���=�)��ũ��ʖ�ڭ�����ԬR���zU�L�-�5�Aw�o'͓��+��փ�@��s^���-rvɽSVN�Ԇ� �e���N�xv���sci�Ԛds+R�YA�:9c�-r�`YK���)m���#�B��a��lJ6+s���%�(%+�4p,�j�/�mMWv�E�t���I��Y�YDT�q*Ko�=�F�Ь�o]*S�]pQ�W���r-��ǚ��c�%s�c��[y�ԧJ�[�l��T�.�ͽV�`��O\������v�E��k�҅�n�f5��e�s;C�k |��f%϶�#`�wu�6�㎲�%-��'F)�h�B��:�7���M��0�ؔ���(���L�D�7�38>MVa�6^o=��%�z�0� Lm(�[���(2͍C�vus9�`�t7.�JWw:��'i��qc��n��C���xc<�P(�![݇R�J�f-���`�y0��g~�g�o[:�����3U	�-��a�n ��
*KcMW��*`�&h�ti�j\u!��J�: �>���wvz�-������̂f7����:�
(� ��l*�����/�eM���O�����AD�`�@Pjֱ���*����!:�D�T;v��۷o���&)(���*z��*,�h��(��
J���۷N��}}v��Y�L�Ơ����2H� ��=�!���x������ǰ�J
M�QY�-,PQ!UQ%L�9ӷ;v����|&��;�/3b)bJ���
��Pgx�TPQM�n�>>��v�x�QT�r0������UK�d�4�R13���<x����yTP�IT83�5E%$�KE�n:v�۷o�k�Z%*�fA�M!�u�
��f�����"��s� �
ih<̚��*H�b�(����(�-1��y�����|]m��ۑ��]�!�۔~=���9Ė̒��"u�j����oE䵱`bP�%��3]�Ͻ�<����jo��b��J��n���vJ�}v���� �ߜ��m�&ԩ���:7w�m�$�ǫ�:$����,�7+yS���ٖ��s����,�w��%��E�/�;�X<#\:{0���?���
ϗ�(zy ���}r5�	�q��<9[����/8��	ZGX�EiR����u�P��/��8����,���~d��k��u������%3]�5ԕ����<��ڦ�s����w0�c4�{���?��!�"�DJ5%�f��mWE�0z�mf�q�5�WbX,�	XՒ� ���|�p;[����kz��y�����Ϩg�n��c���Ƒ`�n�w���m��}�%��ln�=���h8���W�}�`6i�f=݇�A%�?W�Yl�M��x�2�ލ�q��Ϛo�!��ge��)�c��xj��_L�..�Y&u���ErK.w�ytT<���&zE�����W^Sa����EU�8�*��Oz{�������^�n�R��Cƻ-WP��g� l�;��Q�����G.��|��>�9������v�������<�;HWܐlQ]�=Ͽ���ӻ3��G�*C��8v�9^ Y��CA��jUt7���3�hܐp�l�M�C��d��ʸ����1=.�8MM����*|�8�r=u�6�E�]nк�w������<�^u~NO���[�����[ںSN`���i����UAm��6���� �k����T�ڻ�6��p�m�s3������ʵ�ůu���g����zsf�;��wGau�K��m�<��dt�]+%-D-�^е^�������3c��q���(�+�6o�:;6C���8��g����9¸�UM�a�#6�s���+@l�uF���[�;�ɸ��⸶u�%�_m=
Q�E�>�D[X��뉞>l��0��&��,Oh�fP��w!�y���ݽC���'�>����Q=��o6;W�G��pH��	�b��t�[��9���Ō������e|M�a���vD�9Y�؅�J�-*��+|�a̍q̀�̑��϶^�r@�T�]���%�T�hV񡋉��C���b��Nq�/xۻ�U8��W�RG���34�%�n+�R5Çm�w�S�o�l.���lQ��2�	m� re�����#z��!�#P���=M7�]���:]���b����N��� �z�1w�:�>	a91S�\��i���1�"#y�P}ӈ����=�Ƙ�9���i�@�aU�^g��a]N�v�� �Q��� (��Kb5�gI��d�����=�v��Y���CԍM�|�]�Ǫk��ȱ}��>l��-��#Zgg�*;n|g��H�֐�ko�vC"���=T{���<3�LD�������A���eW0�,�m��p��S"�� ���N6LU�n��[�X���i����l�uFO@�y�v�P؎�9rva���K⏧r��V��s�=���g�u�zqޠ\�2�I�Ͻ���NPI!@����~;pܪC����	��V���==��[5�3N�#fn*r�-'g�,�q����*��\��ffP*0ϵ��;���;M~~��w��K@�w{��(�7���du�����E�̨����Ucbp����I��P�ڧ�U���vk�U�� F��*Ф�`��O���c3l(�/�6=0���3��oSk���F��`lݭb��Μ�7$�\�i�ǐ�1n�}R\)�ndJV�+��&mH*�/9�y��1[yý�4�` �4��x���ϛK��ް�m~���w];�m?�BG��<��f�l���}���[x�Z���c{�\�>�pV�)_R��Xdo�6�h��;3��Wk6�ׇ���?@��yȹZA��ј���h���8ݷ#on�w�f��!��C�d��T�E�Y���%�m(>��×A��4ڮ��a4u6��ᖱ��tΤ����˟m��m�a������v�K�fa䨿�d{�N�{ٰ��)O���ʇÎ(��f�t�\�=�y뫤��[�\�1Z7�>�_�d2�y�ZM�b3a��z��v'~��ӛ�u����kBD�&(�������^�� 2n��ڋ�cb�	Z;�}��d�tոSB�߻E��y�9͆s���ć~B%g���{c���*9��$f	�����LaE���Y�<odQ����V`�	b}�M�^�oh���G�Y��?��y ��ʻ9��Ԯ_*U�"�,�������$*}��z9�;�;����ma~����׌<���B��X���w�T5^f�*ٖ�-~-���p`���1��]���l�Å����O|^*r�cʎM�7����|n���c5fQM���x���I�x��u4�U����=S~���(�e�Z�m��x;�nNc_t������%��DR�x�|���X��,��B7	���ȵ�1-��3"=�E�d���Vd�U��*����Q��k�3ot����̞��w�����焲�[�]ǟxz��客�!n� N(Ŕ���˼5�x��(#w-��,y�[�`�o2�w����C�ȋ�X��u�|s37`�z��`V�@�Q�ٟ-��j~�~���3m���9���M��hȺ{�y����vN�H2<��A/�`˯þ�Q\����G��>Rso����.D!���*fzr�@��%�Z��]�8�0�9�(MȪ�M�>l�{�)�k�yx��}B�����Ҽ�k�*cŮ�b�l����:�|��q�w��ҩ7v]�{2���ݖ�UȺ��S	Y�����-C��Γ_^�R��f㠮�ɰ�)+��+6n�ܴB(w�}�MfQ��S�)>
���1u����gt{��,7͞�4��t��®�������O�4�����sR̝wd�Q��5�>ѐ��0&%����=���:��H�ãMׯ8��i�8K@xS���g4er�e���C�7��
�L�����&�kWJ�Q��o9��#7LF�#q�a�K��!Y�D�*��۶�u�}Ɉ~�K��iS�-�z���K�7��Y���U��H/Z�x��ey�9�gqW{8�h��Fuc����M���@�k2� 0T���)@�;~���LF��'=JDe@�@��,��St��P[l���*�Lv��J�����vfj�O��ʩ	��9�=X�G�̣Ae�WUgoua�8r��'=���[	-m�`Y!�a���3a,�J\mmmD@�m��20����`��k0�s�p��D�1�l�Po<�(uL�����B�nej�+9X�1*ɩߤ7n;�^��&H��Ճ.�ܜ�ƻu��q��V�#S�۸RN�$�MV�F�d�Y,�B�u��{�`,�][P�3+�V²���{���a��셶v�0����+:��1'43��g��S�?u�O���Cc�F�y�vE�r�Ho_[o<�S5d5��p�W��Ğ���żJ���D��y���	�>��񭭾��foJee-on�#j��h�����c�޸Rplቹ�|�v�tY�����:��wl���[���2��z�f�3m�m�@��'{;�����jQ��8q�Pq��{�,$q �i���A3>�v��f��>��-��4]����_u"�x�\�����p�7b�57X�xvLj�^��gώ&���� @��қ�3�^-��csy�N6�wI4���e��3��ֻ$�E®�Z}k#�.�
��w=KgN��ww`��d��Ӫ|�l\�0t���v���F@d]������F6�8VƬ٢-%��w$�do
9RiG40m�bz]�!����_��S�v�q�c1�S��_5�B9�q��qw}���0u��-��3��Ne�K/f�Y�ج��-x���ԫ�ֈ	M* :@��U�;{�ew��x{�SS%v�ÎS?3�4�ବYc:��{N�/�����^�8�#sz�ԛ�2i5Ĭ�5J2���f���;��o-z�V^��R/)q�5B�v��S��o���hE���nΣ.�d���FTz��V��s���VeMJ�"w.6�p;.�@�b���k��y��1WНT��EWRm�]�[��$�7�������t4r�v�ڡ�r��Ty@u�u�����0�
��p�ƥ���y9���+Ք8�"��oV�u�_��-��z�fE���2���zF����*[ܕo]d��7Rݡ��#K�w�Pol�����#�.�[|�yo{\�P��X��(����f�jw`V�n|�vVsu���ƥo_#ގW*�N�咩{�2i螖��3S�z��-7^x�r��צ:+�%f��t�仩HR�͹
��̮������^O�4��c���DL�>t�UmT�&&��F�a��3i䣆ҠG��۽���Խ��*@�9���ub���]*���N��k��V�9�$�kh�C�G� �޻˵��R�����[ϻ&�j�Vn��� A��ޮY�[x�Q��Ck�,�>�xV���O��i���^1)��<�'�g�B{�5O�Xc*�54�e�7r�j:���<����]~�b��}|�f��W�^p9�[�`woÒ�����6��ff��/;A�=��״RW�?`���T��c�y;�\���vj��3��B9WH�4~��M�k��^�=���c�HI]�EZ���|�ٮ�w�S��{���{=+�S�"}�{�-qnR~=b9ُu5��;�@jU1|�B��W}E�ty�L�!\���[^u�hɹ�\rf�cd�2%�O 5@���=t'M���f��D�],8������������%sj]�S.����c�g����=��5�4�����>Eka9���myT��-l
vg�/�#�a���uQ~|�m��|�G1wo��-K��2rR��Y����O'�Ψ����"مTg5KI9�ԁFS�)��R�M�fűٕ�o_s�m�xsv|�QR̒*�!X3w�y�U$��(2��,��>ҽ5���g��4~����唜�CAcSt�l�{5���T7o2Y}ٖ��K��g\��6����ː����ث���zl��_^�;�:�|k��>hۿr�i��E\Pm���T{[��k����yJ�[
ق4�̩��,��Q���?)�0����ݭh������ӷ�M8�fMܔ+�V����f�����k�8��P�Z�s�P��zn�-�q��3#�3h�(rw����-�(����:,�������!��Sfjoe��0^]��.gq�ny�>�H���h6�ʛ�Yٰk)�.J���sC1+��7�9� �0������=���D��cpi���!�@pk�J���M���s����z�§�S���̈�t!<巹�UB�)p3�%��劅��U즑݇4nk*�Ά�/�e�B�"&�Vz�#ۂ���wTYf���Di�>�Z�4:�͆C���;��k����������3 ?4AW?�E�W������G�'��=X��i5'g��41�+ߘ�.� R$DpA�e0
 �"�! �* 	 �*������ �z�T0P�`�dA�eQ@� @�d@@�eT@�`D�A0D@�e@�Z t� ��� ��� ʠ�� Ȉ�� ��\�% @�eDP@�`@@�d �aP@@�h� �4�@0� ʤ3H�) ʌ*3H�) �&��bi�HQ @�D�&�%BV��HhB `��	�hЃ!H@�
����R� �,�$��2#!JȌ
��A���d��&>_��� 2 �� �N�>������?�������%�/����u�}���?���SO����ˣ�<�����`����]��?����~������~�����o��ҟ��o�?�E��~��QW��Կ�vBjLB������å?�@U�������������>���}N�O�� yؙ�ޓ�O�ƾ��
���""�C(�B���	J$�@	�	@��@3"ċȌ,��H1(�+@�"2H4 D220,H�@,H0���$B4�J0��J1�(�B	�2@�(�"�@3 "̃(̋,�0,H,� �@��@� Ă�H0@�H��� D$����"B�@��,���H��,ċ,�B3� @��2��!(�
�- �*�+ � �2"̃��0�,) ̋2�ċB4"@�+@�@��,�B��2-(̃B��@�@�)
4�@1"ċJ4���R#H,�"R(� ��-�R��B D�$JR��  � �����*�(�(��
ҩJ�@��J�$(�*�D��(B@�(� �1*P�P	0�B� 8~ě������E��
 @( �����������	I�������_�'��|���\N�?o��w��y�އ��'��	�={�>
�O�O���_����W��@U�[�e?Y/�O�^������Q}�I����D@U�����O��{I�i$���3��W��&��N�[�5?����@U����<����S��Q�S�O�O���j䟂� ���������؝%���%/�����-?�Kc�oI�G��ߡz������v *����5.~ݟ�t.��<�ɾ��Ca�??�$PE����M'zQ�|��?��Ɋ~�������e5�c�$@B[M�!�?���}����o��G�g�#�hE����J�Y�l�5�6f��V��%B!��؛T�I	P��b�EM2�"UJ�y �H̡�fbl�fȥ5i�V�֛2��lh�2�&f��m�V�Fck
�֣mPV̈�9æC�N���V��E21-�R)lklm��ٰ�ZT���Zو�YB�[m$����V�Z��46j��H&�.��z�% ��   ;N���I٭I�n����u��ku���n��	�֠�1w[:�$i7]:ũ�U�ٻ+��n�mj,u�m��YӮ]��{�"��Z۷vZ��Z�� �:B���B���z)s۝Z�v��vqMuv��� �c[v�I� �5j*J ��wl�thS�t�6M6�2�iU5� ��2�A�[j��c��
��t�Gwm���ذ`\�EB��S�P���ֻ`v+���P�Q����)�ۀn���N����u�QJ3n�TSt�qN�[��dЮn�[t:��lJj4\����-[T�6���)� ��t:��'H)��J�t]q�n���J�\�S�!�N�Ea��;8�4�1�k��t��mmB�m�[*�kx �ʪ)K˸(i5�����:��c�4 曧"Cwm�v�5NJ5��\���]��n�vP��΄��Ҵ��5�Ŷ�� ;r��	���T.(��7@U5��a��1Sw3��η5m�wjS���D0� WAuIѨ��KFԱ�[6� ��TP4\���]�N� �7U�E[h庆�WL�r����pڀm��Z��6�t�t�]:�q�[j�s���DX�m��� ǀ�&�8����[�@;*�X�`�w:�tk��tv�mu֔�as��4%�U�v��V�	��jR�mY1� u����]p �f�ەB�ݜ9]�fֺ��t+Fݶ�P����GB��,ф�f֚*���� � �   S�	�T�J0 &�	��C��)�4a04d�E?!)T�z��0   FLM0�O��%J�=F�F�0 ��M0� Bhh)���2M�=F��Q�OT��iT�Q�����b2i��L&4��|:'��2b+k�}v�<���&ъM��V2�ʓH1��B��U�MqL�ނ��^Jbq��K����A��ȁQP:DUJ(W��DPP,	���w_���������ݿ�ߙ�DJ��m*�����!X+  ���״��`����[V�[��HUP1 tx��:��P���ʜ�qrQ2���v�I:a���&B�I�w��=����ǝ��E ���JL�k��Q��D�̊4�N���B�H?(-��!�!!�c.'�#$܈��`�`%�ё�%#�'�&Ȋ0H��X���I�A�pA�,�$&ې�`��,�?Bj2X��Y�� ��"�$�\l��~$�������O���>��Y^����>����s��.�o_�wK������� ��T�w>h�(k+�@�S�Hݖ�Pn8�n���(��Ma,_��2��P��ȯ$�H�5�˯ĜH���',x�^�A�!2�V�$�!�u`K��R��b����q�O�md���
���׼��;�Ɍ'��@��iV����,`���^���N�G5ee����x��P���׿h�H�}ɮ�f-����	#Z��kkpK�U69���&�%x,�xP��k�qh�u��V�-	���s��p�����:aÕ"��i]F��B�.��\6���3f�����=v2)�䂻�mS�ܰ.�+e������������j[�m�YGZY��S �W�
UX-L@�x �4Cv�!0S�e0iz�PT��n�[8�6!iZ���1Xic�-�C�r�X�T���5�ä�{Q9{%��7*��!����^��m]C��^ ͇�5�lN�W�#2�u���L̎����C�2��f����K�͒��M�'59b�ͱ�d�M�owvy�	����M՘��֐˷d^+c������Z��є�L��M�/�ܬ�vqKڋ��f�Q+u���n�;��!Z�&Y;txq�B��I�H��JX�^��r滬�[t�����jc;a��Y��*P(O'i�"���q I�w/���z,����71j�&����?L����A�RQ�V�%��F�eA�3+Gf��I퀜��M�Aq�Pz�jzsn�B�j�5��ڬr�ݘ����{��Q{[|,u�r��]���Lx�y�he5c-A"w�6
b�YʟhH�ZX���5lk$�lwV�,��|v��V{��l(E�F��%���95�l�ø�[9y�-�"4rP���Y���o���ʻ^�WC��F�巊�=8"B�i6�Sfj�i9��k#&��D�ý�`%�yJ�L�w��7ˠ�x0�B�5I`�D<�+Z �]ř(��B���*8�U�;�����P���L�Gf�� ��5UԸ ��ZQ�,cX���24�$��iҧ��{�is*��>��@nv�)L���]��m�Rq#!�-�Bf�_4E[u�fbN*V�m+&e�(\� �,P�)�ӽ��p��W�;z�b�7R�P���CFnKHd�W�G�z�N��ys4M2�8β]`ؿ8��H�D6�.f=�!�uy����ųfP��Jf��mD���6�%9wxv�8bq�%K5t��j��Y�`���=̎.#�Y��xqB���O
fʩ��`��XaXÈ�Y��=�"�JW�Mn[���9�L�1� �N^4l�H�&3W�EGVHR��5��J�^�GE��彘�j�J�7�p��I
��A*V�n��̵R�um={J�]AY��rK����x���<3��[B����KW�0 lf�G��)fe�ka^���TouvQ�t��%)@mCa�	P��0_�����G3Kڻou�6ڒ�E�f����r�Xhf�2&[�]�t%�[D�ɉQZֵxZܫ�6��V1^�Z���h&�3VA�zb2�4\�K�i5W��B��2CḢZQZ�dA�Uy�F��L�6��n6�#"������ed��l�B��R�qdu��t�U� �&Pw�ݸ򵿛��$�X��st!���k>GZ7]`V'����u7D�����N�1���lI��u�Pl�9���*���yQ@hc�9��75s�*�0�x�iҲLFW���#��u�f湂ij�׽g�*U�������F�=h��c��d�Tx\���F�swr&�X�.zse��R�:��I��V	�f�4L٦G���`��Fହ(�L�YQ�{uv�u�D�)�w�wYIl@�2�]=l��1g@�Y�̹�n�G�	�^F�D��.K���Ǐ��*L��٪��`4\�wKc���ٓ.B�ѹ�с���y{�$hiV鋔Q�lP�wi�ֵHU�����6-Uz"W��˲,=�Mj_�DnnZIE��{��p��T�y����F���Ȼ�.�A��;�fGo2D�0��H��f�6�(�Ze�ۊ���g.�V2�n�����at�$�w	�����E�Y!��.�ŊK��(rke�q,�H����yX�`�o��v�:��J���9,�rk�&���bX�s0<gW`��]EXK�̶��/M˭��,��	zn�5lMi�Y�����h�T0U�6<Ѵ�A�\{NY¶#&������.�+@<���-�[y]��N y�o���:�sP�P�yt+��#���4���Wv�킺��|�7�����kV�hu��7��Y.��Wrk��E��U�u���,a�.�Ӛ���--\­Ө�2�8�S��p��`֖t�Ɩ���fn&�g�,O���-AY�ܭۂZ�f��%K�6����a�V���L�
�"�"q�gm��Q}�͖��f3N��`c�an��Yg$j����p*w���m◧b�Kf�	��̽�(J)�u�Tъ�䵦fH]�A� �MJ;��������K�*)~�i*u&+�L�rͲ%ݸ����h�E�3 �JA�^]+ئSXsc:-;˥J�R��3/0����bط%EYf�+Ɋ[AL��RX�HYB��VhP�����e�b<FC���-7�Ż���GN^�Lh�鹕�PJ!���F���f,� �杽�څ�Q�v�ڥBe�`Q�M��-�t�PѭR��'�6��)��ɲ^��Y�+�R^o;���"j���5�}��,�Eam���F��V��.
��H�:���tk�n=�wʼdP�YYP�I3�FnR�+xp�*���hҡ�"B��,ݡ��*2<?:�y�RӍ�9�o2��	wee��P:��|1J��_ehV�і7٪�(��^�Q���2ܫ6�WgTɷ7o�hD;��-�H�o0iō���3�����GS瘾�F���Џ&�xS�r����Si��盭�L�����S���֥�K{b����ٕ��*�%�6�.l�z���+�
�R���5�n�u�֓5���m+�6���7j�5��]���ۤő�b-I�˅7n�w �^��4B��)7Cv�jm;G\W��o&[�jO�ň�4�4�W0�7*Xu"�QU޽�h�w�gF�mVS���ܛ��S��,�q���e��^h-�ź�Q갉:���,+3J�z�$h��b
`���=
���P&jX�3j���J��OX���[�TytCa֬���0�˴G[�i%�r���B�;��Z.�Yf��=���3o 倡MW�fY���%=���� �GjԠ���9�B��-�h̄��X����U��%�觬J�1�7M�� RV��7/n"<��H�0PY*ֻ̱��5�	�渥��5u+f���hF�F;(A�k.�������'RRZ
_A���^�0U6��"0�ْ�6LF��� �OA�P��4ܛ���9�Ѥ^jf�lT�	�t�wBU�cu
�.I�6e�Gd0U�Y4�vE��^\Xn�r�`r��.�䧻�q�B)Cr`�yc�0�r^���n�oƝ��J����":pɶ��4����M�)Q� z��KRJ�f�^:� :NlPSзD[M�uTL��Z�qb���:CfY���X�j�r]n"���Ey2b`i�4ڳ�(h.�d(�ia �RG[:Ve ��W��#+!��kYv6�#T���P*��e-
:�Y�!�3pmJC24mlˣ��vd+���,�Mr�<cl�ܩ6�ҶPQ�F��3�J�W%[�6�֞�K-����,d���幕�l�-3�'�f�XEe�-��[�Wd�+%	�����{���W7[�j�J��8�n7M����v���)N16�וx-������m��"R��y[3]2[��i��o*lܫ�(�n���'pR����r�7lF(1z����*���#J���L�5B�UE�4�,�bb۔7/%�aȄ&����.�ݲ���i���b����b��7r�J6^���jGZ�;�S[dТ`�`$�4(�d�X�ʰ�t;���R���fR��Bf�¤�emI1��J�O3b/K"f���Ŭ��Kc����(<���׹ 3�o\-�Bmh�){��L���T���M9��D��!��ݥ����2Z�qfʅBK��mlK-b)U6���9�mf��5(./q<�k0f�^ �'ɰX
|�T�a�j$#X��L
ɹ�޻�,���XǇY9Y,s�������1o��\�H��&�Y4�Z��/]<
���K$j��ChN`*UM��+���X��s�l���̉ed��6�i�yz̤�G(P!h��m�t�e�,d��=�8��� ����z���H^��c�71���e���SN�nFW�P�3$���']�a����qV��684{�nMcw3 U�M�f�@� �yWx���t2��++K	�L9(�R��֪͈;�@��6L�o
z�oF��)�JL�KI3OeCRl{r(�cx���4��p	lÙ�@��n�ׯ.��5V��R�P;,a�h���p^\!�%�t�)��*���Ui�}i����4n�L�ʹpmS�^��YZR�B\�dbMccb�P�R�&9J���/���]����̼'p�^[�i��C�(l��l`*��t��Œ�kZ�HɍۚI�2�/k0H�y���k�(�-̆��R҄��~zY�<�� 񧦞�˒��h������)�]M6����],��a�Z]횱DS��v����n�e�e=|��Ѳb@fAzda;1켹c1���5�4̇JI��
�����:��0�ő�	�mG��x��:R���5Qަ�����0M͂�jo0%4�8&VJ:U�[hc-��Y��nnV����3Fe
��O(�������Or�[<�(�%ܚ����P�P�Wy�5�̰��:Y�*��{>��ww+��j�Jدu�K�����[�I2C6�޲��r�.D���;����N,�uI`Aދ	jZ1<Kr�hNh�v�lU��/l��Jom-��p�[ ҧ��Yf�.�1d��,!YNf�d!��AxhՖU4�hC�w̭�/\g\��6]JiK0SɭQ�������$�ȱX3bċŎ����r�YV�-ZF�S5M�������6f�wb�I*��b;��9X
LR�n�
�37%7���o��ۛL��+��ڻ�=i~��1FѢ���fV�D��;�T��l�Eik��{��(�bg8�xeV�� ���8m�5�&@�V�&�kJִ�H���"FK��E%$���!��M0AE@��AlĉAD�,� �T��$�2H�L�"a�	I@�)��!&�	6�H�J_�����4$�c+�M��`j&�g�&�H����P�[%Ŀ2�Q��b�2J,D6�-�q�M�-~�"�ԔQR7a'�G��E`��G�	N�|��Cа��ڝ���BA'v�C�K�.M�}���.��q7��ّ����N�� A30��x��dqP�r�+ �H�>S�,Ox�=yf�r�>,P��E�p���bA 3:�_.�q��w6�� 띅tԸّ�1i�{��nJvoEn�(mα>��;Vv�էT`����	� �8MdStw}C,����D�k ��<w�19�d�d�u��	��q�N�d��p��)� F�jE�୍�ʐ �Z������;��@�-X� Ƿ��O�Ah�J5LGn��J4,�b__Nϳ`��=�q���sz��GuU��H�k�fR]-�(��]	�0���E8�ɼy�k�N�����L�����&��1M��k\YMvK��@<D<t��f0�؜���E�m��U�z4�Z����ꍍy���[1�n�ʕ)��u��ѲW(rr�f��!�CB��*�ef�W�A�z��j�NYOmۄ�fIfddPrd����$��-���%q0����4�7C'�6+`pf����f���[+�s�V��z��\�
٢c̭@�yaܜ�N�/����M �D
�vc.�Fgi|���{|�e*��4a���ϒU����J�7bV�7+�ʥD�-�G�[�v�ר���m_V��R��&�!ةf��{{)�h��};���L�w� �3e^e�+3VV�h�͕�$��iٺ�c��6��;j[�&��gyl}��3K;2��x�jM�M����3�-�bR�^�C�tƺ�*�\2)oq�ݩx�혊@n0�>0�yώ�P<��e�R+�mW�`�K˸Э��;&,��p[���{y}��橷��`fr
�h�H.��<2)+�eޥ�<��Ɯ�Ѭ�J��="��R���Y��e=����5�����Y֤ؗ����#���b�ene��]R�\�l���:�Z�������\n����w�Lg�H�i�L\J=�h�	�U3��y8��Jy�΋����\صEq�]k�wj)*�[�8�`qf��c`��j=*k����`O:�L�	4q�g�㣚v=�"�rG.���i��xzz��嚥hQn^��@�4��Yb=��\	w��=: 6���j��F���1���ѭY3%��'�\��q�޾�@]�n���1�7�B�p��1s	3)]X)�k���X�Gnd�v�{�H$e�YȎK�����V����Pf(r�iUkUJvmdw%�����֩�_e�t��^c��������]�{("�L(	$���,zCݤ�a<u�k3;)L�r!2���c��u���J��G�,kmt=�j�X�]��q6�Jͣ[�&�^5XS.o\���<-�q��HK���vp�m����fn�Wʡ��}6��:��:3��f���7�i��3�9qT����ӏ��7R��Jsi�w2K���Ջ�Y�����}%��b�����W�h�Y�t:m><N�b]��	q�+���z�� كs��0���M��v�7�J�5����M�A�,Z�lڌ�Vؿ�k�u�,��qE��v�ȆQܢ�L�eV
u*����MCZ!dOo���+8ȭ���tN����i�ع���E/�deݤw�f,jk���B��"�3���˸�r8E�H�-��.����x����`YQu_^M�ב+'t���G8M9՟7�i��K��]%��<�vI��K"���Rl��0.��4�ჲ�Z=������k^�d���Z�C;
っO��̊5m]�5:�[ǙF�92�"�*M���W�_��6=꘩�E0ӻ��&,4����;v&;#��V��@DK6�	���L�{yi�]6equ�M1f�9hgꕎ�+RSa�2��lq�{Qj�l\��fuwt�a��;D���1r����~�]/]r�9��|x���7�5L�~��nL�l&j�w6�|����j�$B-2ej�3���~�m+.��J;.d.)p�j��㕜��弽�Q]�^[�m��2U�5�A�k���N�Ix	C�'gUeے������|m��,�t���a=V,e���D0��U��d�z"�)P��r�I]��X<�S
���ӥ*���^��,�p�x6�� Ca� ��C.H%�o��IɺY"wۯxr�'r7��K���٧�,qmkK�-����h3�E�L԰�5j��p`1K�ʻ���ܫ794��lk�O.���k�+��ު͛�]�G.%�ls�bl59R2)�/����Z�x�E��1��U����cB�A^���2�	�Ns׃�nQL�'I3q�w�Zj�7����z;��Ӕ:.WB�n⫦Eq�-� ���::(K��`ܮ
��  ���L�n�����V;ܟ ���h$���<v��q��&FjI��J�+���o%���WQJ(�䮜���:��+.���H��s.�߷/05��	��p�#|-_[��KOE���]��l\t��X1�]R5���6�K�:dY�V#�j��ҧ.��e�j�Fr��:L�vE���zӼ��ݩ"�ѣn,Lԕ����Y��rVݛ�E�˄����0��o��`�÷�b���͏�x��*Ȣ���!�S"$#)�]��é2>Ԉ�����y��+4�3������r���l#�^|ovξM]�[nQ�i>����r��=��L�97�i�X�T�$��8+=�f��ZD6��μ��q#�&�X��$��"�M�:��8��_�a�[���1-T'O�� �����vƄd���"�bvݱ�z*
uc�g�eA�D�&�$��P�o"��K��
��LNX�5#Ż�
c��Ѫ�"I	gE�N��e�[�p��G.;�9�&��g�I'pGLui����=/y#lܙ��y��n��y�[�!��x����ܾ 6F���Hr�1D���bz��P�'>�#Vl��Sw���s���p�6�@�kc�(�&Ԯ8j-��[�c����9�
��M���g�e�c�FAΛ[���� F�[IN锐5�4�wl[2,m������t�v�P���d�p���%�B�^��kb�ţv�]89/V���]ҷ������{Z�j��u�H4N���5w�#{��Ly��3��@��Y��qGc���K��n�L4l*Za����ۼ\�/��\��E4�-��C�<  H�۸1{�or�mM������ĥokws�X�D���T�+2�q�s.�Je9O2�r��A��^͡j]��s���gR ��c)S׮l�dܛ`AءZ`��y�'/���K��%�p��W%�Vm�/c��ڃ48vfڳdL��y+X��խ�E!�6̽�cc-26��@��f.]	�;�.���!e�@��ߗ-�r��S��[mw��!O
ᄣֲ�Sr�t$��h[���&���.���0@��(j��*j;��:]nv����j� �f���]�i��DS
�j�M	˖��fc-�wq���^u��T$�F:����ϭ��3�:���h�Ɂ΍d,����Km�]p�+Φ�o�D(+��>d�a��F*mmL���xj�M㎗ib@�Y8��-=Y�8��m,�Bu���@��� ,$�i�<��u'ow����t7S�ƌ{pA���l��5�U�4�܊���@np��;c9�Ιp��4�� LȻX��HQT��6U� :u�j��t�3y��4+��*�g<�ڌf�H;�O4s�5Nmd͔�GI�SWjі�2W9�9��u*ut�]�c�1f"�zH[P���`j��gM8�(�k���X4�I�6���_d�W����$Y+{��_\�{�j����2���#g$׏�T8�%�v��\��'���k��Y/*����ۍǹ����F��b���8'\+]TC��Gɫ�e�4N���a���9�B�oG�4F^�	��w�橜g�86�����B��,k�i�Tm��IS17�.��n=2]u$	X*:p1�2�Z���m��)dJ	}YP�=�O7��FK�w��ےTW���wb�6M�]e)ңή������wsi#L�㰢��q�t-���pPkV�k�ҩ�+��c����f2��EHGZ�z�[Q�|t-�\l�ŋ"�ʪ�Y����K�Α��@���۹m��h�v�Q��g���%(yV���6���H5��#+�4��j���}B�<(bǽ�Z��)��ܡ&Vz��i����� A#t���琛w�e��ݧ��la�ְE��N�7����oP�Qd�ET{l�N�S��tn�d��{����#Vb��u��fI�`�i�W�ed�1Nv\t��Ǘ�e�7�C#m���FmQ���P��@7J���O,]j��(�1mK/������8�e���`Kiҕ�W�����:{�@M{�|�g��O���G���5�39��ޗ6낖ED�Wh܋��۾�e*��k]#�f�AaҮ�\/VRRb�[pG�U��9%��d�ëaou��n��˛H^��R��K��ۜD�B�+�U�^:����X����ĭ����B�)\DWF�MȍJ{*�e:�We�ԫ:�9ү�+τ��;�V<��]E��Y�ց��(����T�)fpUz��nظ�p40(TY�n�|]���P޵&ȇG'g��s �fu�&��B�WOd���Q����!ډ�����h��9�}�X��<�B�fgZ����`�� fV��CU�bp5L��ec��r��Y<�k�Y���d�p�p�4�蕄v�z1Mj͊��k����[m)����Y�3���u�YR�	h���+� ��#ݫ&�6�:7|�3�K9���D���^@�d�Qƪ@��J���T��M��ŘkS+*f]�m�K���P��\��U#ۗw����5j�����]ҕvh�\&$�Tla[{����V��X��I�Ae�[+oZ��^K7��J���H��z�b�.�)ٲ��pTrrͤ�˲�{�t��7�Ʋ���_z&o�r��s~V2E܍�3L���d	f`k��{�������j8$�wsS!�B�y�2cW��f��
�ځ.�r����9-��$��$�I$�I$�I$�I#�S2v'�p�GP��L����Y���H41Nlf��%�u}��6�� ^���Y㚌tѕ�jfR��|*�x�9(�B{���W�z�Y2g+����X'�T:��X;|�2_�\W9/0D���3ϗ-5��=�a۶��'�(
��'Txi���X�8�VE��3kSZ��K	n5[q
�VQ���2�uj�.��wK
]��.6Vm�_=Wgv۫��R�"�&���B"EM�cm�P��p
:X�&�_�+. ���:�[�e���L;S[c��5J�T�݊V&��j��7YZ��{��t�Hd׺vc)�kWf�Ӭg�N'+�-1�EcS)ٮ��f�P^����,Bj�T@T�;�s3�-�T_��������w�8��hc�}��ܠ���;�w�A���6.��\�p�i&ž�	'`"�l\�?����ʑ�mw�]t�g���w���ܰF���|��f��z%s����	�����Y�fu[F�I����+%�ۦ;<���B0�Q�.�{�=[ ��15g��R2�k9�hF��Y��ͫs1�2AV+(/�	�d� ��� \������3hWf��3S���<��-q��rL8Mc�D1୭=*=W�@P/����:VJ�F����������u�vk�q
N��O�����1JK6��������7Bꗤ-kHeX��P����x+N�S��3��::��{�G��h��3*�͜�XxD���knu5��ڬq��̉��C��v+!٦V�c(ze����Xf�3xm�.�φml�pL�ŗ��_b�E��RY�\�y.ۑ����4�_ic�U�4�fl}��;3}� O;����J�qsڈ��b���6
�LM^WE��[�,}��<�N�a9���;����sMV��<�eȃ�	L��r�]D�zI�Z<[�p�p��J�d� �-c���������9��L��vD^#��iں祲[��T�d��lX�x�����/n���ݦ��©V�cSұ}��֍;b�<��y&����)�=ۃ��i�8Ҳ�q�"�k'u��O�oZk��쫶�HL��Պ�k�q�`�Z�S�O^4E��!�+�"��{%�$�7QG"�<:�M���/Eդ!���!�eک����y�;i����*����Rӱ�ef�ۙQ��^��pV��p���5�ܽ�-/1���6�.��/h���Y\�z*ַXu�� ��϶�[�@���WIb�ۖ��+O�J��I�;�����#	;EV�]��#��f����я�q���Z�y�v��j�����Zg�b�T���A�6�яOl�=O�����r�������������x�)V��D�%��.���.Ֆ
꽅���������L�a�޴W�2�2c�{�sP�A��볹R'L�%�Ҿ�1��$�n��ZF�%2�!���˼�ᶨ"i����펡��G%��Ѡ�u��VS-ڵϷD�c�ڔ���m1��-
��"��ad��K��.�@<H�9��F�!E�+�����\��Yr�q�k�ϻ�qh��� �;!��.]��י�2qͥ�fi��`뫔6��G�L\̔��]'+���QS��ea�*�e89��(t�1�n�kڷ|7�7�8%���m�H��O	�7oMe�M3��h��jK`���\v���@kq3���j�Y���,�+�hnRf>�bu���g���Ń�[s62�J/%f����+����(.� �f�����k�p���P�ln��*zZ)E���T	�p�Nܷ��=�	+y�[�l#C���yHv>n	�w6^j�-em.��Z<�W�.�5�z�&�U��:6��cJ}2�^��{ݕ��*��%̟7��i��T}�{nVܷktDI���g�1�T�J����J���i=���$&��'���kS�J��B��i[`h1�Ͷ3��+B��v�ó��r�� ׸t���$�IhI�owv"+�3w��괝n�S�-�!8�^u�x�u-N��T.�"n<u*�
Ů�F��٨�Y�E:cF�{�ogƁ&̰�ۚ�M�I���r��Yd��bgX��>oiT�2�M�n�rUk6�uJ�h�
Z����Eܺ��	�yjЍ����YW*��j�9�_s�G��U�R�Tğl3]����ɚ'l�� ����Myfm����v_-�Bכ��PV�w����f4%�Рt�����bV�~�f�-��w�5��Tz2�L�t�Y%�2aO ���QЛ2a��z�Y2��G�+�n�pd{��
9��LU���îݺ���4�.,�~F����ۤ����WN�5�cAS(��7{mtr�x/�ٵ����@��Y:�Kt9j�����������P�yz�ؔQ��z�/5��N��绊���4\6��o�]�L�뺝(m<w�A
N/�*�.�ԛm���$W�����EME�/6�AӖ�J��Vs>ʱ����P���*���*���MEz�+�1e��T��3�Yv��O.�Ui�sk3 .�E��U��� �g���{}�,��� f��J����+hlF^�t�.7���d;��dͬ8R�]H-u��#R���k�Nz6^a��@�Ne�(���m[�S��r�Ͳ��5ӹ�T�3��q�x���q'2g���Cr2N-Df��y.63*��ȸr�� ��I���'�����__Z�L���aeK���������u��w^�eDZ�UF�ɔ�,3s�]L;+4�ۑ�w.��yb]�|�C�WU���8ﻢ�L�v��(���q�
����5G����t���q��u�^=Λp�����oP�[��ui���^��:��1���̒-	S���WKD�lg*Y���Y����@�3Zj�d�/b۶/���մ;�K�z������:uUB�dַftý���e�e�|F��%�1�K}�_k�Q����S�T��J�#B�0���+�k�"��g:.U��:6f�
)��gs�OO�Z��7՗u|9�蜱��*��o� ��,,ᷖ�
_6��״��~�{YB�2�D��0X(:���|�Va���L��o�d�wg丹���Ф��UiQu��3vU7�Bz�?/w$::��h�=�V@U7kP6���k�v��kS��W�i�?��b�2%�~U@�!����4	5ͫ������?=���Y;��V l�}�h:����smWr�YQ ��v��\��q�:r�PNy�B�_l�������[5Be彷B�SPud��+���6Rr���gܧ!�)ګ3���;!�"
�iqN:8s'K@D\򲊓�
���ۯ�A9�QUV"c���$h����w&$k6��UUQ���h�~��E"I�5��j��fw:�]+�V'E˸t���óMK�6º^β�YL|Q�]��󢎷��&��?.�L�`��X	Sg�ߡ��^�A��X���%��,6����K�57���X�^r�y8���rTkSz�i �wSrTz���"�\j�)��^S�Aݼ�A6�����7��	�̕�{'�����}���F���̒���UY��k.��y�AX���[ cn���S)�\I�u��݄B�R�fhw�orb��'�1���}@����P�3xPͨU�=�]�{��_TDU��m�<�����8Rb�57]t��;�í$o2�Bc��®�����Æ\�Fut��K��E��n��-H�hK:vuL�u��&��qim-ݠ�:t[66�D5%5(Lj�Bom�:h��0謠+����x�%��U��N��}v�~2���Ԙ\�������f��M�`뙕_���G� C ��Bۥ{��'|�u����*�j�4��n����O�h��X��]N���H�ܚ�n�w��b^�E��Wh9��V�o^Ú7�����5�W�L�ڪ�40�
 �Mu�5]���;2g�ʤ�����)�,VD�==����᩠���'�`�K�rR��̭s�m)�d:~��)�M]o�UUt���ϩ��Ψg��t_��~̜���W�ٺ��k�Q%8��Ò;�YU�s0S4��#e��%���w؛Z�d̎`Y0�[��k����@�O2�Eo n��Jt�o�X��W`,�b\�^�i0sC�K2F�b�FI����+���#�"�c�dV�;4�|5']N��m�_9���'\)��~���8(�tl�B &F��0M��$��ˊ����cjdޮJ�m�����ۋ�o2g��8�_*؆���n�n�ge����M�FV�����r�K��q��o��ٸS�_8n�0G�v�},睪JwwU�����%�0`�5���K�yFm�{�Pfqۼ&@��+���i�m��Y�(Ɋ���ذy��F�`_r9���w�}ۨZ}�U)c�42+c�j�CJ�v1��! ��0\�/Ei��L��Z쓬��B��W�ݝ
�h*�U�i��:;���Ql�lky�z��}w��ӟ1�[oa��nt�0����!v;�W}%u�����C�y��u���a��\8�Kn��b�ڕi���U�*SH��C��*y�s��(�`G+�]�yo��ssQ7�
Ů	X��3�]3��z�l�� _U�\�
�Vv�Ɨ�*�x~�~���+C6�/6�B5�]�u*="q�L�*�{�����z\�����{�Wٙ�jL�G���p��8�v��Q�}��P@�T�ŵ�bq��u/Zb�9;�Y}�¸��ݽ���v�W$t�(2�s�w�V��0u
���V����s0��8��5�.�U��U���������O�P����6L��R��=�o�x�����
ޛ��̒�_Ff���Z� �=���W�U�j5���E��g1KWi3Z��oCT�t|��bw���;�-[���t�k���V�Ur�*�<K�f
<3�.�p�酰��K=���e0�C(V��a�?:�.��@�<����Q�vaС���i
��LU�3�*hM\�ڹp�f����vI4���]�C@}\���V/����#6[{hsZ�m�˖�9�V��i9�����u�4s���B��ꕏ��&(S}�s����em����7x]η�v�e�:,�\�JY�ws��2��)lݹ ��
�9�^��zWVf1F��S*�p�3.�݌�)�z�e�HOmf٘72X��Q� �DŬ9s,]bh��:�����o"�����D��YlI��ie�}��^�h���fv���^���s>�v`�/)'K_W}t R� ���Gsu�Y�g�䧛��ݹR�S� �]4�!|���_1V�u}�;%�f��x�r�����:���o-���d��72�eu\xGL���J��B�Hj͏��%_wZ�T�b�Ne,Yu;�r��nw�[E�.i��/�w\qʗ�V�5��B�+9aM�/�No$/��Zx�sh��i�w�N/�n�nn
n��X�ױd׉)H���١�8
�e�31�1�]*�\[N�U�+nu��uVqcr���WoJgd"�{V/`>�n7��vQ�F��i����LF�R��.��q8��]��,ԧM�lh�ȇ�T��u��+�X���'W�p��MMH�9�VՋ7���O��A�'IV�F��&���{�����Y{[�=�)��3�Fq��,�|�x����o�r�j�#�Dj�JE �����ud���������pH�&�`�D����A!
d����0?�6bL�(��$�Pl;2�i�	a��`j!!�	p��A������܎nu��ͻ�M q	YCC�$�V��nI��>��Bp�WH��N�O��=�}`��u��J�ج���5q��\�P�%���5]��+5)��+�J�%�Q	�έ���B�X��<m3���v��:�PQ$��!p���6R��ŜZB��9��m땱�e��r�࡛��uIn� u�	�X��5F9�3����/)*�˵h��i�XL]�#��ԍ;U����T�?�9Bx��S����8ּ�~�󐝗ύ��p��T�I���{�J����d�Ǖ�7G�U��|�bckUm%5�l5��EƛV�c"(Q\Rvv�u�ӹ$�4U�y���t�PV�4��&�p��=;u���,��6�7�|"xC�;��wkWe�5�^a��cV��S�1���r�:���uh�pa�lA��0V`F+}����r�P�j3����ۗ�<����-��kiV��H1�H�Z������������L���e$i�pe�d�c���?}r����]��te��v�ݑ�{޽�12k�s%ξ��v�d؟�wd�J9t�J�hHf���Qӛ����$�2hA�}w��\W���wK�7���:�st��{�^{�>|����޻!�/;��{��]�.o*��ڣk����n�����;�Ҟ�v�m����k�r��ޖ�^�{�����-%�W�uEr���^��k���|�{jJ�N��:i�z������ך�����;�/�{/c������w����ݨ\��v��+޻]$�j_]ni{���"��w��]�\r�͞�i*{ޮ��wwO��wg���v뻝�^�{��&�*����\��uwH���/N��|����E��{����w^�ӻw�{{��g;;�����Ļ�`�w�uѩx^S#ON�9�=�^��v�ܮ������H��;�]���`�4(�9���(׺� K���˒/�K{���w]���T\�����k����=|�$�(�"\��%լ�ѫ1��٧�Yz��֗E+�n[�o\oM	�O�<��d�����p����V��������{�,h�
܂b`#����[��CEG��Wߠ�wp}���~��d��K�d�u���]�%�f"G)�}֏�%�Kr��񗇵ڼ��Ę;}<����2&/��<(01S䕋�*�3 ��ݕNfu��b��A�X���CA�@�ڱ/!�˨X,bʽWWcķ,���ቡu���H���Q��~!A�L�l��Zt��^.��M�X=���m�υtƒ��!3�<N����+�g�+,�Zr>k,m���{|EN�3IG������R����y̝�<�r�*��D����o�=�4����y�ک�[g���+���O�]E�>��o2�+xk�JnV�u�f/|�yN�dA�����Ε͋��;��0"�|���|=m�Y*kw�떭�!]T�K)�w���L�X+L��~WuC_��c�bRi�׺��\�[��%����Լ=D[�������n���{�a;:��0g-&Vf_"�M�1���T���Ӣ7���������LN��b�ڋer.��|�����3����u( v��{���V�>�Y��\%��Y^�](��F�=������Wxߢ��'b��V .��tT*a�*�pl�f��δ?���P��� [z�fk���\�tf�`���Jcr�Ӝb��A�`�14���:�j�r�t'��	��NNp�o��ԥ�K�L�^���?���L|�l4�����������ڣ����'8�^�&�\{{uW�H�N� ��)'��T+����'jd��W�>�J0۱x}l�Yk��g�yN��
b^�W���/�s��vj?g��;@���\�[:�^����Ax���!E�'�H_�Oؔ�8��@�h�}yavF�OU͵3�iu��'�_�l?Li������DE���B�T���5��!v�v�ϐ\9�M1[kO�1]䥽$��(��K�����ÇT�]2d���Wa;�>qT�+x�ܨ1��3��ˮ�E�,۳N�j�yr�.�ys!�+�֌���	��>�dV�o]mj�M9q�¦sВ55)z��^C���cG
���(m�i�"��C�D�Y��wf�	�����B�l�;��_��ȉq�5�R���k.���w=y9Hx�Կ�z���\�_}w�r��[�!G�dp�� �����Tw���X�d�;�R��|�84b��[F������(�n'�/[�6��'ߣ�BW�����^܃K<f�#Nr�D��?{�wU�b��Z�K��y	\�ʆ�����͜n�yƎl����X㚆�'�x�׋�D	~guQ��3���Y�d���MN�n�c�p|��"u�������=ʊ;�(F�a/D #M��j�佚�&�'��D��8�E�i]u׮Dt��er�/�uz�iJd-VfIG�x_9�<]�wo���ꥦ2��#W�R� 1��zW8�3���{�
�*c���YqE�q�p=��ͱu>����"�
�s~ɕ�:)�$��ӂ�h'�!}�K�>J��$;ֵ�.O��z����4��W�3�c_fYFM�� ͥs��¶�F^�ˤ�/�,��t�� %'R�f�^���2B�3�ƿ� �VÌmq0÷.�ծ�F���x�el\����ڡ�q$`��(�W���<G����^��;v^n�����{; ��]d}]�@R�\6�2!�^��B�Q��ʥr�6���p��=����(����U]�'���P4a?xhC��r���GҽR�
�|�TdӴN��ʯ���J����Uo�x�@�_x��Y����_z�t�ݼy��h�yx�1.���+��6>��B"��"_��">�Uș��l���+�m�hz��|ɾ���6q%�!�&��xF�$ضgc�\S{��YCo�3����g?~�7~X|Gn6|n�zQ���!���,�m��eF����ǐ���0��c���� hD�;��x�	k��ջ�.��%�$��KW��Du�*{a3�k�w]�g�q��f�����8�Ӎ�d.)r?}e�/�ٔ�v�9�ef�:
�j9f�fۥ����T���.�*�P�e��[x��=	��F�wH��� p�'l�RP�b��T;h���.��1A]�-
�+��ݩm7jSt���T��A�]e���r��o@�!�9X$�Xn��~�Rg��	�lK�8��}\��1��������tz�`3��ʬRV<���]!�h-J�9�#;ٛ�z+&��V��;g��L
�>HW�Pϼ:i�w0�����?m+�L؋�g��Ӯ��R��O�8X��gG��������r�ו���]s7R����~�����;���F���q���]�2��X@�0GM��lwK¶���M��'``?����4|w�]��L�=��������Hl���׈�P���KW��,06c�{�ⱄc�$絙^�#1�6{�'� �����z���H'�
������5���}f�c��A�:>S�U�zz@�C��������%��g��wj[����2!<�r;Jr�=�I��V�k}�����y|��-&W�'��4����̱�jF�,o�1���Q����������0�w�e�֨��g(Q:�V3H�o9;�Ci��#�ct�Cr��i���J���r���Oj�54�����3;k(��'G/��&;�ӟ�
��Z�!���ׅ,�L��U�Z%n����wvi�D)��~K�b��<o����+ʌঠO��=r������w-Rxa}���(��g�`���{�J���y�?�X~�t�+��fM�z����92+�<���5<-oP���痴���4UV�Kާ���Lp�!
��N����_|t��_)��e��U���m�g��,����~U2@4��~�+�5�����!�\t���3Z��
��PӼ��z��7o��=�>�r�x�'�BH��l#ǲ�܂����xE~���0���\0S<B�<3{����B@obueG���ð��-��r2��0��w�^��y��+��H�>��]i>0[q�@˞�M�|�)��xs:�z�\^�`x>�A�	{�;̜���������a.!�D�B�������!X�=��Z�ڝ�L�RǇ�Y3�{sb�9����<���ةY=�.ɇ�d�r�Ը\�[���u��<�6��Y�+!鼜[���|n�N��azzq���5��T�5���fsG��L _�nnM��ѯB��<.���ʀDtG��@�/���*`��E�-y^]����q��z���k�}��U�T<�Mi��$/�1�#�rC���#�N�{o�U�W����n����1\/���5@Uҭ<��#�||O��*=����8ߺeԿU�I+�hi����}�i��,�h/���W� F���j�k�x�w��QA��©{Ȟd~Cǰ�Ev4p���?_e����b��\�Q�k����������5�����v�!��X��tU�j�Hm�Sz�����3^�#hVRNS*����ۭbx}�<`��4�˵���W�k���������e�(ڿi=��a����H��?4]�%����F���ҏ��.��.�?) ��h��x7	��q�����{��52���|�ѵs�Q���G4_���=z|b3��uсؿ@V�ny檶�x�|��{���:�:�a9���
N�|��m��7mj�o���Z`�6���U��a?et�F#36ez��B�5/�Z�mep�S!���O�G<����x!�4v1xv�^��kn��{���������X�K�dڂt�;���5o ���+��\��X<��TO!���� j?��!���u�$j�S��=��+�P2�1����b�ס��9�/�C�y��_�������q([���wt�Q�^�X�Ǘ;7�Yh�,�2/�ƍK�A����_rO�Pj>IJW��>ңg� EULT��t�R�8����\�$�Իo�����Ǿ� �k�/�2B~�7|�h�,�)�X"��v~�]�;�j�E}�:��1mk�U1�]	��#�����eh�x��h`a�e=��r�'<7QP�O�x��ҡ�Sz#SX��4�#��{�*iq�#�/��6�8��2�X*D��~u�T���.,��>����h�$�ٻ��?�>��"ۭ��>��}�|~�w��Ү7j����ǲ�|�?R2�B�P��pt�a������a>#9#�ˤp���c��}:�I&��]��F�����aՁ��cݝv[���q�b?=궻��I���4??t oh^~Pw�Y��4���T���wKO�=+�ePV��RYZ�g�.P����NJ��E��R�z�9zɾ�=y��/9�>C%f߄�"�Z̚}��o��M�>q�G؅��ڧ���yXWБ�1���ƓǟGQ���P�ʮ-U��x<\z/��{�vg�<�Ë���3���2����?^��>r��ۙ�9Cr�$����6��~~���LI�����2���R���{e�A�i����l4����x��XņKsU���D1v�{%�7�ű�	��o�}�0:�V����p�j�����u�X���@�F�j�a��JG��?7۱��_��Gp
�H�&W�U����O�>�8ѥ���Q_]+c�=�Ofyged����4�\T�vK�(����46��U�W/
?���>��^8m���$��BIW�sk�߼�xU_��Z4t��A�L4C��!�/yU�+=t���n����^X�B�$����׾�@4��C��;�@(H���|p*�|ׅ�����"�����{#I��j��c�_Ob�� ��Zh-��w��|ߺ��DedZ�3Hw��� wk*��ea��q�p,퉻'��sy�}�������U���T&Pu��H\8�'>U���j]�w�Ds꽼徭�+��H�lɵ�N����+B��E�_�f��#��
������{c��߅�;C?1�@�x/K��:�gH'ŏs��EM��I~����Ä3~�*��*�w]��CÈ5Y�/���Oo{����[Jϻ�w��B&�E��da����B��=%�C=O������s/��j��+:Q�H��/����dv~�Ha�Mz\�H�D��2���}aC�n���?G�^lY\��{�կ���I�W.f��ߦO4�ޞZ-U�o`�+��s6�G1���9P_o(64Ev�=�wQ箹�ؑvA�k����G�ނ�T�+�~�Y�9	z���{l9��12#5c��)b���7��=I1ݠ����x�{ug���n���T������j]u_E�[�8�N-��澻Eԁ�@t^F�׼H�~]o9AK�q�c)ol��ZB���&e5�eO�O���z�>�	���&n/�FB��[j�t�@����jC���Փz���Ykh�ˡK^Cw;�͵"��n�;:C���;���\�q��WX���X�cx[�3)�.�X�"�(a6�\�Z��ٌY�fK�K����J�U�Mc��v��eM�a��fb�+b��Z���:ٷ��V����!R�܇q����9�ٹ�<`�]H�|9�r�Q���4��ZC�݌�{�;Ul�c�3NK5��n�LT*��||0�b�2��N�u��7eHK�\"�8�4�b2"��d����Oi�|]��И���P�	�6��t��ʷ1�}s���=*�xxg��*),�������w2�]�3KR��y�;�c'!�y�ʓ��Hn쑮��{�%�d���'}���H����Y����(rׯ/(K�ӡ�m�]�D��
W3�3;�wܮV֗H�)Nכ�}w]-�w�4�x�W&d�\q�D�J�x�`��J���݂��w,Bjn;�~P��hpܬ%�p|��ʋY7�Y'C&��JT��_oU�c����`��T2L��)�s9#o��I���D�41��,:i�]�Ȫ��q�,v}t��E0��^�ws��o���p�`�Ҕ�{�\�1��3�]�(��à�Ƀntn��(K7�{�-ҳ�,����鲤!������b�Uu)�!������j�NpL��h�*	��e���j�ű�}���F��w:�:��Wl���1rt�I���j3�.��<�+��)��2���{�`Qcs8������_��Ѭ �\�ެ�Z0ޠԮ��+��h\5,x3�����������PJ�53w%�t��<Z�`�M���ʧ�X�dN�Ɔ���9��^8GR�d��e�f[-�|�pb3Q%]Ij�
c+�+�x�"o���@�9�����Y�h�~+:l����.��YjR��θ�ta��\�C�����Q�1U���b�U@mdan�u���kYI㙅������	�[Jf�t�������3� �w�#lr̗.�d����C��3�#Vt��HN}p˫V�X�\��d�νb��-wp�k��+%>ɝ�"��t�ԘI���x+�=z��.���8s
�x�kbr�.��z;|���'��ܳwg�y��1�C�k�}��������ş�w�p��']���c�)Z����_�'u���\�uǻ]6/wK����#Jwt��,b��$wi�GwQ�\3�\��T��\褧]�|_>:*
U4�Ҕ�^\<���A0e.nd�wK=�ǎ�.�����I���������uy�Q�5pѯ+�o*��v�E!�ŹnbwW4d����{E�+#��G#r��$��r�wr�s��y��M�+חM�W*L*4k�t(�-ˤh��7N�sW��� ��A  g�b	��OWk�6[%�j�&����+�%��6�AޯVF66�?>�������{�-���O��Z�ݲ[���[�������K��_�.j�s�u�o⾚�r�����Z�>��_����_o��������_լ���e�w�ު|罼�$AH�	o�~{rߊ��m�_=�j��o�����_�>֍��W�����~<*�wA��-��K����W������o����+�����o-�����������|}~��������j�����Fߧ���J���o��}*�.o�\>�yo�s_��>|ן�;W�;y\����k�����m�_��}����]��Ul�?}�Z�a���S]�i�0@�k����[�����k�Š��r��~{�~�~������^k�so��nno�����徕W6�����7�幾{��W-���m��{��k�r7��{����Wѳ~�r�i]�E�������'�������W��\�Fܴ|W�����_KF�k������}?�����_>|����v�U������W(#�As�?3�$� �!eC��8�����w0���? $?� |ЄG�_�}��|Z*��������ܿ���\���W��忊��o����k�O����ן��ѿ?���-��������%���"Nǐ��>��i��.j������l_J�k��o��o7��W�|[����[��[���W-������{���_�W/>+��ث���ƻ����J�o�r��v��ǿ����8:S*��}Y��|0��	"N������۔W�w�������5����+��?M������j�9W~��s~-矯�m�_�|���_�W-�z��k��5�}~����~����~����x�m��>� �@��?Q'�#�[���o�Uϋ���εʾ�/��Q_�������_��m�~~�|[����ڼ�|_�ӵ����h����uR����Q��l�>�fp�fg��d�$�Io��y����G+�������so���s}7�^U���A_ֹ~��W�_�+�����m�~=�����_����z�^W�n��m������^��S����w����B�x�Y�28B#���k�g7UE=&��������H�ݏ6�8.&�z1`m�Oh��yR7QĤ�pz�<a7"���rj�ߵ^ں�-٣�DW�a7$a�Z��8���[t3[f�2��:����];+ww�MY� ��� 4�ţ����o��~�����Z?�~������Z?^���W*��~_w��-�����]_��h��ܷڹ�)�t� �H���)j�p���a���������?k��m~�~�������W�\���V�}���m�W��꼪��u���m}����oګ����ϟ����}~��0eW�|�t@D�%����E�"�}=�m���yy������__=�Oż���}߮���������|Wƿ#��C�����iY}�\��+z�r�Q�ul������6P�q�T��>�c�}�;&�̝�Y�,����.��c������y�/v��¿\�O�xT�l��.�"��_}���3weѸ=�(���z=�Ke�����ѡo����g��X���=ʂY�(Fȃ�p��G>�w>��j6߯ӊ���6��7N��
��h��^"
^[75$�EZd׊��j6}M�=��ΟW�8�
�s�8���l����=�9�{yH�LP���B��HLvA=��*�]��)�D�ޯz[�'�FNĽ�O=��3O�X7�{�Lz�t$T?�l֮!�Va��ч@��]���O:�hOMz29v��.�	.è��^�:���u]L����,��J�ߵ'�r轶A��/��
]�+�����wz
�.����Z��_E���р\�kri����I+�"C�7�;�4�`���xa���U��(�{��/r�{9��ףq���F9�1�)�]��7`��oǏ�l�s��)�-�X1�߫�g�3���h�B_̓^����#®����J�ݫ��K�����ܞ��6~R���:���t"d*�'�/���+�ʋ^��n����RM��!����Fgf��DgA8��~�D���_1�j��&�����${니����څ`lu����@Cu�W̐�������o�{U����ݝ�[�<~�{ެ ���}Y7��l@�.�Q~^���&#��\	��ͧ$reW~�f8b�?c�߹����Q�:�"�H<D�����)ʗ�O�R	 )��x��]~P.�e���Y�X�=e�:�����98J��������kG �[ڦ��o�B��
�~���h�!B�+�NH��5�*/wL$a�&�qvg�r��f3�Uc؝�X���|l�^0z��� �9"�RtJ���]q������o�q�:4a1�ˮX���+6��Y��T��1�]:����f:E��5�����y��[b��J���̝]=�C+�w<����\кs��q��{��ʙ����J�}�/;N�(�h>hhQ��\�U_��b^��ޯi�|��J^�g��r��1T�|:-�3�kf�Mז�l�)�L�P1LKdyC�yC�<���v��ȷ���w��{=�[��ߍ~������y[��I�Fi���
;I��m_]�tnz�l��<>���Y9^�O2��bݹn��<'�p��'�a��|�;p\���Úz{��qͯ�y�+��T�ޮ�k"B�ر=Ny��MS�5���f�M�s�½/��WU����R�Iw��,y_
���G��ձr�ޚyp^U�#U��]4/$sȐ/8ޥ�/��K#;������Q)�v*I�	T-w'�nx֪�����U�Qom~1eɪז��,��1�G���@�V�r���gє���T�U�[�D������ԟ��G�	��C䤘��CPi���k��ڬ~��l.���ɧ����D{~q����S����v;{�vԃ(�[�k���"�2�k��������b�=2w��/܇��u����.���NmM��4MS
�i�:Ϫ?*��)9�{0��G���>��s���V)]y�.�1��_5W�\�`��A̬������U��=������9{D��ʷ�73�jX�T�=�����G��}�mPNwp�e���şs��P��9��>į-�`��X���GP��������:i_��>�]~��\4���z;���eX�UԠ���i�1^��c�ZȯPre��O����'�?t��6��Fe�������{�W7J��g��@��GQt�k�K��R�G'͗�&R�QB9�"ˑ�Zod��wN���ޯ1�#�Y��N��`M�HK)(f�!+�Æp�����Y�/�;��_�  �������@�>����7~����s��T��^9���y�,��T\^��ի�hꟊ��&���������4�}�2f;�gs�&�޽�A�n����R����\L��:M�Vw���`�s�>�]��Wef-��ު29n�{�!?^5_,6���_m-٣�� �y6Oz+^�J�Y����K��ޥ�1�H�����U�(��1~�Qٺ�K�cۖ}]zV�b����~�������~�_�-�'���'�?I�J�&7x3�y=�ֈ��U��>QW޿��m�^ġ����5s�b�����,.�;�R��bxa�;G__�}4��b���U�z���y;:� 8�U�$��������q*�/" /_z�e��1��t:shgz�e����/yuZ���Ⱦ $b2�7C�h�C&<y\f�G�&f>��EDG���Y�U؅h�.�Ks
�Zy'5�Y����q��u���-� G�^��=�����:�W�_�4�cՖ�p��"�fS�7=[%C��C�[�����UU
t��s��G��~�o�����ו�U���}*��bi-3f=\��Ѕ���w�{�$)\9�9
<=7�7�%�`���E��l}=���>WH(�鱵�dQ����j��@E����u�����t�J5�ftƔ%������.��5���	IBԢ*uh��}L�*�D�19-��W���nz��l�/���\v��wGp��S��]O�it��+���W}t����)-��a��N�ss���[�.s�����n��{��2�F1C�&d<���h�����O���h�����=3|�����_���Ng��>N��U���d��
���+l�v�u�dۢ���oo�K�O�.7����~N�h�!1�Sv��T�-�!�Y過�qh�\]{N5��٠�^����FJ��X݋�Gs��D�g�W�:�d�ߧ]7����t9$1�m��Wv�*�c���}]���J꿫����������Od�{*����+����.9i܄���d������U@�{Ŧ�廹Nq�u�o{���k͸G�W��^6���B�[����Z��7ہ��{p��3���M�rn�����DΡ5+����"��ȤZ��]k�ƶ;��`���)�)�w[�th^���՗ؕ���/Ȼ����ѷ�n�������L�0N�kE'��ߔ����r�V��ׅp������ԁ����"��R: ��|<o��<�����7syeZ
��<;�=�p���
��Y@�yfnR�:v���y.�{��{���#�]}!����N�Bɸ:���5�����ν�_D�k���Q8����`�AqL ą;���T����f[J���U���*�N��X�@Q�0��H��>�d�U�e��e��8z�J��J�=����=�X��x�蕂�N�N�a���xX��f=�c�U��㛈s��}U�UWg$R~�Vݿ����9��Ec�<}�tGM��|��
3�m���t�z�~Ƿ'��C�O����hϜ�������G���4[�>�~;�`�����2���{�s���C<ɴ����K����R�b�J~�KC���Y�G�zo\���
��<�2�=�#�H��3��y���k<��y�lw�t�ޥ������p�u9:�gU���lF%�Q�u�χ�zߖCѱ@��]{aR��˱4���Qr�}{t�-���f��ZsR]/z��(�y��w/z�����m�He>.�Խ�ڼ5\�Q.���
�^����_mv�Q��^cޣ�l ����ݠV�٧0C�:�׽&~����f���fA6�����TG�[���~{�%W��N�Y3��n�M\���Y�Z���XK{u�Z5�TĦ�T�Hg����br��/}%fp��k6�%�lN�X̢ۭ�W,��2�ج%vv�����Y/�ho5I�}����ܺ��~�X�E�$%�WrUu��Q|T2��e�7�A����%e�k��P-H�S�_I�r�����I�[ok����Q������<5�_��݈�W��+��
)����=�E��/���>��w��u�(��g���.{:�Ov+˱G/j�HD^�Ǥ��ޞ�Ϸɕ��X1_����&{�y�ҕ���==�J������?.�q^}��u2���=[7S���>�G��2}=ٱlW�ː��#�K�7�7�nms387�����oΐ<~��5Rf�ΞdW���/����v�w����1�}�g�q�e�{c��������r�UT��X67(�U7I�{�Y�Ѹ�iŞON��~���; ����D��h�1 �'/��-����A��}��/0���zӨ[8ux%�Z#O`����gtduh���|�;�Ї���?_<|���*��q(�p����o6k8�b�5t���t(vLt,Ǣ��]b��,�ҕ�Kb�7�k+`;9��]��] ƃ)��.���[�"�����ۘ8q�ō��Q:jM��u`��S�u��.�P۝�B���E�ge�vGF>�#�p��9+���b\N�V].�+eZT�A��j��`�&�0��r�](�ə�])�uaNkh�O��)Ky��i�Vɽ`4(�krr����7�s�p��h��(U�,�ך�h��{���s0��N�٣�c�q����Ff���c!�ǡ�Y��Q̸�J�+�����Lx�L!]v��j����v⽺��c���0����<k�����r�gU��8���<]���_\x�T�L�G0Ԩ��`PeMVm$�cngвR}�á��ѣN�t�DK��ww2"�F����WS	�`տ��n*��DR��M��j�O�h���[kh�<���.�*֕u6�`:w�er��T�R������źv�e�DC�CAbgvj�ҜW�2%�>�Ŏ@����N"AI�H�$a0�/�hW���{j�$_~@������gZ��/�S�K�o.�G�kHߺS�	�^�Z��Z0K	��=j[[$f��.�2�����D��>��dme� 3vn�]�W_bN�h:ή0�r�)���lǽ0�f����l�>��{�C���<&^�<�\t�\xoGy� ��Ǘ8%�W ���ie��g�t^�Z� ʏ�[l$��=����z3Q�ϋ��^q�e�GQ�-�\�GwcsRgWZ�8�sd�nw;n���̷q�W����\iX���3t0Ӑ0��M���`�2�G8�`�*���u�ff��P�v�̆���V���>�x
��2����2=o$����n]� (u����1�鳘"�%�ݎY��P�ette3>0*�M�qh�WX�ݳ]I@��yr�4��;[���x�V.𡻚��:�:��Ib}OsN��5yl����G��ݭ�m$#u�wt�p��f$�tp,.��ʑ
T�C,��֭�8J�{1�]���C����MALi_<1�B�]
�?[���
C�5�I4��b���4X��,�ϝ�Eb�4cF,EB`�,Z�r��&���#;�mF�:�[F+�M��=�2����0�H͋sk�3d�h�[�s\�ذ�6�TmL�F�1h��W��r�|W5���*1���CW5��%&��F�+ssQ�����r䖾�$ōE�d�-�vQF�j5$�V������� #������'���h��1���\��u`���T��S���;��ZR� ��#��pg:�Y�`8�����;\��ﾪ������$�P�����)� U����E��䗏+7��I����ޞ��%���2ϫ����ߨ��yo��xM��@�����?"�=���zs=�g5��Τf�[����jA�xR34�ch�Q���҇W{��N�xa�}ϻ��=��\)��d���Ou�q����hy����
8�Ю{����z�R�Ǟ�u���N�P��հ;�:�bTJݠ{j�)ƗY�E��a{|Ϲ��s��W���At*z���~�b��N�ʺ��P7z"�eK��ao1�F�W=0JF�(�~�jBN�~.��0Iڹ����p1����v�H��WB�l�MV�}{|"Ք���ԃ�!�+���=;+I\�Gc��*��~��3�?�P际"��h����W4$�R.�e�w#�!	ʶ����;iǶWS���Z5��/��?L��v�|��[������o�3��I]���p<��y[f�pV�@�ЭW;���F�u��}��}�|V7$�y��K�
G�w*?�PF������s	�c���oH�A�E��`ڸ�O�Ԅ�'�<<d��_������
;}���K�������Xc���e���5>��C���ݡG���]��¬}�f���wPG��.e���)�W��"�ɯ�Z�si���w6lEyt��E�����ޏ.����|�j8~��[��ߞ.�������v}�0=b������kZ�>�+^���Ƿ�'�=��Hv���6���)�l̪��~��i�Wޫ��=ů�d��o*�a�*��DJ�y+���M�E�5�|hVAZ�f�?oN{�j��JL��T>�Qe)��Q�F��{r��տ}�����#��\�)���>>�YX�v�]�k�te��=�n���<��"���}�N�Jռ�8U���c�R���m=�6����f�������Tiݳ;��q��C��g���8e�-���5�\�
c�ss��U� ,+��ܕo��.��z�m/��Ԩ�ha�fh���=�}b����i��9S��`����	��Q&4v��_�jm�E{���Rw>gM6~d����CAP(B�P�ɕ���n֨�k�>���ٴ�K�Nԝ*)r>�K�f��^f8^�˴���Q8�.��5=J�7�X�~�b�&�sք�V,n��@,O��Z�����نm�̯y��P�]�.+g����Ҷ��g���j:1_+׈u5���_�Ɵ,�B�tS�j�F(�B��Z�����c(.Ë}x�������Ƨ���S3W���^U�۟wA?yv��|)r�ܲ�eB���ޡ˻�|�إ���+��s8Ñ��[ܫ����on/�|�h2�c���Y{�>��ͥV�D̕|.]���\GR�zn�S�չ��R`��f{���u�S)�c�y�֙:Y7E:� �A��\Z�۝����"D.V�hP#�ﶿ�}�uד��cW�N*S}ѳa�a������{nE�W��rs���Ok��緂�J��qwǨQ��՞�������">��ub@{Hk�㷇�m�p�V�o����ܞ�8�_Zؒ��$=_E���M/�긏S�`k�～�o�}�qe�<��߈�dyw���;y"�O��B���X����:c���`M���}9
/�Q��)��V�̈}�r��'V�`����BG��^h��{%�cEr�9Τ��`���~�Ȑ���x����Sᚲy y�R��_H��΄�������n���csa�/?��к��M ���J|!�lZ���sww��t�</'��g8������*;�3�8-��F�/N� I�H�f7�m�?1}��!*=�!>j�,{1׺�?:�S������(��Q�n�3��A˶i},�#�A[��Q������ҥk~N��E��$��0���(-�����R��Kzݵ�e܏�����Q��������r�,�E��uލ�6�x����~U�5�W���rs97>�}��]g/��(by���G����{�]�L'y��������= �=�R���x��et��H{��(S�������(+��N�n�W�|�>��G#���ڰ!����ag����#�������mK~�a���}G�6�g��Ѵ>-)���+��v,�9�1�հ��}��n-^���m��<�vS��s����}HZ�Y�f���cU���*u�����Y�ۿJ����r�]��:)���#�b��~[���~>Y����Xٟ��o��7�w�۱����vu�v1�XU�΄ɪ��(��旇�/w[��d���7G��ًj����L~g�!��H<4�]J��3fD��o��÷vk��]q[�ΆA3��S�p �Ә���غ]gG�Ros9�H��e�H/��%��6�k8�y�/^�b����ʻ��������͟n�^�m`���}j���u����s���g�˵׋N�h��J���=�	�;M�����=^��>�9��v�,k���&��x̀��0��>n �O����3��+=W<��@���wz${�������P4�/1�V՗�=�����^K^��_�Lא��.�Mu�ג1u�an��t)p�51�xj�^˨������Z;��)�~ͫ���}3��1������A��/�ql>�:xX����{��S�W�_���P�Y�E}]+��?ԛ�A�n�c}�cṱ���{�6��oow�zҼ�}�<o[��X2�9vQ��|��Q}���p��8��*��OU�y�M�?z1"��y5kd��?5-�O�^_����+��潣���v�˸m�E�~:��xY��טe$��"�Չ�3y]�:��Y������M������T�l֋��U�n�l��4&Թ}Y�u�?u�L�;��*�F�d�G-Nr#���}�W�tlv��}�k_�_^g+�!�ܿ+������ۛ]�m*XUm�����ISv�W�=�b��G$�~:��>���)��*���1//T-c��h���˨��������f��ch�R����ٷ_9�|��?9^�2�*��l���SKl�^��};�u,ܾ�~�7��x۰�\�i(Ȯ��|��4���S}��z�~���F[���/e���i����ˈU+�V,t��wW1�] f�y�t�� $'�r[������E��`����G���K���S�]�UtU/e�%�=��bӽ��jy�W��׬cl|�����;_8|���!�[�Ң>	zW�R�]F,�蚚a3�}Y���;P^�`��$ڳ��X�u�h�a<6�[7�r��k���.�O{�z5�v�Ec�ӡ�0p��[A,�+3+�·q�/ј&�@�j�3c�:Gv�681.C���/;1��{b��J.�c��y��}_W��}����,�AO����Vuq�5�MO����q@{�K�d���Z{���b�4!������U̮]&UէF�KVk�0�r���g.�Q-�o��aT=<�y�n��dWU�����#�:Q������C^U_v
Y�|�XW���ƚ~�|�ﰾ�����R�Դ}���w�(e{�O+D~���_z�}7�V�N�^-���s��R+9��Bx��	� N�4�;Գ�oO�6�V��2��hv���/��x�w�7�_ۑ4~V����wd� �����Q�S�g��}�"�M��J:��Y޻�xM�{;�:g�Q��
E!�+o�������{GxL���;*Օ	Dw��3m+3�n�v�9">����9�=�㾞���5�g�+˾��#��e��g�W�Sa� 3yty{�q(�Er���y1,z��}�� �L���@�J�U�9�)�ێ�@��� ,'VS'�\kF<^� �k�L��&b��w�(�Y�7���3��ha��ӵv7����^�������n¬�? ��Y���7��ʠ�+��C)����J^�u���'ޞ_�dX�i7 �A�[�Q��W?\u=�����+àd_�(4J�zwú�%%3/�k��lD��[H����E�Oo	S�˻+��R�K�����Ȅ�R�uja��*��Y۾�;��^�״#�=	ahk)5'��1j̨�ut�igq�zg_��.ݸ�a��2���o"�U@��y����7ߧl1�����گ�W�o���z�{� �d���bU}����k/�zn߶��
E��)s�HO�|8��Z�HǳʆC����HM�������f�e��P��y�hu���7�rֱ�뫻_v�myj]����Vx4%��zn�b_a��\��.�Cf��E<Μ�U��zڱ����&6i��1hDЩ;J���V��9�FG���`�;=���w{���3S���p�4E��}q�$=kz����͚8��djoD��{�z�%�]���W�_UU_97??����-���Պ��ܯr:���R5��2�Si[��_���ΰ�c�}KG��O8ㆱ���ze�~�z�%���鈵G}}��/=��~�/�
�]p����}�����jWݢ�{�đ�G}��������	O^�tV�<�]��ɮ�A���w�w�;�=ʦ!=���[��u�+���g����T!m�"4l�L�P�|�9�=��ա�I����_���r:����-�����F���>������V/>x�v}��O�i�;�3��+\D_�к�Wr���jm-��ֿj��<U�Wt=?�/�w��Fz������TO��z�|�����j6�a�U�WH�U���n�����}u���I�o��t����~����I�0P�uw���H�wZ@���{��s�n��3z��;7�[h��t��
��Y"�}s�����§X�Fq�7yf|�9PŃ0)�l!�K�`V���`Y̺v�� �Ø�S�̻��}���ҝ�cG�o� ckۊ�u��z�Q�5䌘d��CQ̂9�~��!Eq��ZOm�e�$����wbɺ�ب������f�f�S�-�"�_u�QXˮ1�E%+��8��=4� *d&�R�=j^Ӆ�£���L�H�Mw��}��]�ؔ�r�!�$x��{p�{xi��N�t�3~�Egt��늬�a��[�d�����yL�
�c 9x�1�O��^�2��n�8��eM�/:G�IvOP��a�3>�6s<�e_v��X�6�:v��gl|ݵk���qmd��ykffR{�=c�����c�)�Sn�pf]���+5���)���+"��"0� �01��᢮S�G�>��1����C�V*i��WaNNљ���n5GyQY���	/D"��f�f�ޥ[݂���]�5@�C/B:ʇ�����{w��A��4B��S"��JY�I�Merܥ�}���2����īw�飫sN�,��w*��o�oۏ�9Sg,��Aͺtâ-�:t@WR;�S�#ٷ���S�.����Tx��5�T99Y75�M��S���$se�s;�n��N �3O\κ߮�8ju�%�J-VŖFK\T���C������K�[N���,}=C�Ҝ���>H]���.��t^F(̣y�^��L�v�	�����c�`�܆��إA�ˣ.�aS����M�ዳ1u���*�6��g�]���`�6�	L%�sԠb:��K�Ό!Ľ@���#]~.�[���ǘ�	�fs�V�݉y}���428=f�C����#��̽ά�3v�Kz�+:h��m�Z���K��FΙ��[)����þ.S�q���5i�.�p4μ���f�cݩ鐲ю�Yu��Vh̙��W{��Czˀb���V�pe�N;�r�&cK�d�3e�C(^$8<���:��yƀ�0Um��~����}�������_ῷ���ƍQo���ɷ�[���ہP`�����5b#lF�m��QF�T�Q-�kATX�X�b*B���A�r�b���+�ۖ���-�#m��cQb�(��Ab-�4��F�� �X��s;��Q���汱c�j-�llVKh���-yZ�ʮE�`	�A�QG8}�&���zV��|q��@�uhL��)����lU8^М0&W���;��W���}��y��>��Ǉ�z��������VP�����s7��d}�3zo��tN�m���J�mz�����f�J#���2��Z�N��zU��r����S$�[]2��sQ���Vn�ԗ��彗=X"�}[�k,Mbߟot�ȵ]�j��I�k�N�:q��`��O�K:����}ڣ!�6�/�����Ej��^U:*J�������
�;Nm�r���ݾ��\}�͍����~�j���7�	K �T8�5�ۛO�9+*�T���=v��NFnFнj�����a�ݖ��>�)����K��>�JF��{�܉|Gu��	�p؏�E�u��"s����P��<��4�W77��y!_��y�eY �gV����x�)f��ˣH���'}��+��`0�ov�O�+�F�WK�4����,6�tކ��1�Wz�b����q����w�Z�^�U}_UPԟhє����V�c�vq*����@����)mČ��7��
��o������������������3G����h?eg/�K�����KO�s�����Ց5��s}
�u{�:_^Oi;��S�<v=�� �Uc{f�m[1����}��Y��!3�{�~�z^���Y���D�bͱ2Ws�{C~�	�ޮ=+����{>c}�I��;�!���t�C_�����1�k^��WT�:�{�Xx��sH���+�q^�{��l?��g޻=���ϝ?,�߼�s��[�+)�{٩z?���ӧP�U���`п�VYCV���߻E�y�=�����L��_�����<�z��T��Yڷ˨�rdD|�+�=瞪�҃�wBb:�n�1����/r5G^@gc:΄ai9J�=����}�_��J�ҡ!m�5��[y�d�-Y�H�5����/*[���s`��V]oW>N͹�l�5��Na8�ɑefVʽ�l�s'��Í$/i91(��?���O9BF���Ջ���ݪ�j�����K�l%gFLF_FhX��n��uXK��ʍ��Y_N�m���4��>�����k��J_���w�w��Mn°ѸU܍c.{w�m��3̹���J�ݴU��ݳ�C���yPL3;l���U��{#����=�N��=?TH롢��l�鈹���/�+:Ǚ�S��|oy[B�jP7g��yw���v�x�~iYظ����^/J~յ� ��������{�Q�ы|�h,Vb���ʺ��T�.��x�+�Q�F`�M�JF�p���js�����sڵᾔ����;s��w;�C/��Ez��z�`�'�Ӭ�u(�ǏV�H�3�����j�.-[q��c�0��)?_�߽�A*��(=��'����[du��,RN� ��̥J\�8k�*�MR��բ�v���.vdJ�d3��s��|>z�s}ܤ�+�K���8�%�;�*��_�3տc��kӾ����ٳ˓鞦��2��i����uu�7�e�CC؛	��ov?T�O�c��z~��e�^�`�C���DW��#�~�q��w���o��5�g�s;҇�IKʰ>��P�vug��7~<"s��/�<������k������BBѹ�Q;�5o��}�-@=S�׭ߝE�A)������eϡ��.�`J�6y�ĭ��r�^I�D�%�����~�)���i����2Z�e����hG��{��Q�V���lL%_�_��##�����>�B�Y꼾����雇�0fE��y％�x�=��wt:'���Z���&�,Jˁ�ؙ��!(�m^�y��o�2���c���"������yfq�VX2J"�n�����My��X������͸*�n��Z�ׁ�(I7����.����ӳ���C/2�8����U���n����B>�[��+��_�c_Bs�0۸�t^N���3u�ţ5��L�i��|��i/�\[�g���5YѦ������y�L?X���X/$p���yg���
G��3)g��Nt���b^�k�x�G�)��j��~����O<^ڱ3�Y�*���B޾�;�Mp�Zkç�{��C'��2g�)N���-�%[��r}�˸�2;�k�Z%v�}j�F]����T���aH�W�����ޓ𭏺�����+���^���V��>B^Oֹ北"���ῼ�%-�}�s��Nv�^)�}:�0�w�6L	յp�?Dz���U��I�=I{�q�:H-O}����҂�����_w�O���s9�����h���5�3v��V���ѸL(���28!l^��nN0N$�V�i�U�mX⮝�"��� ۘR2�!��-��b���3�������ﾯ�o�)�{o{U1u�M!��g�%@�\ES�o�gc͎�j��kՉ_���w�R�m��oR�M}[�ې�	}�v.��D�����\�n��i#��ԋ*M�%��SVf~��?8���j�I^�\����k:(h�|�#^��{�5��R~�+�4n���rE�����{T>gp��U�=�~�����-gԝ(��%�{,�ӆ+~�i�3��<'B���K������� ����Ս�V�{�`��;�f���7OǷ��;��Ɂ1�\Rp�'tr��\��ں�=�Ќ�F{��],�9�ǥ	�+8XV�P��xOa�f�FQx\i�g4v�9z���z
��½C8xhz�&y��8���}�z��4�~��jC3��Q�_,��~��T��0+����VƷ3w��Z�v�Z�W�n"�a($�<:;�S%~c�n��gr	-i�MB��B�Y�m�k!r��E�S�v��e��]b��w;B4*a�歝J�B�彎v35�@�p#�������ڥ�{�_z�zľ5��N��ީ����G�AI�q�V��Wt�Xζ}�r��w���/7=������C�?3�ߣ
V�5+�ܣ�j�����Nu�����l������l����B�G��K�W�ۯ~HGٯ~ޑz�/��*���'Exv�;���~�Iw[�o�W��r�N�m����>�s��i\��Ŀ|L%�7[�x�/W�V�_Z��gձ�ٕ�~���j?@��9f��c~ͭ�t/z瀐{����=��_Jn������=�?8��k�%��8R�M��%S���wW��������*�N����ǅi�]	R��|W�\��������0�h��1Z{9uA����>Ԯ($;R��l�C���7(��_�0M�*�}�"9c���u��eS�M�#�Ғ����f}%�)�w^C�-2pb$�8)'oz&��g ���p���;lU��y>{+���ꪪ�}�=�{%�M��CW�h �4m��n�(�����{�;���N����ዾQ�%WEqm��=%� ��o�no_*H�]p��k��#9�Е���}`�-�ˠ���}�w{V���%�Cd��ͥ���O�G�o�6.���R�,��Ɯ�n��"��C�����ڟ��ӨN�OE��4��n�Z�y��s[���^��/Oה�㈱�+��;;gw{��sv�P�C���T9t��T�lyw��ME�MO�9���Է߷��k�c(�m�ȵ{0[Sܦ��)�|2�dj��ޝM�����UaI���-S/�uy����n�r�wX������^ߦ�R�k�~�fΧ��R�����������I��7�5�Hx�b�(���U��v��m�YQp�tۣ��5��+�蚔�IF�^���v� �/2nv�� ��bc(c�v8w[W+�@�l����PZ�R�������	��n�������xI��🽾~m[5�j�"^�wz�]-�_o.�m��A�h�;~?�VU�ݷX��v���!g7�z���c7�E�O�lM!f~B�˼�Q�C�m�����U���͹��Q���Ԡl5�vG@��Fߧ��>�w�[�s
p���ug�p;~z�j�K��������3�K;���(O�DM�4�z�n#����/�a��^�wZ=~���U������G���٫��=��c�JU��di�6�9�j���2���`��[9�	��\מYc������d��ܲB
} {�4,�g{x<������~α��E�BA?z��d��ޡ�9˰��u���5}���T{w�P�nt U.�����*JE92Y}pd�C;���+�Nu]�����Γ�է5�,�H�9o�e�g�`����C�BS�:�j���຀���1�:��x�t̬w���^������UVa��O���ݗ�͔�J���S)ΙG\ܦ��>���ˑI�Y��u����\&ߜ\o�W"���?J~��4�����V�Y��шr�v�QS<��\)��>s�f��S�ͯ/m8��@\q�pd��V��|x��d~إ���.X��>������ϳpz~x�^V��n���?�ڃ�ܮ�_z��'���T��Q�,tcw���MGg�wY��}bＮ}����*�?p��ڭ���/��]!���
��)Ph���T�[�Sy���X�_;�,B�����\w|y�r��p=�]���;������yFy��s�_MeH������-޼���xH���^��|��B>�]�5�s���W�d�L�)4��,�	)���F�eHLP(#��$ ���	�`a7K�+/B?k�6Q#�Kͻ�9��M"��)[�[
Ƃ^i��ʻmu�j`���ˢ跟mQ��A�9���Nʻ價�Ցm��&�95������Q�t�k,ml���X�s�>.�]̔���|��&k�l��N�t
\ۘa��üV�V�ekv9����zE��P����gG��P��m��@�W؍ˌj4)W�E*!��D�a���O��1�,������>�,76�t����"/
]Z��j��a�5���v��ٜwn��r�B "gk����O+4���z�p�0�w�P���t��! f^����[P��6
�
�3\��e�n�*{Q`��E$&V�o�_C[J�[z��:k"�jl�t꾻�|.
5.�Y5�9YR8Ҳ5;�-�7g����9�]��j�����Ǘ2�ut��K��]p6��wT�֌����+���!�C�����Ft�;j��+��-s]z�
�R�:��k�n��V���Vg�}�/jY��hnx�q���W�]���`�"ō�]Z{NI��坳5ʨj��6��#Rd�����o(黷���rB�
aз3T��U�	ߊ馇"Wt5��x�������&!a �iD
JDLF�����Z9M�����Ϩu�*^�[V�h�N+��gC��+zA��D֩]�X^~g8D)p��P��h��l�v�m���n��dL�gS<`7N��;@�4"i�VN��A�Aզi$3V��+��g�����0d�3�Z��6��Rɦ6��w7Gs$���E�ǙlWP�%I=/���A��d�u�ݹ%�vFP�%��j����䙹O�7��_��H����0d�l���EnN>��q�V1W����h��2n"��u;3T�К����i�s[����sVt��٦�ٛ��������ۺ��p�'	���������ҩ�)k+(�'�V�,��.H:��#��j2n�ɝŃ̢��7�n�p���> T���o���cTڍr�6���]�K�٧�hV�OT�;���j5��K�1\l��5D�|�A������2]&�b�+�,S��,�=I��.�>���°$�دB��u��_㫨zF{FukV�V�>޴���$v��[���m�x�ᩓ��0!����|�2�,�K�u�k�GX�]�I�
y���jRRB^+o{�����Y���E��F5`��Q�U[��sV�m�j�yjlc�EE���,UF�Q�Kch�r��b�"�X��n\�sm��A�����k˥Ƌ_���F�ւ��X6��hѴ���*1�yrѷ�ʢ*ow[E�b�/6-Ci�?
D�I�6M�GC�ݶl����@���
W�ե���Ag0�#�
�r��T�DT����p(8���/��`@L��ɾ�d�5�el�Е|P���.�k����T�껸��W�Ľ�5�7�<�?���e���+���0���Ig�~�s��]p���!��@��Q�4@4�s]�G�����^���z�-&~���W��y�2.q��Ǹ��%cWz�W��\����,wH.�<�p�ړ!q������J����>�hu/�b��({{F*�Z��NήT]1�3��<��#}���ӎED��(J�r������S}�]��h{��]�;����$%�S�W��z�No[ϼ��w?]��5�]Ѱv�&��MO3򟳿Gu<���+��~�G8�-m�;�z��}2�|��Cc�������z�ц�~;�g˨�d��@�����vz���{�c�=�^|Vۻ�mǖ".s����J�*T{��ڼ*'鎻;�WR{��F(4kUq��)���V��w\�Boa�W�EW�[�ɪ}�Z�����p=�j���:�8��� �� ��%�eZ���]�)���¤[DD���S�1זS��i��I�I)�N��!���q�:���:U�n�WZ��m�uZ�����GJQ�A� ����~]��6n���S�=�z�ڑ������JAB��j��w�W�ݺ���z�ǵ�M|�+�.~�8TWH��k&'�ĕ�mՊn	�ߒ"�ԛ��3r��ɫ��k>�:^^����P�Y���y���=ʾ�& ��N�gyq܄����t���KS��&���`U�\�i$���8Ы����<�[�����T�f�E'�ةt���F��=�)��?�3軟�V���z���#삗E+@�fnu�cÆ����<�D&�*�ƥ�ޕ#�v�r�e��#�GIW����v	D��$���m�)87��;2�@����Xy+G���Z�c�y�>E���zބ���(O߾�뾽��[�v~OJ�k����vmt��w�$��Y*��gq���%��[�B�jͷ�-ͭ�H���]� �E{�;+����S3\���{2y���u6^_x֡��>�Ԉ�a��t;��W�1Ǐ��_č�>�i
�J�j��:�F:��(�3�0��I��k)��E7�S�W�0����<TT����քn��O�Ǆ�S�~��	���Jj����N�q����������3�WU�K�H��-��WI��X,�D޺�ȇ7���r`��P�͐m���~��{ ��B-��ng�䝯mUg���F�3�CC(ƥc���(������vW����Yu~��Z<b�@r�pd����y����Q���������Y��[�#Z2�p;����PL�B��©ʈ�n�c| �2
�<��2��%Gq�8��+��p�|���1��BAZ,��Vo6���=�'Imᾧ�Nܕ*v�)g��_To����nY��T�
��+���M�(m��N�{߿D����.~�ݻ����;64-�*#�I�'������ȍ!��S����k�T��^
�ۄ�B�Fz�h��:�&�{�M���{��M������b��}�k��t�~��P���R�yo�����W0�ٕ�������/L���;㺏��	������*o�=i���]3ʬ�M�7����^j�@����kD�����]�7�:���M)K}��=���~K�u}�����1�/��M��O�߿:&����zq�d�I�V���d��s�����nm8�<ş_�s/ΞPů��g�o�_Muޫ�Mnu�D�Uz���q톶���eep5bG�!�����]�	�]�4�Y/6��:9�i�@�i���d�n�Ir`�|��H&�h���D�[����sx6�
Cu�j�й&�f�V`w�����}Bu��/����}��F�����<ӗ����>�����^_��1��
�b�I�^�uס��z�F�]�C�a�\�Y�C�'��<����=�:���et�`mwC6%o@�Ў��b���W�����[.��+9���.>`�X�(kB�}�%��9�U�8�"䦏g�;�s7��w�/P=@��[�*.X��7d����f���{�p��l<�l�7�e�[ڵ}6�|������y'��;0�c�{������g�l٥z���o{|�9���T�/b�s#�C=AJ
g���c`A��藺k��L��Ǿ�n\륺�.������ת-�Q�{����V�YOQs�����/s�������cu[g�ld'�P��c|Nf�6b㻝�
i�6J�䱐oM���pC!�3p%��
�e�}x�q�;G����d�P���^��KB'�VĪf�u:ڧƠ�R�UU�9/OD�~�����}�<7��3�u"q��ֳ!D�������Ð�^ݪ���T�
G�V�ݩ�xʃ���k5f_;���ͼ]��Nr���o�}��U+���})��B�5�����!��>�'�ڧq[����ŷ[0޻����X�PCˊ����G��:�IOh�Y��Vl#�~�m�B�]��t���<d�}���� �=�O�B"7HuUpUPs��N;!WM�WS������_OW=\����U�Q��uo�藷�ȿx�8��8��f=����J���Ρ�l-jl�L�z�s��i.��=k/�xs)����|\����&sz�mߺ��@�����j�o���VbEr���W"�t.��WѴ%ڬ�����/�ī!��#C3e����!�Nq%����k�n���T��L[eJ4bI���b�2�R�"���̍ՙŎ���*PK������m������`N���>��۾�x��������9_T����dA�o��W�pj|�R��O��ݒl;�)�qY��l��ś_Z���c�=´V��N-�跧��鎟��P��F5y�h��X�����8�9�Y�Z��K�|�"��5�>�6��-¬J���{(���Eα��gM��I�S�l��ӓ��U{�{�}:���������~�s��2�AW�p�{�\���sM()=���W]�=�ޛ�ǌ.F�d�QS� �KM|����W��V�K�,��~y�f�2��<�*-8d��CYuJ���}�|"�[��|uGU羥��S��5����9jt8�|��ŋl��ȝY���m�����_)��i$z�����>�hy��07��|�/t��{~\U�@u���=�#��-I�Qު;3n�O�J�m�vv�JuʖV)W=Qw3P֎yjpI�� Er�gr�#�ϋ�we=��{}0+��l<�ևm򒪿�����%�z�̠�:�L[T
e��nD�����!��3������z��of�_p��_�]�T�&���P��o�3��3�kv��y�9�ׂ�ʡ��1	�����@�=9ʩ�����_S��G�wf����$����X�����/��L2}.��}�$���ӎa��_���߯:�U������E�q�� �qUR�W���N_������\vA�_{�ީ���)�nq]���1P����hV��Z��腧FLe׽W�^��>�y�8���d�h�+��Wm��	���&�����y�PX3���/Fy��^o���CYy��u�߽�U��]��(��t߁W7��y�\�^8}�-�Ņ����Lؿd�{�{� \�'T��x�[ﳭ�:d
�Ŗe5�h\�s�A?0�MF؃b�9�V.]BnkT�0+Uw
c�:�OM�ȣSit��U�Ɲ�׻�3_��>��~�.�V4jn�����C���B��4�z�{=��U������WN�ͧ�Ԡ=��J�ߏ�P�S|p�z��.�/�&�{%3�Tԗ�1���ݴ뇔�}p7hё�m��r�{�9�!j��vUy�{��S�t*����pz����d޴_�A��'�kَ�$�@>ɯ)V�FX�ߍXOO��~�K�BvO-�7�u6�EEw�Y�� ��>w�~�|�{p=C����'��,�r�B���cú�\�"&���YW�����^���ju�����B;R�Q���Y\�K!0b��d�{��dz:qj�מ0��w�6���
�JO/�hP[E<ּ3�W�����-��K��vtMeC����/i2��m�zL�z7�7z�"L�"��#�4K�]�,�Om;���]�܅\km)�7�M�tY��׊�H�%/�ܖ�V�{Vm�%r����4HjkN�Pf��@2om(�D�n%���D���Ro��9Nc�pg��g�J������y�t��d��p��SĻ{�o����k:�	�B�}�#ۆ|���"��U��d�璇�XW-��Yc9�웜�Iy��HA_� LY��>�+7u�!W7}��19���c�,lL�s�l���;�r��zo9u]Ru�C.�ժ�y/]T��N#e�A�T;ň���}�v�]�qPj���y���i'7:'���97��ɮu�eJ���QYV�`�<�,k����luCOr��Ğ�<Q��7�|3����b��K�M{(Y�j���������޼�9|�I����U�F�bb�T5����"�������e����i��yO�#�Ґ�����������h���pd���Q;T&H3�	��/�i.�c�}��&��ǢY��z�����I�Ԟ�7� A6 �9�ނ�q�㲳*E%������ٓz�&+u���]��J�8B��֫Dމ�F�5��e^hiW_sW5�sY��GU�x*��j�oW�ޓ��N[��+��]�r,�Bu�����g*V�?��dkإ<'S�Q������7;;w�Ti�WY}���rR}�I2슒��؇4ᛢ���֫=���l@��{%I����,(^Q�Y*���[�ƥ-A�U[�8�|��J�
U�NV�H�wnW9�9bqu��)	]n]��^N�^�5:T��V�V:]~����B%fm�¥�j��ޜ�0�1�玭���,h��;������os�y.B�_�ތ-Au2�=�Y�Sޡݠb���/��)`ޚ��wgKɎ����M=�k�ss[����-�
��&��!YJ��.]p�:3��AY�ې����x�QJ_51O{��z�
=��v��0�	�:�SiΣݯ���Y��ydu���j�5�7"Pӡ*��ق�'vvA�dŎ���/�ή��nt��6�n[�m�s)�y�=���*z*%��4��$2��F�5�����D?Բ}���B�"�a}tw~�	Nv���
���Z2X'r�Ɇy�[A d���V0.����W�J�MҾ������MfV�E�#���ՠN�5��	y��c�c�e͉�v��t���8�mA}���L�#S�4�������e��K��}��i�S9��2mU���
̬��v�\
lYR��.�F�tr�R��bЕ�}� Y�[nʡ�B�ĂP]����8|#$�}�9��	���|��$q�o�3�Q�Ή����b�4��;2�:�Q�{)3z*f�w,J�A:��7����"������f�ɛB3J�ɦ>wuċo�^�HRO�;����2��^��j�q��N��!�u%Brs�-�Ez�oZ�|�--H�vn72L�@�Ǎ:60ن�h�vT��[�X0v𚫑m��uI�.
n	��72��!b�%L±>�)����qn?�R��As��ϋԅ��s�����+��b��b�XڋO����ȯ��Qo6��o5�sb��\-�m���6�v�ˑ*�k5\�*��Z66(�\�ndǚ�p�E����Y,V��6�*�k��<�n�,Z�`���(��-s\��b�����]�m��ۦ�h�A�6"5�7���ԅ�Ds�H�O��~t9�,�~6�k�OU��t�N�W7�-�t�-⫸v��j��z�����ޟ�T�M^�����ҿ/�^�-�A1��+�=>@�GǮG���O��1�����m���f>�+,/VP��T~�yuw�dn��Rb�f6����EVUb�8��>ACn�b��Z���ş��i.��S�]O�w~�si�:�޺�c�{�?l?s+��^
�O?-�j���k��uvIS�^�����闹��xs�!�؜a�і=U����N��0�O�		SZNyuR1�h[���)6<*�* �+W���r�	g��U�k�M� ������x}g�c�=I�c���3��v�_6/�M��қ��r���gK���%�uڏ����[��Cܽ�O���w�d�h$ו_g�n�Ԃ.ŋ�szhE	��"�yX��q��׫\���}����a�v}�Sg>N�0v�VU�ͥO�fβ�6�>9�fa�e��+1S��R��OӶ�`!^W��Xl�i�����gVH.�i��j��RV��bX�>�82]�ٕ����d�9Y��;ow�N��򇐞���׵�(W��_,��Fh���<����>U�ڌ���@iR��۽;�Q݅�9T/��'�uQ}kV�hZ�����~�S�F����L��FG�w����뫨el{��ھB���ZY����׫˗��c�5x�J��ez���zuu[��6��K.�����W-�.V��_��)��9�緫ψ��@ټ�J��yX�;��}폇�s�pi���N�:���5ݓW�B�cݗ���8���>�L ��B_1�ƙu7���m=�H�Ƈ):��}��l��f=J/z�;��;��V���Q������
�>N����g���p���􍜴;�r�g�<�zǨ�_�x���~���b~�b�K�`� +b۹]�!P�V{��T$�׆T� ��:���?z?o�`���nrê���d�c2l���V'PBv{���Ә��F�U����/SC9Z�f�m�g����U�#��;��K�v��(�?ʣ[�J�����'�~=��)\�+��~�=k��4-���^����:s}�t�
Xs�;Ç�\���к�����ݽ+N���5��禢�O`/������X�y[�ʜ�$�OjU�����S�y�Ցu�^B���p�w�9tj�>�({�{��ܹ�Yh.H�X^�8߾�p�����&���+O]�<�[�7j~���ڠ�f�]N�\ua3�������{��m��-l�u���uj�ժz��ݗQO����
�h�v��C\D�r���������z~8\]����M͘t�No�Wǖ@ٸG.!�?O�}��˃�t'#�;.cWO�^nc��g���[�x���g8��^����B��Zꂶ/K]J�q-�w챍xL	-&��/ʝ/�e��e񭼃d3X�f(��K ��I�N�3���C)5[���YDN�S��CK>)�n��G�@�<k([Ӡ�/���v�n%�+���d/<�����h��s��<���@��>�c
�Zg�[�'�==�����>ޚ�o��$��d���QY������zk��j�K
��(��9��~�����.6��'�X
%w#7<�����eg���S��;��˷2�n���SYv>�t�3�1˜��.hdצc�뭝�W���pC[�v�kp��{�qs�s`8{�|+��f�)���'�����~^3�$1��>�n݄���������˗��O{#�+|��AF��7>�GUv�XB�����f��/�j�wK�\Ϲ}E�b|Z��Җ���y��r���{=���Of��8b����WVtu��s�y��_�>���2=6_����ڟa���J�ݵK��߮�3W�(�K|�%k��&�NVqWa<���]�"�r���h�r�C��)�v��B��z�v�h�]���<��m!���(a�(�����SfSi
��'��r��Ij���VQ����ߎ��a�o3��o�}������楻}-�]R�W�u��V��B�xn�;��m4;w:5]�S9x�6��ݮ�^�t5��x�үΰP�<&�ߔ��N>~��I��Rz������ ��_(�p�ﻳ��f��{=Ƒ��U��W������ׅ+q��3�ko+��Z;GUj�L{��f�R�����T�\�μn�"�{]*�����@sQ����
�L�8����R��Fm|c*��(�[���7cR��B���cr��4/��g��R�K��f�Z���ug72��>�?"�}3Y/u�aE����Cl�����~�=*�߾Y�!>��Y�w�/���י�Fp��JB�ԧ�G�Y��fy�?(k��~�<`i�]p�K7�a�V(�	�;��@�&*U|K۝��t�mu#�j�[°�W��a���V� ����{�`p�Sb���NV���c{���T�j4�)k8�tâ+�,_m�t��T�OWn�6���V��F��u�}�@V!y��郎�ъ�t�+E�E�n�O�f�;�<�Y#X��9 A^��7��Y�Q1p�<
��w�S�s�/��Yo�q�Ҏ���F?vU?���MϷ����O�����������Szj����'���hƤno����1�q����My����|����p�{�.�1�����*+/�_{.X�h{�I�T�"J+��T�lj��Z[���:t��FN5�E<�<|���������g�[��3�crf�=6�����zkn˸����=��͌B���.A������+Ry���N"~	�4�.NE�a� ��[� �_A��f���_zC���KGgvx�KJhQ�0b7R���'[�t&9��	�����N�i�f�E@6 0�B1�	�:��I���n	�����B+���1�e9{�@Rs/&q1�Id��SGU��G;"x@*���B�3�EM���[M=H]7yx^��\U��pb�svm��t~>Gd��a���^Ԋڶg�a�m����Vk��S����ԣ�����-J�5�����nI�~}i�������}_z
��O�����O��y^w.��?�)��)�=�#<��j��^�*n�Q�w8���g)�m// �������=<7�����s�䣫PJ�(��o�X���A���vx-u���$���D��eׯ{��?O�O2gxoǲ~�=F���:}��#3��OrL׹%=�z��S9���H1�GqzuV�j�պ8\�1�,����㏽�������(�i>�Wp>��j���O��m�}���kw�B��oq�uA�V�!�M�]�������\�yyA�X�h����b0��%�X���c�@y���D�5���,c�,8�����N�cQ���{]s�t�m��s��zaB����e�V�Y铪�lc�p�0\�Ҿʹ0n�b�˹�B���JW����Vwj����_�g?c��NZT���eOBϱ��Bm����V��uX�Gɡ3G�w�E���ι
ҡz��l��GDP[�o۵h����)��T�C��|2^mO5�IҠ{Ǥ�j�;��g���C�'�C�Du�
��1�C��={�JQp��o�����l���.R:�ahUz"��(N�n����^���g�u{g��x
�B�;ڦ+�]&Vxd�aΓ��^fn��k鏮�$[�rc̮AgD����/��L�� ��]�q������V��
[ �J�H�T���<aG{*o#=�c��~�N>�������zz�:��{ep{s��z�!6=꿽j�+]zMt缬WQ>��~7@
Z�e+�A�{ӻ�!W��u?^{��s'w1�"�#�Tﴌ�MZ�^��I�r�������ٝ�@:���Gx��Iy�<��Lb�4C��X��o�v�y�{>�ا��� [F�e�\�u�^ؼ�H�d}��}��uUA7)z���+x�Kv�[��L�`>jg��wiW���im���̪B<��-5������������z������*�e�@�5�<����{��ә���'�J~�U�8���������:B
=�tM@���ҩ������|�ϔ�E�)Ӎ8�*��o_��t�F���_�cϭ���u�rN����]g�ןB!���1:�G�Ťm�e�k�D��{=S��pMS�bba��K��s:o��^�; ������Y;�<R���v�wlyJ��WA��H��c(n{j���k{�}������ƪR+���Ġ���^��!*�1Qf�)�^�B�3��F��R��}�����G@eu줧!lVM�6���A�6��v�NS�L�*�-�{_E���46k�v�7�KU�S�Q�d����Z,&۴��Cb��]�	�7ԝ=�ӝ�Gg��W���ɶٞ�ׂ�T8�^�8+��bv;���}=^bg���e�?�VC��w��={(� �����5� �Kh��c��������E��_v�-��P�$(�@����R�d�]X8�+��F����
gzӷ��U�,�x��Y��^�W�`��j�r������#�#�+1nb�=�7�yR��1T�9U:����陽�OEk�iX�˥t^�R��^��=u�nP~�[pw�Ly��~�[��n�þM��~��jh:g�(f���[���OOet~�x=�4�	F�N�L�����S��m��p�29�m��?G��~�}����EQ��|�Uh�*�?�-fy����ݬ��O��������0~�8��܅�,��(�HJ�A1�Q�(C��ğ�ϩ���xid͍��#j�>@>G2�ڕ;���}x�r����[xqZ�YL��pꭵ��;�P��X9B�M^��J�́k.�}��N:�Yz������<)]R��im�j��0�s5N�4i���˨��a���(���o�SCe[91m��^Rn���-�%w���K�j[]�â4�b�OY��DM�0fT-����&H�d��-�ب�i��}�C2X��J�+���r��+o^�\�o��i�8��:�\��wRu��	ǔ��_h��n��1-��+Z�B��"����t�)VX��3��k����"����X{mB~��%e��Ud����$N�[#|�&L�e��Ab�k�B�n���M�ݲ��P��t�����i		��f�P�$f�E�s�j�;��>[K�eI����w:�O#m�!F�!V~��n}:T�ӏG_K�����K��d���X�Ig
Ѩ8%A�>Ax1��Q�����W��m�����&A�c�ӷٛt�Э���(���{>]���e����Y��^gQ1L�d;o�CՒ���[=ɇq8��P�c
V��K@b�N�\�ꙺs�AP=��Z��b ��iaI(Yp"�nĜ.9D�,�ٌ"� �˪�2N���J�y��+���:���Cc��]G��O�Z�m����jC�E�/��n�@k���0d���u�	����vծ��?O�177�o<�����!�E�7I�[W@YX1B��w��{:�3)�S�m�$ �hW3��d����/n6���Ve��|�:b�D�R�vA��O�c�FA�M����h�|Fۊ��C|�|�ncŝ
y3]M8z�.�е�(�H�[������X��ܬ�u*.2�s��QÔ���L�[MS	��w]���Z�i��M�4�\ª���,�[{J��6��+��b���u���T&f[k��tcљL]�#����\�:�u;Fu�$o)F�$��tL�O�u�{�J'^w@0�#V�1{w��Y�Տ���d����Գo��-���L��</f�v�DY���}2�.�tjsQo�&�VH4�]��u������4��D[����(c3'4�&�S�Ѳ�����W��]o�q
�'%���ĉ��a���ـ"�8�ʖޢ-��Σ�a��gpl��G(���VY��o0�G
�:9��r���6�*���{��0H|y}o6_h���o
�@�Y�s��r�sn��k��ߦ���6�ۛ��P&Ж�9�lb|o**�v����&�-r��r�5;��F,��-�\܊��yF��܍_;���Et�� �+��\�h���_�yk�v�xnW64Z5s��v�.c\�c7(�<ůK�wsb����v��*G� ��5�.����#��!88漙\��̔f�`��E�pp;.d��V���}_W�=�Yz"|��f���?�iN?c�3�>V��H��O�ׂ~�h�`�_�^N^����/��~�=Sc�z��|�� ����(��.�����*w�v�in?p�����O;V���;�K�o:y�]����w�����Q�Mr��Ӿ5z^N"B6V//h�I������Ͻ�Mg+do��>�=U#�nﻪ.WT7��_�c���s�1�3�l�޼�a=��fz�����5���ٖ�K��C��aȰ�
a�Yr%��0�����b �?�>���.���o�W]��%LoC1;�
v��o�P5�_D�p�դ�>�sꁌ�R���a�H�P�?U�]������=�N<�OB,�&��=R"ugfUm�[���5�%�֩�!�Se��W���7���f�������=��W�5����4���B��k��yk�U�&��f���m"�,�]s&��g"u�a@��z��j�M�zͷ�B��+,Z�ݎ3r��G5�N�!���Q�@�-,l��}�M=�Go�����uWk��tv�ZޢȆ8?ϫ�����������Y��:�;/�	�����@�F��9"�7�ds�0/s�t��1UЙ��)D|>؀9NrI�5��,��$^�
�e@�yn����VtuSK�򰾩�ჷ�o��تG�]D�Yf���=���%����(d=ុ��/8�}�f2a��4v��i�j(��W$���u]��U^f���nq��i�\�P����V��d�q�B#=�����>|�qy��*
�,�����l#�;^|Sl��
=���c��+�=�G =�wO�C'��Zz��p�eW�;y1�Ωm�ݍ�m|�ķ�7���W[���<|&_{���}��+�8�F��I��?/X_H�|��(�<�bv ��U�s���󁓫�sp�A��tJ��Ǩ<w1�K���8�$��件�1~��}Mtm�g��dY�D��2;aL�sےd.s�P����`�Տ�ni�媧�M@�f+�ټ7��?=���_�y�:9�%�w!�$]��)i
C]��"���6ba�w)L�J����ko2��Wcx������%���R{+���  8]�Q�5'Yt+宋��D����r+��s��ym�ʝ�k,>,{Ҷ	
�uY���>����ʏ|&j$(q���Q} �O7v���y�E��ѮF`�S�O��Q�w��,8LDP��'e�>ǣ*�i�s|y���r4�_w�/O��2W�Л��V��d��QC�}2�ej��^����G��������齋����B�j`�����9�¸�zkb����̜����y�]�c?)��]g����9V��r�f��W'۵�8���Ca9�-�=^a?Oz4�G�h�>�l�[����*�J;�*�W�>g������~�B���L^�s�~&�b��T���탋�~0 .!W<>����Ui\�5����ǖ������\F�ޱ4<�[$ȧ:��@��#����W��=���_�O�xi��Y�]\E��M8�Rm*.>�0f3��u\��Xɵ�V{��|p�
�ڿG���ʉ��X���-U�ܝӘ�\�������`/qu�x�=��X��Q��ˮP:�Z���v1�aV#9��1pͥ�er�c2�\�t�Aʀ�H)���[>�ʘ�ܫ���D��o��S
�c���R�,��*C���7�r�����J=T�Q���ra\�
B*�q�]J7a+�0/愷���CG0���=�gz*�W
��b�t�q�nYV��b-zE�NyUqD�펯�MA%r����3���нq��{��H�[B��7fWU9�Y��U.a4��N8�$Gf��c\������U;ǫ�����@E�Sju�5�n��)Wb�OR���LcI�����,�Ci���P����L{�9󽪚�76���x��h�کQgN(Q�!�/���%H���H���D���v���r!+�M^�|a�|�ÆA�Ι�Q��5�\�v7�O�<��sٮ��yL_T����,g�_W����>B�ퟘԥ��t�>��7��������Vd�-
圷9���6�l�%��<������9�����۫~��c�(ZT-ZǷ�W�i�J���3]���>�F��F^���C�6d[tr���x�h��A�h����!�6���=�}��3���ZxA_t&���.��Ob;t�WeI��P���fv�?��Fޝ:�����^٦�R]�O�VGF���_����7�0vmq^��A�s���e[k��	W��>�0�-���EK�<uWļs��ݬΩ3�h��:�:���>=��f�6+$vB7��itJ)>��Ɠ4��yNH��Һ�ǫ~7��^}c�&��:1�ê(��O����j,l�!m�U۬��d³�y�Ҭ����Q�k>vEo��b����͞;l>�Sܟ�{�W�;�G����U'*e�
�:]�H������S��˯z3�O*�񋨍�nME���v;v��\��A��«��
N�ȅѷ���� �q��F����.H�X/�k��~�}x�\X*��\A���;��N2�q^�N��91\!��:��V���	�Bs,����08*NnI��zA�<r�~�2)L!�p3;9l���Wk��:L{�Gl5D�1��.TG�O�Ir������i����%��ύ���%w]�-	A��8����^է9�� 5��O(����l����̨�3iҷAI�e=Q�q���,��HX5�'$�6��a9�K�\j�9�*|��������RQ�������� R�a��U_t�9�ԦYA9�R���9��||,j���5����of�:�͝��&϶<bte?:v�S�;���S42&U�6F�y��J���%�	�}�֣J���i��U��ϫg�`s���M���sc:%ͯ8{^��v���g�|s~CT��*�H����!�E������΄��ZTJ{�ﾾs�V9�r���{3)��1Y��.9t?H=I_ә1���JI��{ݪϟ�P��T5�<��(ßnI)t��
e��8�8d���i�9�}�S^Zu@�;��E��w�|rׇ[��:h�7�$�n~"��V��~���g��|'������l?������_���ܹ���}����3K*�y�R#��w�QAʢW���\r�k|g���"�g����%�kZ	�xM�u���3�x����=���Et�9�}Ls�G�JC(vм�$�[Y���9x�C�*�9�)V��n<�_��1���}���A��.�i��ٵܥ�3k�{��b_C�V���nn6�uAw�U�7���Ⱥ��z����k�#�Ω��U]�e���T�	��*����'{[(����}��(]�9���r3S�s�<z��w�K|�x��T�T�UJb�R\"|c�D�
�Ӣ݈ʃ�y9���W�	G��S��e�AN	�k�5Μ���%t\B9
����c�����}���de����z����; �RM�02	f����7T*^�]f�\s����vT��}C�8���,�ƕ�t�@�Pdcr\#���P���gk���/�1*�z���
��B�B�UF&���r��q铷�kn����*���Q%v�B���j���kW���~>�*���[/Fꈌ��l�/lm�̆ܧ�Q�a�|��[,�[$��MFH�^��J��,�eGL\�rO��9r�1Uz\�AE8b�P�p2BJ�u�(�Qke�y���~Kʝd0=������΂�_���k�G��t���Y8?P����n2 OpE}U�Gs��YuC|`���Y:���0��Np�˔�6�Qu��Z�+u>���*�I�$dЪ����G��uLr�2!c����/f68Zk1�������gL�����;�v�1��e��f�1��r_B��%P�f��H]��P�ٺ�KK�ۛ���~�f���"��R��.<�����ey�8��J<x���{\��}�ٛ�܍c�/�����/>��o�����.���~�O�p��7Y�\����˸��W����ܞ7�"Ϝi�tҌ���q>Vf.��.o�|>Ϻ ���s�"�K;ΰ�Gz}{6iR��*�>u���o��HL���`򞟆{���E�a�ד�E\��t%�ȅ��ٹ���(~��8K+wTP�W�H��N�v��=:h%�����a*�0yyF�� y�C��������%�Fs�K�l)�(��A�HO����(ND�*��F�/)>Ƣ=��%�}5ʻV�KޠL�jb���t�5C����S�1�j�lt,M�<aoS�g�s�5�I-	Ǆt��i���x4tm����	�c�"qO���?&��L{�p*�~ؙoja{&�Ugm�E���~}��,���ɴ�䇞��Ӓ��})��8 D���Rj�֖�L!w�iB���'\$���X��7F
�s�<�W[�&:ه
�o;j�U ���X[��w��#�|>�8�6�O�+0�D2����P�	T4Ќ�sb��5^�
���|����ӥD?B&~�V�J$�9��0G���,�G��1:k���������#sX���w�d#x�1A� ��.܂���ȅ�����RI�������EC�Q��Mz�݌뉓�e�I���a�����������_�}gY��8����s"}Tٿ\�B�ϜP�Ӽ6`���B�o��r������j0��|7$�M��8z(&(��A����7�*��d�Zʿ��V�����=��ѥ��9��L�s��]���:P���κ_m}����53�/�A�3�b�b�C�Z��1SI��Uʇ���T��O�Dч���R��y���װ���+�й��*�O���f�a�������N��\�j_TӼ���+[^�B�̆ �gvf��P(Z�+ y���2Ϗ�%7��_��9d)ي�b�-�!O]M�NKoi�au��M��{>�{��Q�EɃ�n�6�e��:�ֹ:dLˮ!v�D7�mNf>�.k�g�=N���V�R{.m�;V���g+2�E���3�@�qc�B��˓�}��#�%ڥ.>��d>��/�ݵ3����*<�^K_�].�D�NLه�R��0p�"���WގQv`uÕM��Lq�m�M��?���ί�"4�q,���O7RO}=D�0x�$�UL^{�B]_O��[��ĺq������J�$Ï|���
��c�J�t��[81�������au>:�J�J�jf�^���s0�RbY��YA���L(�s�mC&�c��>���?U��LC9JlѳF����ˠ�z���ή�����s�ӳ�������IDP���1ꡐi����?��Oǜ�+^S$e�/^�,w��[K���-�2E��Q�mB�+�2��[YЛ]�oޠϳ�\��բ�D�59��tp��#�9��:Y�9)��n`�|��8B>ɑ��S�'�C;�پ��O��je�1��w�Z���*�S�F䒩ub�33"���H��C pL��7�?˩]_΂�-M�����u��+1ޑa��h�Q��g�h��57�Z}�]�����`a�V��C֊�E�������Nڍ�J��a�ri�2�����
9�EHԲ�Y�A�wIp>�+T�[��e���{��EQ��q�������A��X�� OP��y�pj��5̬Ҧ��!N:�M^�RA����9��{2�յ=(k�Vذ����'o�:pr �ܱk��e��}��Mt��eh$�#e�­ח���:(;3Dv@�}Z�&���5�>�Ӊ�]�0Z��ov����q���`��*n�C/V^Җ��`%ð����ۣ�c���dkڡw���J9�\�)�#]K�[�恮��s�txP.�k]�	f3�*oG�v��6�������q���ݨ�ˏI.J��_.���5�����`!�8P���6���}�\
���UڹZd�gh�r��wN��{DD�k�؏�E�gq�ٳ�zխ�)��)qZ!F�s��h��䓏X������k�5�Ք����U���Q1���=�x�ѴY���.����St��%Y}d���;��6�d�|�Q�.y�e�>�	�H�\��y�g���]�a��t�
�Vn_7��RVq:��!��"ޥP��y��P�,�Sa����6�V�-�n�+��͋�e�`�+(;��ԩ(�c��� iJ�0�bj�3/&gj{��96e��H]!���e���,S}���	MD.�I�8޾,(�Q��Ȓi�u�O��I��miμn���B&�������N�D�_�M�x�VT���[���0�4jC����T�MI5�`5]4�Խ���P��97z���ה��v�q��Y�u��nM��� 	E�Wjf�Rо��!�@do6����auC���0�W�� }�j�t�\��G�6�Һ�꛶�Jwjn����ǅV��2p���/i��n�0�`,\6� �Ӌr+Z9�Gh��Hv�h���m��w���q�/l͡E���y2�������3a�Yg���M�u.�J-�U �2��py�R[�С(wA�v��h�f��%^&j�L�jZ�kn�wf7x��ۉ8��}M�=����h�S(�~hN�x(���~?Q�U���]��n�t6�ѱ����6�ͣ�nlD^��ng��k\Ǻ�{����v���\�\.��w]�mE3��-�^^U�=���c���Aos���+�\��o�_>{����r�wv�������[��W6��[��^h�Yݮ���\ѮA���.V�wlo�;*�yp�.nF.[��{�ޅF屃X��W�r�4UΛWwr�g��NV����-aU�4�!ȸ�0POh-�.��eq"�T��:��w���*�P1Y��s��S��b���ϟ�3qx�C���?od�~����p�����f=���y�	�S�X������ã��s�Ek�	�n�nZV9�yh�-OQ=���dӤ� \?����^�5AoW��Շ��Z�0�Z�qR�i=�`B�� ɹ�B���N@�t	�Ӻ_/�q��|���ldF�=W(��XI���� 7ا�P+'p�vD�T�~5���wB�s�9�~��#������j"çGЎ@�>�%���]r�g؝}~^:��5�W@s��'�A���t"~�v���%ld �|yU��K�5�oe��R6IsS��fk3G�zU@��6&;SrL�`��هj����b�_��?O�(��� R�i�󨏤y�M�qt4���z�i���Zo��k;@�bJ�D�4B���G�qD���,�Ν#B$�������{��S~w�D�t�X�f�2=����:�fKd��25ty۩�����k���ݮ̦��n:�����q��s0��p��l��z���o,Q���֪�X�˧�&e�@����;��%��D�-ě���?W��}�M]UŇ	�_��iT����`˳��v��$����Fl
Q��v�#j���*'LVę��Q�iޟD�B�>{_`�!�8���h3�I�㈷9�3MP�WPl�Ӆ���;k���~Z���O���Hc�J�.�yX3[�eWFoM�6l��3�.��5���7r���u�g����x�q��=����c�fy��	�����y�_d�
��F��g�+a������O��o����Ds�]ǟ�ns1���,����2w�oz�7��fJ��sϾT-p��.q�"cqOn��)�6�M��E�NtП��x����D�/�5�����}��ڸ���/:C���[~�<YΛw�5�(�r����?J�zb��A�����Vu��j�0�=���r6�З"�<�FT�IU)��눊�}l��Z��-��QO�G��<����Jm��w˲a�w��)�u���H��}�.i���3S:�D�L�$��b�f�D>!�hQv�V�[���\�L�����W��J�L�d�ds�b��*�wi<��9�Ȫ�h����Zt�K��;���G�y�C�DKR����xy�{g�7{�ņ3U�K�=��"��S�L�!I(�Y��|z�쎣^����.�1�t)�����>*G]��B�uPg�"�G;�i���<�Aa�Q_rjɗmƈ�F�'��3a�¬�4�
��c9m2�7]>�Y�k�-P�1�LÊP�8Q��O�L�mH���t�U{�pb&�_z������ȿ�8���L�;�x&%i�qC\� 9f|�D�)[��`�����1��p�r*�N��VE�E�R,yޔNr�g�ڐlt��P�ȏmʉ�n-��rCVEa��բ}�r��
��-�d�À�>�:|I�r��>eZrX�"b�en�zO�8d&��_Y��t�ȅ�Az+�H�G�h��,�:��-��ާ�X�G��|�vh�ޙ#m���uK<��b�r��׉�VY�}v�.�CXʖ��`�u���k�dh���K���Ŋ�s'��ha�+UΎ��d>۲v�Mw,�D��Z�=�lGx��U>Z�H`ʶy�o7�P�����Nto*jܩu;�����%��w�$?�*��-@�W���_m�����}>�tɾ�~�6G����>���	�j���1��-�C�Z����2��_s'�;mK�ו��7��Fx�͈���k�:��j�O��;"
ރ��Q�_]*��;nDɔ�T��6Pr%�Z���T���-N�y#��M���p�?`�S�Q���/͙�c�Jc�CLzr��!q;h==��]�év�K��s��9�{<�����P�C��ʏ�P�}�����}�P��Ʊ��^��ߍ���N��5����J��Ϣ8꿢Q'h7Z^'PL)'A��/���=Ʊǵ�M�Uu�_#��BZ���d*UF�nI��E2�&|�Nb神.*�����J�s�Y�ư:l��أ�1�Ҧ������R�0]ǂ�e�������.^-X?~��?��tz"�QTϔQ��f�t�19!�T�3}*����iӘ��Hc��&���`���>;�0��4�V���s���ټ�i&�4ثIX6��(��$����e���Ǝ}�O����iй��]D�DS��`h��6���5/A�fJ֭8�u�q{.A�.�F��Ռiq8���>���/�+��?��T�����/���&��gQ���N����U�C+�7��-J>���4_�or|�I|��,8õ�ȕӆ��9.��S����*8����c��Z�;i��,�G�*��p�@Ή��dm�*�V0�������ީY���X���7�B�x��×�ߏ�lS���C�A����8w�}TT5jQ{�XMF�p��2ec�Vv=:x�'�W�s΁{���V�s�@�1,��B{��w�5��^O�Џ�f�$F�Y��^>���Z����?j�lo�����s����ن=�
=�և���گQ��ռ�/��Qӑb4�?k��(w׊�D��Ƭ������� �ޏsz�@�;$:���a����]H�UR��ԗߤOG�� 7�u �'(�Y=tph��N���n�� ��t����H7$oWP����\���}L�� �d�\���{��q��]����*�Ѵw̢�S�1�w%��F���@�9lm�Ӧ������5��O[%��O�����,��U�q�R�p�#w�G����w�������D��/	AFh���_7'������t������L�fy-��&���8�Ee��
��6��O�<z�j H�*��r�ȱ-���ݜ�ʡ���Nu���<�jA!ڛ�r�g(
j�?o{#��yګ�S�:�ג�aLz!�9��'4k�`����d��{�GD�˼��b�wSK�s膥�]4�8/��A���8���yt�{��n="���O���<����q�s�Tp�mO��|w��qN7���Zr#wX�����}�(���C<��Dƌz{����1JU��7̏(1?��Ϡ/_�5�{�/����ˡ騔�x������+vU�@ej�o��{�z ���4k}:R���v��3���FP^��h{�}q�G��P���0W�yP��=�m-�1bb �,#5L�
r�{?y|��K#�������kTJ��;T�n�ʷ��;|�'5�Q��N�&[��,O�@UJ���YVr�cm��7�g,��l��҆LX��b��ȧ݋�k}wϦb�q�����s�~��q����?g+�����`�l��2+���N�x���3C��a��G��EC���"t�}�7:\Ze�_�����r<&$�c�z8��dښ�F(t��}�}Ӆ��Eʐ��T�D��;b�5d�#�ZϷ�y{�ΦNe��7F8�BϽ,�^P�W�ȅy}��Q������L��B)J�Y����X�<\t�Xd+O�Vd/�5�j�[�l6g�]����xv�MA&��a�ɀ�(:��/��О&H��y�.�ޮv�C�̹鳤�t	\�P*g���_uWʤ��:�zm;>��^ޤ��
��ޘߢ��y�ǡ�*��j��g��;�#�^�]��k3}z2�{'��z�{�B�oGM���Y��Y�9���j������;��Y���8h۹͎Q���i�}�(�����8��$D�q�!]�r�ǔ�����n3�6�[x�j�s�>���4�q%gmz���d�69�Χq���[KO����St��#�NP���m���9���ү9���vcw�kmU���v�_�8-�7���r�dXP���3�yX4!ې}��u��[���[+s{��o1_�ɉ:0�V�Zd�-	^y��N}��o6x�U�:y�}��^�za��;Џ(�4wa���.��#�SJ~0~�`�)4,�=��}ύ�4�H^���@���Q�_v[����ug�����>?����_toz��F� ��x�GV���>�etH����wp���[�^5�I�`�{�V������Q�P��gqӪ��7@Yxy^�J�GW�粅�j��W��"�2j�1W:}q�<��z�UƛӘ6�-��p���jl=3����bFn��)���3dU�2Ջ�u�cu3�]�>���?���S�[�O��~Pw��\{*O���q��Q���"��:���q骟W�nAu}j�6��8��]%�9���'�z�ھ�~��;Gם�I�R�9�6�+P���P�e��-;v��e1�ܝ)+�F���G:Ռx��)(OQ�j^-q�zu�Y1�SIݙ9��B+كpH��}7"ԡ�eI����sK�D3x�d��s�|��Q��7�%���,��=V�",���iz��!��&�I�`������q�Z�k�K�3�F8��CΨ��0���s�0`��qZ[2�0)ɲ☮P��PC#s�+�O�F=6�a1�)�W�<�νU�r�����
?�-G�L�>��l�l����e����yy��풽��g
sܲ����v�ح�52�f>"{Ia�sK\�����4��r�@,��ݮ7�4x-����0�+��e�q&�e���[�H�YU��ߗ�O��#�3����9��"ܦ�Z�;���N�vT�0_/������+�q~�q�z�X�y46e���CM땪G�
�Y�S��䒯B����o�߆����[�R_!���|�+��ߎj��,�\fD���{W���k��PiŅS�w*�w�3�>��X�l:8d�a���]���J�Z��V>?�O�!�3��MW41k�,�oj�\81�t�9I1����Oz�R��M�w^>����;;k4k��Fʭ� YΏ�j�Bfwe��G��#ݼ93��v%�Ӄ���)yU�1�'[�d��"�(&�r����D@�5+�-�����o2�s&ˍ��L���i�2�I]7
xXن�A)w�ɭ�8�}��r�����9�����x�[�Δj�+��Hߊv.��wIb���_��i��z��R�?j����C����k�X��͘��b��.~��]֑���x|�F����W�oś
���|��ܞT�tA��|�����dW ��Fr���=���
K𯎿�)�(���V
iE* hz�Ú��Vy�/{o_$K����ڨ(Ǯ��Re����bF�����"��.�������t��q'�r	��K5�R�. <��d*��t�ws4��Lع[���1e�뫍�}U=VC���8�+8�ЏEρQG^�d��(=�w�;�H����z'>�T<���a�8'~�}����V�5�h�_�B?�M �2���D�ƚiH�l�R �lG��
_�*�$���H��A�ulIb�'+t�F��th��۬]�Q%#՝bS�I|��2:A��閪ܠ��϶[崹�R�nI��'7 �z�v�5�uшW,`/a�R
J2��ut�f%�sBV�Z�CR�
�ܿ��ʽN8�{WOڮ,o�+|�Vq��k�e��8��4!�B�R�"�II�2����,	Eh�`ٶ��'op<:�ڋ:S[�,
ڛw�t�j��B�k��5إL�Yt���*Mu�<޿M�b�mV;3�����![��Nս/�����S��f��z�˵qF觰�y@^h�}to�$��8,�!ы�;��gŗ��]v9�n���7[���9�r�s�ӝ�&E�8^�T���]��^��=��n��K�9OKw`�d�&�љ�Z4:k��[R&0�+]�_B���|\�ՙcM�#Ւ�{����ϼ���=��v��.���n�EO��՜Ik��݆K:�S����Li�	"]�޼3gJ�2蓧�7ְ�X��V���wU����2</m큅���`\bm[����C����RG�񜂂Z��D�钲�Cҕ�fCcq���"��e����n����Q�P�x	VK9۝�S��qu5�/��B@��!f#���BK��h���q�)�8����	X�ߏf���S{�T��_%4���,�ި-X!�4N"Z���w5�A�H�\v�F�+d�2�ע�5Yc.a; kf�]�ˤ�|%06���j&�IYA���f���O��k-���^oS
io��+�A�!��H!u�gV���ل�7��'�F���1�Q>�hӵ����$Eoe$O2��z��R;w�zC��wNe?A������.)� �b�}o���<�vO��Y��kǙ��4�AG���W��p�Qwas����ɘ��<��ѩo
+�狩�D_m�����^S.�\�4� _���A��{���pլ#��呙u�ˡ�s:M�{�ae��U�0jn z�LٺVQE��4�����0�v�	��`)kF��ul/N�fb�V�����Bk4�Dg;�ȫ��V)WٔeK�%�^L8t�q��\�J�!��U1����܏y-J�W$����B���߶�I!D+��/r�e�w���a_���˕�{�G�N��'������E�nF�ۚ�W.;�&Ms\�d���m"1��G�<������uʈ�����H{����#nh�u���ۚ��wcnnr۹ɻ�$7ǖ�N��j�nrӥ�|[�<�wr�\�l��M�����<� �csr �H���7�����^�hy��;������yo/97�h��� �����%����>v�]t%D�ܻ�n�����\r��;���'v�H�H$٤"9���H@ݾ>�m���W���f&�kL�e�/a�.�՛�a���vk;p+��s{����	d����t����˞��>������I:�g��qa�ĕ�{���z���=tm�E���T�_u_��#���aڲ�+C(�E�M�.I��zUn�u��니�0�Pˏ(����!�+2Ul�F�^�o]y��ovP7��<�:^��R��~�xn�2c7�ngI��u@�nyE��g����o?*�)�o����~�l;ܯ�0��G��z�%���R��&�~G�y+����/��1�9��սBo���s��M�>��Q���Q��O�btc��^���k�M��B������.Fϕx����ٵ��I˘l�ǎ)��z�\���n�������*C#}���:{�
�S�%�ȅyD���.!�+��@��Y�9���=Ӓ�}�?���O���	cP>��	4��W2���fh��SN_�WE�Q#ĺ�aթ�$��6 ,��"D��j��8>�`锵;�dZ^��������Uc���4��nC9�3��T�OүOVͨO��W��=j�'��fR
ˬ�c��Z�r��c��H��,a���+#nأMWw=�B��pW֋r~��U�L�`�[�K�sq`�����ջ_u)���vu�Ƽ]Gz���ƺ8١�dgD(ϓ�y�Hn�w�\���Πb��]o��}�5��~C˺���W�'$'R�t�8E�p�H��0]��3z3̈�����P@2Ŗ#e�Qg*��Q�E�V��0Q'�C�����I!Y~�z9�|��	�#:hEȩ����2x�E���g����I��v�]q�k69M�s�rXy"%u}�Q4l/Ld�of�
�os�9����D�o���2��[i{��tIw���\���FXhW���3�7k�"��W��%G��g2��]�WS�aT�}|�v��w8mC�((�A씪p�\H���"Qq�л����y�~����y��[�]6��׶�9(�@��G_I2�n{��<���X��w§�4K�(R/o?��tߐ��1Gx���0[p����[�~�=�Q�� ���:q᪆�)��H~6�w�g/m�r.�����;p�N��h��n�V�����:7�Ok��.��x��X#�]�E\Gi	�B�d�R*��[��S�w�{�J9E�z}OJ���;�����;��̟f�t�_��3��.�!��	�r�_�催��O���O�Z���Q��je�*��G8�J��;����̾|��`�ؕ�>(��T4�J�X�q$�Y"t�eW��t�������8áx�mq������|D�ʒ�0�z��!�lX3Y�����3B��Ւ��+��U�ݞ�t��c�lS0ܪ�}t��`����Q'k��O��ܓ$��}n�C�?V�vx�@%��;������#��wdns�c`2��蘟#z�Z��m�說O.��SOJ<L�}^ܳ���zQtꃠ�cdRbYX�@3d5j��d�PP=�#���~s�E�~9_tٚ�6k6Y�����;�d��v*Բۮ�+X;��Q%����DM��Ί�9fu�g�z�#=>c�9��{+l����[��7���
Qn$�����l���$tƍ�pw|:��YU�H�#
���tp�%�㠭��l�7��P���H���l�.C�?g��ݢw��06�Y������Cq��ٯ�7�77/97�#�W���{����zI󽠏�U!�6�;�D��W����k�{�nn��+���\?+���Pw@c`]�ȏ9ё�x�!��:���}QfyNo�_pwJ�ծ9:Z���!����s�]�{<�o�T
��_l�މ8�9�<}]>u�LS�����P���Mln�魺�&jw��|��ļ?:�co�pt�J����Av{^��w����;���L�\&J�@l뺖{��w���mx�7M�h�.񑣵�R*���R���4;�U��-M�r��D7;�+w�m���'F��:-�G;��y�q�;���e:	7�K��O-������^�Y�M��p�7�p1�<��9BZ�0���v9f�˘Y��uWG����P�}����l��xr����N��}o�����Q�I;bkF�A��{�!oUlA�?B{����s%5�/�ز��,]��U ��	"$K��GX��qU;�]�[�u���+�.���l��yS�^�VA\l:���z�^��x(d�ܾo���jn\u�6l��B��t:���T�N��q�cw���i�pi6{���`�N���NCSD��6r6���������+e�U��{ �5��j_Hh����`�i֦�ڵ�q�<�P�o������V��f�Y���J;h8誯y{�Ԧ m��'a���r	LC>D��C�Y���~����S*���M����k���D8ߔ8�CfJ)Ĝ��.�Uƣ$,����t���}��\�~ꬌ����ę�2݋q��f\X5q���&����EL"���r��K�>6��:�LYD�:z2/���6���T5Ō�ﾲ�w�:ع�o%ru��DŜ�a�o�k�W�E��%Ez$��+},���dƞ)�{V(�O�I�����Z��������P�LϜS�����𙋚Υ]�W�O���ƩE�g�rE򟮀�>r��ޥM�,G�!?W��#���?t���7���\KÔ�T8��Y��U��4e�+��)3�{�E���ݵ{�z���h�sމ�	F�p��ޡ}��,�nt��T_A���g`G��i{�~̪�Y�j�Hi&�gҟ�%	;tj�ƥly{H��Y������j\I�M��Y��Z�^9Y��__�"�ą,v�+y�0F\w��w�O�O/�L��ڢ�7��)��Dm�Ζg�7؅S�z��l�lV�G�r^�v������;�O5{;\p�[��~�~>ļ������֌{����:cK������ʱ���b@���4��-�>��=+�>l��y��
��1�)�D���7nj* ��@�PHW�u"{��1K4�X{Zҕ����Ƥ�3�Qb#�IɔO�n�p��޽&`u�������K��L����ݵX�G�;�����u�Jr>���{�Hn
rO8�e�f�c7}�����4qzx���-P���r)�sT���1�a��eX.Aβ4�������O�_״4��7�g�_d�P����w��D�JQ$�'��;;�
�����x7H��Q06�NEȪ'��k"�/9��L�bS����<�����8��X�,PnxmW�;�ez,���5�B��y�"o�kȉ���ub	1j_������M��*$���A[͝�EC���k�Iq�qOj���h[K��-�/Ysmo!�3���YDZ]����:q��AǴ�x`��Ú�2[f���kp ���`Y��ᘺ�Ҭ]E���v��: ��3{��6ڭ�s�l�9���<��;���UIz`��G�g~I��z�;h�!�����w�Ԕ}c]	�)@�ǯo>�*���=p}FW���x���?T�$�Z���W���}o��nzݭ�߭��9������0����ϒ�,���A=���	���5zl�`l�]n��w�����A��(x�=�w�q���~s����JܪJQ5Y�:}q��� ����X��y+^����q^���ʨ�'�G�W6O�e8��2G�ab�����n�\e�>�Q�szj�UԄyJ����94�L���Ze.َ-�̄�k·���.�A�F�K0ۡ�V�&h�>�/�s��n�H��nU�2�C���.���)䮋�UEL�E,�I��"�ƀ�2V�"�^y�/o�W�	�07����{�1U�::g�3��2{�M2�Pp��YE�b�=�"�~����w'�}{ZD9�:q��S�
�����Ml�VXQ�J�М��s6�t�S=_F�3�e>��ާ],:/�S���8���D�/�[_K�x��k�lϮQV����K��k�C��%7r���m�(��s��V��!�~����裂*4g���N\�\��V�8k߭��?�P��5�"y�"��"WLf�b����-�������#��c���ꕇ-�L��T2}ҋD�3�h��/��(����l�}ޡ}�/�y�gnwTk�U�$�PG��Q�q���p��D�8hweAǞnk��A���Ŭ���vs�.9�= ��΅��f����BGzy��к��O��{�\ڭ�ك]��O��(��?[�b�zjT
3�~<���X>��)R�
	��w_�>�[�W����Fr����n���Q�B;�(��Gx�I�V��cs|�]84}��z�g��ܻ��#��a;� �#�Dթ���������7o}勱���g�==��7N�|��֫�;�>zI���0����1�?߾K��ہ[�;�|�* d�Ij��4W`z�1$�޲å��'ڃ�iǜ�s���/^���]s�N�&� ��OEDd��ED#�6�ｼe9=��a�����6����V�cYO�4�q*�v��W�5�]�^U����������q�y#���F�ύdaWQ���(���h�wz7�hz4\^-�}�N�6Q��׆�������t��>�½}A�(ܰ��������.�#ܹ��yq����S�(��1-���e7Ѡ�:��C�K�g}�<���7�O�1_��W�d������(G�`����x��HX��b�F��oDW���h�!�%s�1fz�|"�,��o�R�����k�k;Q1���A�.((���@��}�����nԫ�(D���[����d�|3�e9Pi~��QU/�-�]ĝ��<m��1�¯,�ՋOt=�sWUq{�M�Q&v�
�Po��qA�0�Y��#W�	�Z~>�.���'�H�1r0vH�(�*�\�d���_�vq����:�}�}�ݙ��~���Q5�v}*)�A�d{!�|���Iy�@�|7�12,�]�b�a���^'y�ls�6ծ.�#�1C�b}�5�:�ܻH۩�� �z}V���I0�Nh�ɝ;���=����g���/V��V�#WMwE-]���(71��9:�2��{��/��������><G�lBkpw�]y�^C�S�p��,�2���ˍ���ՇG�}�����o�鲒�m���I�5>p+k�B��k�����3>)��C����ף�J���+|��^JEٿ��%y\3K��^���^r�4z	��Pš����r�gO�!_|����璹{aX1��{1���?	����-�[��5�l���Wy�{ h��)��)��Fc�3<�X�1oΔC�D��X���=�>��4�GE\��.��vU����1-]N:"૝؂���L����n
�2)N�$�1��LO,;�F���>,D'�.6v!�7Aթ�$��+���Q"'��3�=)"�6޿sE3���F�螏CeHD�T	\�P5*��ʻ�{���e?h�K�.�/�c����f��C6aE7%Ë���.�Rc �0~P�#����(O��~xИ	���n2V�^��\�\����5 ͢y:@D���"��in$a���h��C��(�͗[|�� �m�.)�oOnm�Lu����$��t�'Ůr�m�[@@]nq�h�b�VEk�H���%]���ۘ@l4�X��-�Ϥ7����KX�]�ou�ҥ���
��fg:�BA� �45��[Tr��y�{�f��+��X����°�����$-\�2���[b�%�Tt���$���W8�s*+�%\y��⭌f��G����rY��cʳY�3�
� 52��ν�.�Z��<$TM����T{��e�m���A+�Jsr�%���3*Y���ep��9�Xu���[��39��pj�WV�t�I�H�u������a�8�5����	yvi�0*�����O&#���{����ɕ��0�A��	��fT�=��-��!�3F�q���@�fA;.�'h�:�f��WƔt�òB%��֤��GBъ�r���� ���j�#��{��7�dar�^#�t���H^��"����:�vY�M.�\�/�m��KOl	��7�Xo�>�_8vD�j�	�7Ռfܒ����s� a/���V�Y��}���tSm�ʢ�D^kR��Ur8�5�2X^ǚߢ�:m�h�YBrX���%J�m;���������.�v�<k�j��R��L��'Rܨ���s��F��K��.�)�94._�@��&5����PХ�7�;h�h�r;�<K}�4�K�ךη�t�˩��w��*�H�(�uմ�uL7A*��m�씑���u��N����W��Ѭ��x��29ofK�j��)��:�"C���e��N]Ğreي��qJ�������uf�몮��U,M	�99m����<R��9��p�Zz�"L�\��}5�[����2��В�1\1����uv�p���u�I�7�u�M+\oBjLb�Ph��s�%��W��P�'-`2��qjp3�un�ډ���	W�"��[�q�)^0c:�όҞ��v*�/r:��j��6p�j�SQ�/�J�E3s_K�+L��P���¦6]���������h�'�N�oPy�x�	�=�mH� �z�j��@�t4u)slr�#���Z�F�w$W#����۪�*�f�w�����ﻫ�����(��j���ݽ��jD�Fo.ܺa���٥��S�����TA){�!f2��w�ؼ�����&��D@�
�/;˯v�+��F(N�I����	B2���ܺ��ѽ�/N�����wlĤ��r��R�����rXs� ��h{��4�P�&G]̈]ܗN���&���:A{���"�>/zs�r�]:�'���t�N=�僽�ynl��ȓfH���&��;t�.(�ܡ�<�HDd�W�v7����;�dQ��z|A�e��lX�*�&'	���:`��-B)���S�����`���L�n[����y�6;K�錂��O�8.�8��J=�2�Ä3��p�O{���߄�f�;�/ɣ�cK
�妍�=�Ä\EC&v���$�Vf�o��Q5/� �Uf��L@����*���ڹF�x�v>\/������������ަh��Ig��Y�+b.3�5_��-O�}���B���nu�>�Ȯ��u��ct��L}��3�ކR��8%�B��2!g¨/E �h�������鸎�y걵%X�B@�*Ԏ���p�K�7o�`����Q~��;7|����%�L>����F!�>�3�r���l5���<}c��&��2V���	�T�;��謗:�Ί?�1��.��mt��/~�Ύ{P���̓s���-I+v�\ҤM�a��p�|��2WD��FH�y��·׼$�!�
>��z}���[�W�����8jt���b�s"4(�Ȝ����D��خm&�r�om�n�7�tߤ#^����J33�g�����ڧDT9nx�â3b��e`i�0j���h��T��x`I]�5 wlWy����+����2�����י������K�
c���H���A��2�r+�ǳ«�e��Ug����v��/�=諆z��"b�GJ0�B�Մj��Q]5=%]U��g��}�#��\ K���*�����踄uX�D�nx�fY|&���2s�+�H��$��'hĝ7{$������f�^��Q��ٓ�7$���l[Mg��Z���RJ}.c�ҏR.����F��3�>�S�:�{�Z3���kܾ�Q��:_�we�����('��"�͚͖bi|ڽ��9�������g�*Ӊ:���4{�Z��*��4�g�;V�����t�lnzz�������2:i@�yL�(�h�[��(�[1���қ����j7�ݾB=+h;�F�)'`Ձ���-mb�8vzY��Ï��ߵ��7���Ό�Q��Q�C���Aw^d�&:�ؔ�r_����}�O���&�$�y��'%<6�e�5�-��w�z{ʮ��&Ō�tA�62�ta���2�&�rAGt�〾+�&�q"q��,���
��c͓���;��%��E����o:sk.�M�qu��g�ǖr�,ЭH�S%�oG��~�㕹	�	Va̋���L��|>��7�V�|�DU�e��2�+�s���@a\��/n��#9kZw4Idſ(}�ƒ�~�s3*ks�	ȫ���MO5�6k��m��'!pl��B{�r%O���9������qt76������d
��Ɵ)����B���:���o��+���՝1[!�7y#��C���p��(�{%X�J()��D+>�~�{�W����ُ"g'���?Zʂ�R�|Q�����f�V�osu�=D��9/���x�a�ڒ9a�+�uF{&z<�h����T��/�u���ߤ��FW:s�]d���A"���C�C!K��G�Fh�{���0�y9P9t�S��c�n��r�	S��\��"��q���.���|�cw5W;z`�.�j {J���-�2e��x ��T6i�}@x;���?���]�� ��������sul��_92������;/u�tf���E��C�ǲI6Iu�{�FnH�n�!B*��ED+8�-۾v;p���+����L8�p����.����s*�9H�	�#M].\���a�.!�]QF�q&Gk���S��k�?J��H~��!�L�an##�>�!y�(7��8���y喤���������#�zz�Dl�lH3�ּ�Z�7���{@�p��O���jJ}϶g�2-�������/N��'"��#�=^f?N��q\�^�я������r�)�S���ɩ�.��k<x8�~'�r~���.��i̞�FN�i{��"Յ?^��~I�i`�9Ǐqo�ߤY�֞_��=�.?+����7�&[#�t"���}+c����=�Q�τV�&��sz�)'�$X2�`�jo��5��9�7�1|�k���ʽ��:ܬ���˚����!�-3pK��7�Td�i|{)��)c:Y�.�(}���{ҧ���~�v�:t+�9;s�lI-ŏL��ZF���q�ּrS�%�|:�~��h~�:�?�V���D���@M�Rr��B�v(���ge���Ĩ����eXf蓳��*E4���]����(��;iiT�Ѣ5�!=��$�8��Ī�>�����{ c�T��=iL���C�c�'����@�N�|f��1�w���~�bծ����t��.TEt+��}a�RI9�B_Cɐ�]D���I�ާ�����[��ʳq�b:tݘ#d�Qٮ�G}�l��&Cu�$�,�����`��^�o:�u�1���O	��C�G=&72��*`7�*ƻ���1aEϜ׾޼���̯��QP���[���"s�P����c"�31p�<��X�ms얊eȑ�fjF��GʺW��ۧa�Q�vT_{�/cr���^���Xb�J�uA����A[1��)閼}7^�=ɋ��'�=��Q+�>�� ۟�"%m}?{�*�"BX�
���K����ߖ~�L�q1��Q'>�L��v}�ȥD�j�b�NdB�ٟ85��{}�ח�j�%C�O�\�ld#������Ol�V��ѝ��ϧ2L-��T�
����Uח�j�PKeŦ�I�x�)t�ks{s���A�b�v���6_g^\��G;?e��܉�N�W<RXXM#�X�����o��K_^=Bی�c���&�]_�k�ն��誢\�P�Z|`��;�D~^gƼh�)�O��fi�%B�ܼ����Õ�%����b+&s��-����zÔ$V���A�y��O�Ϣ�;� KGn��=���Kބ�[��Rx�O��O�,���	�nV�kv�>�gz4�"������Q�QB�C�e���BP����b��������������wR��dJp�Z.�#IR���'O{�;[?G���ޥ$?�2��m�_�����㍈�F���HEӣ@�
�b�beoWk�Gޓq�B�H�CPbĎ��3-�L`����'��gٲNl.���1�cݷԺ'A��_�����
�#�+���)����>�1��&�6�?R�9?r�Oy|�d�U��+b������eLVG2�"Q��U�������=�2�?�
?����G㜡foO�r�Q���:�Is�Yg#��T��X�&���Wb���R�����6�	YAt����͙��b�ϐ<u���HD�E��ʶ���5,���tLZ����*�d��\�=�4*:}��� �_k��f�dG�a�SĿV�f�u�6�9ɻ�29����`�5_�Lur�3����r���s޶$س髊(�?�Y*&�k�w7�3�0d{e��(����<����d8��(mef̟c�qX�}_o!pi9̋Q�k����n���O��=��$TX[�T/6���ؼv\�W�{6�������B@��h��ׂ�ous��vWCq�C���It���U��a^L�o��(�D��~B�`�a��U΋������cF�#[�o�����i���j1��Ц����)mXu]����zk��|X�6k;����:�j�[�TTl��2.���!K�����β	m?�.��3�6t�7�����:�t�Q���X����7yұo��\�J��m\��2hЗ�yt���P�����0کҍJ��u���<�l���{��2Y;�;���KqU��[��}��#��~���U<s��\z��^W���;���{	R0�����2��[��wA�n��[���"�]��C��$�'s,�Hk��tQ����k�3"ĕ��>o���hz)`�MښN�Ǩ-Y�U��o����謹A��{߳<U�g��c�Pl�bs�+�^0ķ�}�U&;�Rs��~^ޤ���q��N�t$W:s��/����j�I�����W��g�3;/ϩx�0-��@j9�0���Ը��=/�l�
�e�hxK���Q�mo�x�K�tx����,{�[��q������ɉf����z�-��1�:�y�:z�G.�i�Cl�^*T�؈Q�D%x���/2�<���[��zpm�kM���w��N##����;��pslj���^JǙ��=5=(�&X[P|N9��uF�C':|P;�O�������ZF��?�lr������ez-��J>Q;엷#�
��L�{^t+<���{ysۏ.������o���zM=i��VG>q�^�\��l�]�����=���yC�%l3'r4��Fw$_)����U�{S�>o�1`��o��^�C=�f��X�Խ:'-op����ʧl�9�狵��q����;-W1��M͎�51���֍��t��Rv^.��$��8i�H�r��A坏���"|���|K�������z!��hq������&��xoW?5��� �jB���5�RUc�f���%���dS�dR�Qc k�(��Ӈ6�2E�z��p�u��k�;w��19��b�>�\ѸJ����r7�dn{�p���5J����l�ӡ��T��I)G}���:"�����TKO�J���#���z�;�q���i-Zw�k��ޓ��fZ�@�+ʨJ�:oҽ2V��[�nFT=8UL�9."�B'j��ߜ�wD.��P�ƣg����uy�{����&�C�f���񏾿�>�:���Z�
%��W7�����7���*& Up��_�~Edx١�dN)��<���8��Nq��o�{I�M?:&��<�>�e|�А:DM]x�'�4���8v�x�����v�F>R���̩�f�������r��	�]6�8�^�O��ZO�=gg��Q��M�����{v���Z���/��f�=B��q%��u����24�����q����*g�1�Ļ��*�d{i_6���2n�h��)�.��ω5��=� ���4u���ѽ�s
$#K�2�;f��1g��3�VĘ���O�Z� ڹ��m�V��f\�D�t§ �3��D���)�6�E۳�֥��Q�ݺG��mo���~y���^��|�h?V�$�}�~���S����8Gu�'p�՗���h߯������^PSw�X�w�lg㛱���R�᲻Ƭg?'���xuQk��
�)�0��_+1F�3�#W�t�}��[�ឫR��5�J�;��,v���'5�>�&}^pgk`�7:��>Ȓ�J�����K�������#:,��OVr�O���d'�P�	�܂����<Y���|T9�Nz�=�����6����dJނ
[)�<���!���U���ʩ9�oJT=5-3����λ'J�ҟ�uE�R�:q)��9\U��h.�;	���R(�g;�~^>�U�Nz������D0�־+�l��8��?���Z������N��	��o��eD@T�L��������)�����+'Ԇ"���@M�g)�B�xQ3���;�{*�Wd
*�$����Z�m&�o���o+��v���5�Zo��������V�}(��>��j�ֵm�[[m}��j�ڭUsU[j�m�R1I�@=��X�I�M�Y$I�C�p�!T ��
�DF��i	�'tq��k������Gc�7��%!���@�"A�� ��d�  �� d�` DHH�42�1$�	�d���$�&"�"D�CH�%0�BA$D`�!&$�$3������L�C#!"b"i��&d��DffR������z*CC�8�![Hl��C����hP2�4g�3	%.l�8\oIV(PMt�}�6���&!��i����$lY+*f��L��L�i6&h���m�,ٚ�3K2KD����*f$I+6m2l�M0F�&&�)�JI��i�M)��4Ŧ�L͚l�iF��3L��Q�3"2R ��e1�������}�ֵ[k�(5�Zn�o$�~�$;DO��E�=HBJ����.��S�\@}l���E��#[3�4�@u�����h�'g������G�?JQ�@,�d�u�r����»�d�E0>Җ�
O�Z��*]A���s=Pq� ��m{�u��H���?�\������!+�&����~}��j��mm_3m�?�]��yZ��_�Z�m�sV�U"-��В��v�!	�F�A�᨜OVv��� ��� UDɁqDBOS�1�C�"��E�Q�c$8��x%�hA}�(�7�k�B� ����6�_#ބ����"�v�?���ІQDKsYM%�	�=�n� ?؝���B�Y=���&�J2�r����=��Xx#d~!��7kMQ�/'���=��y�D@T�Y@GI�O�����KY�&�A�,��XĆe� ���(�"��> �Lط��D\��2�Q=0ȲH!�,���>4@. a��
4#���d؃ �(A��r@�d0)�t���W١���6o�s��,��{�V�կʕ���7�'�0���\��W"��@�%�DL�h�'3�AN*t��
�W�9�T�{�r�I�>:��vp5��|]��
���#�ґ��P@IBx��e��y�O���o��:�I_��S��x\o��H�P! ����k���uV�B�-Tj֍��Z��j��[ll�U�mEV�mjƱZ�
��k�V�mX�Ѫ���V��բ��cmUkQ[lZō[TV����I��Z��mj-V6��j���Z�j5��V#VѪ�ckV,m��XִV����mQ�[m�lmU��X����k�Q�Z�Ŷ�-�U�ōm���ZM��k����[TUjJ��TX�V�m��cZض�F�[U��!@(�[����G�A�s{á�H����Q��
�����p���]R$�p� jTJ�d��`���x�26@K~h�@y~b<��q�	��U"����C�����ޱ:���"�ڐ���@��s�:�a3 ��$�s�i�Н0�Ɏ���	UIX�S��7°� *~�@��G�
 2 �c�E���863���QS���w�%®Mӯ���M��J���O
/})`�X�`S� �D�s٪&��.�p� ^� 