BZh91AY&SY���t���`pg���gߠ����    bB��             ���Ճkb�l��X�h��B�Z�������"ՔU4��i�I�km6ll���٭���ȟɲҵF��Sm�l[��fԫZhs�.�[+X(�څ�ŰV�U���Rf,
�l�5�j��m�aU�mj�,&S*V��$�(����[L5�V�Q��   $ε���Fpn�m(Ͷe��s�C���Mp,�Z�Mj�e\�J�����4%����TM��3���Em�Ժ�,ղћj�k+4��;�e�֦�n�Q%J �����ƛ��]�jۮ���:��]9��N�iP�ŵcGq�.6���wU�Uی��f�u�M������G+�v��5��ͭd�`��1�WE�-[i\>UB����E_{:�N���@�ЛL^-�EHz�%�J�wy��B�wk�@��+'��������A^���<JUvj�\�T���E�c�2h"R�V(�q}UJ��78o�)U�}eL�;OA�
�js�kҴ���ry�]���(=��v�u@J��}�C�zd)5]�(�*��x�֔�V�N�^w�+m{jAS:��P �����E���,�-�
�3[瘟U
7{{��@������Y��]�JR�����AF�k�JJ�Wg'B���lpf�j���ѪR��jUM�+�^�$(�Q��RԵ�Zٳb��i�m�e���U*���]>t4>����J��v��T[3N�=��P)S��y���h4Z�\R�5(#���J��T��R�:j���T��U=��x*Q�u����Ҷi�wM�֙I|�BJ�^�|*�X��r�P'��Q{4Jj��<�B��=޼��P��oQ��RGv�ׂ����tQT)�]���C z�H��j��+kkX�Lx8��UR��y| 
9�m��ΘT7].  �9� �x� �.\p�]wi� 4�=� ��Pz(G��l�g���`ml�4�yUT*���@t;��t -�7�� 7��  [�qE%HPt����� ]Ά��7UAQ���,�c#X[-E5�M���B��M�o_
 z�  �F5�@&�P �{ç@��p
�0�4�� ;:�*�ݎ tq�f�k*^�����l\� ���(�� m̗ P��F:��� ��  nSӀ ]�p ׽��uێ�u��   h>   @ L�)*��P  ѠA� 5=2RR�#M2bhF�4daOCIR�F ��` !�2d�U?��SF�      OT�F�TC� � �Q"'��AL�jf��!�ɡ�ё���`��?o�y�`?`�+��������y��s��q����s�����I"I�{��I<$�����$����dI$�'������[�C~��g�~����?�����{�u��[[m��_���<�U[m�ZV߹m�[[o�����"��X���"YRO�(����$�I8Y���D�I8X���8T0�8X�$�d�I8R*#�d��$�Q8Q8XN$�I(�N�RN��8Q8Y
���ȘY��8T����
'"p�NR�'
��¤8TN$�a8Y8P��8X��
C��8Y��8T����R�*C��Hp��Q8XN���8X�
C,�p�p��*'"p�'��'p�G"p�'"p�zQ�Ĝ*I�Ĝ(�,I��,I��p��Hp�8T���d���8RN�H�`p�'
��Ȝ*G
I¶XN
C��p�����DÆ$�*'
I�Ĝ)'
I�Gp��,I�ě(�dI��8Q8X�¤p��,��p�'
�¤�,'
'"|(�,�¤8Q�Ĝ*I��p�p��,��D�dN�$�I8Q�Rp�p��dM�Hp�
�$�d������Paa8Q8X��H�D�I8TNA¢8RN$�D�I���Ĝ,I��'�I��p��*'"p��dzY"p�&�	��p�'
�¤�,���=*,��Ț(�*'
�p�'��,I"p�XN�$�bN	�Ĝ,��8XND�d�
H�dI¤�,�*G
�p�l��,���8Y��8XN|,���L)'8RN��8RN#�p��8X���#��8Y#��8RN�Ȝ(�,�**'$p�'
�¤��$�R8Y#��ND�S��'"8Qʉ��axX��$�dG
C���I>��8T�)��'�b,���RN�������8XI¤�*I¢p�'p�J���`8TC�D�*G��8Y	��N#e��p�p�p�)'$p�()g¢p�*'
'"p�p���dND�dN,'�A�Ғp��,�¢p�'$�,C���,���p��,'
'���D�dM���8T�I8RN$p���$�Q8T����D�H�`�dG
�p�,8XRȜ*'¤�(�(�*G
')RNA��8Y�Dp��1´Y),�Np�dp�8S����
8Y8X�bxW
Y��+�xp�+ep��\,�N�_0���+��)¸Y����d�\,p�8Y¸^�p���,�g8W
�gJ�N8W8Y¸W8Y°�����8S��,�\+���,�Z+��+��+�p���¸W
�g
�g
�p�¸S�p�
�N�F8W8W8W�p��p�
�|)���͖p�¸Y�f8Y�𳅞p����|+�p��l�p�
�\+�z^p�p�(�xT�g
�\+ҸY¸S�̜,�,�*p����a��p�^��p�
p��\+��,��'
p�
�g��,�\+E�g
p���K8Y¸X�vS��)¸W��,�g
�[/8Y����8S���x^p��g
�c�p���p��R�)�,�gK:WJ�*t���,p�p�§��>#�dO�$�RO�A�I¤�,���M��&��|��h�<>�������F�PiP�ŔA�R��z/\��l/Tp�n^�ҝ��P��:V�ս�j܎���Y����*��Th<ٍ���nJ4�W+fE�ȭ7�4U		���x2MJcQ�X�A�AD0����!�\����&t֭v���FT��ܩ�AXn�6��扔|\��J�^���y�L$�"�妳-�q�m뭩�L�L�R�RW�KzHܙ�ս�(<�ӆ���[?+�1���VYT'Fc�IW��#�Q^��'�ª�=x��d(�4ګX���Kf�z�h;F�n)��:������U���!����{BЦdPR��F�4��.e�xr�0��XU��[iiSI��m�p��Ѽ���5�mdL�VS��`�x�Qͥuy��l]8��RI�ڣb�ElUi�!Ta�8�����<�.kUl�ڬ24��H�ި`�%��Ye�t��ܺwY�jd��f�hIovS��AIQh9L�uQ[��Ve֫�b�W�z]�h�����8�E�L*T�U�G)
�t۹m�jI�ʭT&�U�D�c5�Ӑ�۲H�;�n�]��eݧ������b�*�����<*<3+heoe\7�y����\���qUJR��eX�[P'�����l�+l�g5+�1�4�=R���m�1�Py�A�MRn���km���c�Ș����*y��w�N+V�hwp�u��u�,�[u&�]�K���j���1�����ĺ�q�N�K�p��$�������Yu����kƤ1\ep��M#��kdZ�#n<��y=KZ&$�@�6�rkL�b��P��q��FKbK�u�س��E��j��\�j����nhvC	X�ε�EBc �A�W�d�)�fir��-�
^�?�:0�yy��*y���nU�p�,��qlc!�bQ9Y�=�v�4��±��s���v���2��:��T�B)hˑ�6#�GW�����&@�KA�5�/0���Q�r�˥vrιU�����%��p�&�=ŕ.*.�^�e�����!�"���#����Ԋ�ܶ(F#"/b��b�'5��G*+6�ѵ[�˩��YoB�%����Ut��p�12�ه��o���bW�i�.�)N�emc�����X���E׸��Qق�n���m�ъ�j�[4hj2�B4]f��b	�n���oO2�9Q��[�&����J������໽˺�Ќ�2��f�:�7D�+6֬�V6��T�̥*�Asl�/2E?�6��m*�e�Jű�7vӢ�Jf�,Q�Ĳw[���ֈ#&��U�Q���9G5��#��͏D���ؤ.isoukʠ[��)&+�Vڎf[Y7S.�����)S��t���)����F�b��a�d�7-�N�di��1d1��X�Q����v��bF�*�Da�E��_���N�X�)��e����Mķ
˶��	����5X���	��5R�v�h"��I#0��(O�]H����uX�؄�T!�e��Z6WY��1f�l䭽�X�U��Z���,"(�.�Ԅ�����&�*�yf��,�{uP�ڂ��47����٨VcN�L������wUf��
$�F��M�s&Ԋ�����t��ѕ�{.Zb��V �ͤ7+Ҽu������AD�����T^;
<��q��nW�i�MIB*�,�6����a������ŁکF��w�zm�U����n(�)�՞�y(Ev���dʥO5� �W����`�1����{�K�q�~��bېw�U�a�]%��Z�㷡��LQe�@ﶋ�Z	N�ˆ�ʪ�fbYv��@�+A����;�øü�S��Y �R6Փ=z3v=���r���.�T!�妩ޗ�j5��pe]ê��&2:�Kpnlj���Dol�*��-����*4���ڶ�ɛt)v7Y:����� C�B܌�Ac/C�Z��u��G6p5���9�1$	�2d��䪪�8�򤅖P�Z-[n�Bc/)f�#rօKi.�wY�b�u�=�.�5Q9S�v�P�;��P�EX�@�����O6W��7%�{{��X�sv�O]Y����#�T��5ӭ��8V�e�@�UT�"iQl��jEZ�R�e�2h�d�v�L�[4���),����v�	��������6����\�+}bߵL��+v�۞*e]�Z�ư�}h�n�
F����d��������16������w�mF�]M�Qꅱm("r����T��癵hٿ�j�IS"4��Ip�U��pfiww<[ʘi��r��I�x]ǖ�U�;xl�%�vr)u�NK�X�KT����r���2�zю��'Z�n�]��Ѫ8�����Oq<�U��՟�nХHi�t�ۏl��l��ɽ��M�wRg�
j�ǧ^�I��VjQ8-[^Ue�ʅmI6V[��I���۫����*a�wf8S�*hڔ�n�ۻ�lTI���0���.YY�U�.�7�b�p�i�C/+shXo����0���V��A��V�z�ʊ�a��.��u/�M:Ȗ+�g�@�I,3�5ټOT���3�U��-N�l[r�ܛ�C���<8��]�s��)PB��U%�Bޢ�����"�E��
6	��ӡ�[jma�NG�%m͂�5Se��q:�IV�]�Ī�����P�b��m���D}��ޤ���eT�j��x�!b��3=7f�B�cy�Lڑ�܈l8�(U��w�f�7}�fH7&M����H���*�7jνq=ۧQAwvU���Q6��vTی���^��*�M�Tv����Mn�(2�]T��ۀڍ]��jp�J�.�
2�U��y��.��ǳ.�U�;o4I���p�\/glT�֫�GJɑލ��$��Gim��Bt7K�nERGk ����*�9��q�sl�{��]*�1���e�Sr�����\=���A���˹�J�_�H#����)�gfGh^�ZU���`��2�+�XJ���YG-�m�&�%�n�����h���z��EM���ܗO#.�W�{X�h�ۥ���҈f9�B��q=<�EFE�	Gt^#�@]4�bUR��9�!���BtPg}Yah�y�t��َkj�ߕ�0G-57tQ�kE���[du)c�⧍L�V��0?\Ė:F����R��L���VK[,��f������К�˽���/|�fY��T�	)��8���
�dA�9V��=WN��:K�9�U��3(�rՃ�3�P�ٮڒ��ܫE��!jm�kN��iY���9UP����l�!��¨��Hֽ[e�RZ�x���m\4��N�0�PN �kD��9j�g ݪ�����öK,Aț�T�ݧ{�,�����8�+f٣r�¼U����HXz�.�m����z2"C��4H��VX0H�Չ�yx+K�Ya�2�wTm�@d�r�Q� F����Z�Kf�匡��8�C����é@È�#4�+����i3�ׂ��触裡Ӓ^�]x3��k��rY,��D95Ua���Ř����Ss0u��ܤ�t�w�B�J����2�͋��6��V�8q�;�r�<�0�5I��i;1�QAP����W���H㢓T�b���{�77!K0���Qԑ����j��t���m�s�31iqb;��LM#%d&��PQ�ZkͶ��˵2�I��%�$M���i<h
�5Y��sd���&:�L��jQ8�RsE7ln�s6#qY��lK0X��1��B��4��9c��<3)�66���X�4!דu�T����<���m�OKIU$���m��^ma��Ea��[�֚��ٹH�FĒ���v�`�{�b��TR��M�AV=g$z�8��/f�P�T�޽n�9#�r��2Hў1�Z�UP�N'����;�Q�[���:GpゃM��L�����+��:*Y�cT�ì�J�>[�v��Uy����
��&Q�Fa��em%X񻅂1�+%��m@�^*e�U�-݊�i�ަ%��v�#Y��0����nf��M֙Rc�A��`�eѱ���U��Mj�PL(l��Lv�D����%�c.KҢ9@��b��]�R�DQ7�d���1T7bT��j��y�`v2��;���t^�Ͳ�Cx�nQ�ʡL5[Re[eL��ndM��A�Zbc�´�m�6֐s2K���.Hkk	����I�b3�f������SM��ݓM��(��Bv[W��V�dH���ˤX�F<�y�zq�Ò�M�W��!���ێMV�R��(��[Y`�T#�.��8Nʫ���r�+B��wt��k�}e�1�ܪ���V�\�X�:f��*��t�ɱ�n)�v�3n��pK[%�ѽ�sZ�h�Qٮ�^�z�%�G#��z�㦵�ɗ�3iiE�)ڲ�[*�
l�HjcF'I��J��c��+E8�F7fc9�vlb�s%��8��T��a�c�P�TE]Y�L)H��b�ͤ�Ut�(��M\�fPM��5h��-÷�0c�33�nR�7̤����\�bsBfͫ�V)*�>WV,�{��.ԡ��$"N$�l	qR	�Re��2Tg<�NĈBm��1-b�:2�cE�eܕ��"�A�H����.���j'�k�*j^[���U��ၚ��U+Q#0��I��Y�
�������a�nIV^���Rf�����f����fIj�ko��R�Q�h��ꤧ{1�pT�z��57s(e^
����ENnl����%�Z�ޜd�dLc
׮��&$�lxF��h��7A[�]T9a��-^&/U���x��Ra��.��vC��F�`�b��I�X��m�:X
�&E��Ȱ�:qS�����mD�ӎ@�*lY�(\�,+c���WjG���[BnjF�LaXV�[�B;6��)�.��RA��;y
YN)*�Gn�a)�*�Cv��PI%���b��{J��<��j�B�gq�F#�dlw�"w�Q��JcO5)5\���w[F��l`���XY )�<u\�w�-����F�.o��om�H��R�YW3E���;uL:��Ҳ���D���R���S��^ا
\�[+1��<�#�u��$�lچ�*�&hPa&iz���1��8��)仸�ݬ����*�kHLie����_�L��25�b��357*ñy�C�yӮX�"��yx��%Qc��)�Sb��2���r�ˆ���{7]��&K�Uc����h Y�ۺ��n��F����K0��A�aGFb��ub;N���J衵�ng�[d�d��I�4,U%�#ś�5fQ�&OVk8ʒ���-m�TH<�l�lɵv��cV^U�U[�n��,0k1M�(��h��u�d����n��r�iɛbޜ*�%��Y��P�dU�t��Z�c�0�J[���ʸ�5�,�ܠ1�mw�:��a-uQ�hY�u`�Ta�ِ<��wUwz\���u.\�L�,,ڲ�E��56��n����f�嚲�Y�mY��";�Z�1�&[
��B��	������t�4����vWwMF��d�=.LD��ڇF��E��U����l���{w�G�BJ�)��^���l۪��i�%���#$�!�����UF2��:��Zj�f9O7K7�0�v��3-*J�=e��=�um��V�.�#d@�r���-�A��ٻ�!P|��>A��P���7pX�����-1�a/jA�2(�ad�:���⃽
��:!!�w�{mP*�I	P��ރ E�KH,�a�X.�J��	0(�0opN�D�-区���CL���^�,Y�$Z*At�D@���W^o���
�MV�f���6�u�T����m�
 m��'��EUi	�I_|3����s����b��9�,A����~��a6
�W�XYD�X�̄PQ���>2�=b�	4/0D�x��F*�A�z5p������B��!G�,8^����}�oAtGH5��:]��Ub��~�b�6���21�|�|�u����d�_��l ���W�gW�y`KA�(x�D^`��ߘ��.z]z�AY0g��Q|��ؔ�;��%�,��	A��:�:@��<@�4K�na��B��
BՈȒ��@���04��
�^`x�4B�_�B�З`�M~o�	�
���>�c�������2����+��o{��?��@��a6�*!Z�6@�P�F�
�������;�����P�ߎ@�<H���[B����B�0�,e!+>�("���F���j��`�A�3H��˃Z%�9�+���w~�r�����7�tXUA�Z3�SF_�P�*�aH��]�AsHƅ��Z4`��2#���	�><��=�,|)o�@�~pL��
�����$������V�hu��C��p$�D4AG�6�5�����cHbb��1�|6`�c��c
!Ɋ0u�Eq�g�:A�Cj
�	������b���a�
A6
8д���b
|+��x1x�סѕ���K��:�W�4P'ʻ���9����f�:Pkݸȫ�J�2�m`���@���$#����lpT���k��;|:X�ƃ���/k![�L�c"�	lB5`R����� ��/ vD��X�{�C ��1�_í���C�2AY3�5�f��:���#�2	v���s�僭��7�up�"���;|m��SC�oA����#:�戬r�:
Dj��.�b"�p]�z���N!��:�2�rb"*׋�T�,N�g
�"@��Ƚg�Į	�@�:=d���y�2���ë=Ha>���T/ �������A�+pS�l�y�L&�N	i�H�77����������ߨ�?C����-�U��xz��<Xۊ�q="/�^=�r�.�d����9��i�)m���Zt9n��jS2�E��ַ�Y=fg,8�(np����N��iv1��4��81�y��gVh��o��[�]�RU�A�}���A͕���]��#n�f�,�9	P�~����[LM��W_m[\t0v�!HA�A�旂�����"��JG���w֔v�P�Z�6��Z��\;�q���Uuי	��/&�T�<m����Sc�̚�r@⧫ޭI{j�OH��-L/tP{1��Ԧɺ�e�z�����ug���N���Z��u�ظ�sW;���w9�d+8�"���ㅝƦ0�V����*]��nL���:�hJJ��5'�^���f-�^�#αJnwQ�H�(�Qt�5ڭ�L�5�S_W\�]��_���k2���3���x�lյ���&�m�΃n�b��C����6��zn����y��.�kv��8�#��-��k�h���;^����Ł=Y�ikW��+��s��S�f,4m�W�Oi�+��Ð8t:IY��Ruz���hw��r�΢�\(�tg�V[�5����Q�Y/}ݧn⼛�l_-�$]I9�B;Zi��Zv"M��p���ު��ܥ��Ŵ�ᓜ�C4p�6���)�d6DĪ�D��ޝ��=�Uδ�l�Mvd�T�`�7�ԍN�0���.-}�p�����1$"��#�S�ƴ�o4�5�R�5M\ɩcƖ��N�pk�w���\���F3��⥳�\��Mm�i��Z�4掦���uZ���hH�3k�7&'�Uʳv��k*�U�)ҽZ��z�c�mL�-an77Ō��wmJ���T����p9ҜOs�WeN��#�EtBN|&�*�_.��NAL�۵�&�`bԱ�p�U���N��Z7�bڋc�z��hfSr"��tq�*�Vy��k���m}<�)���r��Wf�z�����<d�n��~��GWH.�UǇqhoR��|ݞ��cZ��돏,���-�%DgMFe(��);�ұ}�������H�3i�Y����)�>�J�iG�1�����Z���ͮ�0v����̮T��Q��L�}8��ԧ�N'y�)�C�c"��9��F+j<4�_B���f��k��/���z��]7�2舞���ܸ�[��%Վ���-�[b���i���Ų��<m�9�Z�d����Y��w2_��x���:��ܗ�O;��v�i=pN�fu���&e�n�qrIX��K�0L/\���?-����lo0I
��Ϋ�T*WXq���/vV�\h}/��唾V6_XGr��d.Z�6�Z\���&ܘn��Qc��B�0`�U0�&�5�pgpb��:����P��R�B��rd�7fS��D�ohk�ۈ��WՏop���D�ne�of��[ceb�>�W4�ӽ��Ȱ4�[JSO,�޾�6��ʠ�[+��-�ΩZ�U(�dm��)UC���*�R���XӼd�S�9�G)�س�B!��y��@ԥ��*�Ź��>��"�zqi.㨸D$��q^(u�2{�V���W��6�>�1ކ��$|h��Z"�۽۠�d�h쥭
��`��h�xV��*�����\�U6�0��컕��H���1�ҥ������2����5X�FV��o4�����MV�c��ج���]CI�sB�K�*�*;�H3Q�-��ՙ<�Tj��'��ݳC5wX4/����5��J��\�Y�D�]�G��fMc��av�3V�gWXL����N�N�i�ݒX�J�t���oXAZ�#�9���⬪����*�/�Lz���f���r�<�ɏ8�!1)n���n��������tr�cOu[�:��LT�ʟ]]Y�F��V�Uޮ]E���>��3`�����9ɕ����lHz��މ��u��n�gQ�-L�{�Jj��yήUb����;d>n�/I)+��&櫃UR�%K��N�cb��UY��:��zS7���o�J�k�p���ss/:А��Z9�&���~��x��D��t��ɷT��M�Z�b���9�WB���9�V�NV��%[:�[p;Wˤ��$�	�0#�v��O���@�1����&�>�����bqK��)t���=��[��أV�B��;xucX/:о���uko��u��K|�Zk�c��<�eC�cID-*��d������M�W\��;IU��pH�5`0���}��3�M��l9goj��'%�N���4o8Bb�9{��m�sY��d=Rr_��˫9��a��ӥ;jt�y-s;��ӹ<u�ɽ��7.��Ynv뱙еd&�&G/7*�D�Q�q����pc�Ϋ�捪i�Z\��D���i���epuD�c���ؙ�\\�<Es�|��U�1���5�iKd��f�,Û&�ݻ/Q�f�6��x[=x]׵&�.���l���Vf��|�6ɲѓ;����A�M�y�<_L�b8�A�J�ᙅ��9���N��X�Vv���\�t��4T־�U��Ze0��ȇX�P@�m�[��.��b�e�G/i�ҹ��uZ�q�}�azI|��;]�=2I�����y�v�)4%��N��A�+��a���Q�;-�y�-HU�ʍ]�a��?�vz��W�Q�ˤovM���vؗ�m1�GEv�����J��<�d�4p]��j��]N�	�V��Ә�!���Q�e�|��غ\�̭u[��}�v�[|�N�j7\�)��x5�ƭU�*�;��E��A�˿�՗P:�%�	��O�n��Y{ڤ˪��-��b��E�r�-n��b��&�c8�]�/:�z6��lw��6�}�^�[����8���ԮЙ(ۗy˘���˖�&��n�z���V� ����iͪ�nP]̰�5Wi�j�+�R��z)Q�CM�
9j�>���]�fC��-�[%�:K��L�zV�d���w�R�L7���
̏i�WE�.Wc�����jW����ګ�I���	���7E��\��ҁ�7��j@��6��==N#}:���[���Va���)�A\�r�B&�{p��0���L>�bv�]��f��0�:or�3���ġ��3c�$�B�͡N�ɛڝk��u�U����Ge�Dv�s2�Yʴ��kiW�Z�GU!j��kJ�D�=+u%���-$��V��
���Te��e���i��i��:Kd�c�u[d�#y�f>�
��m}'^녚�RL3�s���A+kx�7y�xBjn�n�e5����u;�Ƣw導�1�d�t��>v�^t	HU[y)	v�2�VS�܎8��TN=֯b��Q4i���1�q����4��{F_*%v#Sn\�й#������׎w��P��#c�.��`��g��*�dQ*���0�=擻��3A�K/M���=U����c�BQ&�d���κ��]ҥ�o���i�(��ꇉ�!]��#�tE�#MmjYcgm�kB��o����yD�o��it�G+�ivd��}ZZ�nL�-�qк���S����0�#����\�֛D�+o�0Xם��Ƿ�Τ�S�wY�� �`C����Ve�y�4���E�-�.W/\x��|n[�yΰR�&����N�����x��T�����T�.�z��Ѽ�
2;��
�s�9�py7��Vӌ��6�I�Q��t��oP��\s��Ws��v\�cR��.�c���W��iP�j�u��-W�WD&�ݧJ{5��.��]`/��:�Yms�+�����z�NV���|w��V��k�R���t8q��_P���Rn��Q���竄�����Vv����:�X�u�������m]r���\��A�;|8��p�[sJ!Z�.
z�����R��1��x�=�5\v�
S�v����rU���UL3Vș+���U�2n�˞^[�h,����8�h��u� Gj�r�6ۨ��*��Ϋn<�jUT�V�!E?$�w]X��OE�d=w�]���ݗD�M%z޼�[::�in�
^^��ص��Έő��[3s*|�L���8��Tb;AU<�u�A�vvb/�+�8��s��d����:䩻uw���̽ƅ: ����N���U|k���/n��T;0��E{F�<�Y��S
������"=jY:]�]�>}��W��3jp탫a�:��[���`�0�M����sP��"�Xq��b�%X�N �ћ�On�d����`�nf�:9�����V3YRբ�1�J�3d�#��,c�#�����h��Xݼ��������v�Q�:��J��-�9��X9�h+���D�z�Xr��F��O�z5޴��ҷ)���]9��#�����Ά��oup����n��yd�����U}�Ϭ�@�C��}�b����\6H�[����ҳl�E"�=݊��E%��@�!;�5�ᣖ<G�ޚ,Չ��m�Kd�d�R��c�E�0��O�we��s�M��3uK����.`��藏�x����A�_c�yd��GFn�f]M�+5wcwρ����K�ҋ:�K�cd�QW��h�{Y���������]��.�3��`u�W.�F�s��u���uΗI�v��ĤE'tÒ��:p��Uխ��w;r�p�[#٣�r¸��E�)����o'^�9v�Χ��ᩋI��q����ֹd�T�tŚ��Ժ���x�픭��+r�㇞�ՐcQ�w������t���J3�\�gr��+`�2��J*)��ѱ�;4sYR��7��M����W)�m���vp+�2.b��NI���+�s�gY+>z��e�Ç�C��(�\.�VtewN��Ӽ'f�����1���ܳOGY4WPZ�B����r�-�D�g�_p0.o1y�5��>eb�m�UE�n�.gV�rv��P��n�@�9ꔺ��|T�㎱J���1��yR��V���1k�l؆�ܙ��O5��i�.��U�|��6ݳ,e��а�֋dVuv�}�g%me��Ӑu9u���Җ#���	����Z�	�	2�12�u5:㞜���^�MOv�ʝQ�����{�������������������������mQHڴi�ő\�<�"�#j-[u��rY�m����f��	�b��W�x�L��V��.UR��2ti�!bft]��T�����W�T$�8�x)���]����y�K�q�;vbv��km�ՋaD�_NU�n>ڇyR�m�A^��d5�v��C*�,I����ju�X���ُ'�:|�6�ɓ���7o�fU�end0�Ak��§u�����x��l.#�ײ�c���5��:Y��N,���Pm�=fG6��W~�S���7!�r��ȭ^�]e
uؙM���{�!Uw�Jt�5����z�i�����Q��i�WEN>aP{���Dv����bU��wN̪�o��%.@�oinu�'Y������T����0V�z3���^2�jN���]r��#�6%<}�=�J���ڣ0�<��ZuHLs�`�ڥ����k�R����%�ꮘ�o]N���4F�]ˑ����|t�O�_w#��-���i3-����(\Z�9ڪe�h���-mR;ܑS�^���Kx��}s���Q��o�wܜ�w�U�m��Xzz>�4"�Դe,6��7/��}���{���C�f5�ٛ�l���u�U���b,�}�����bI��{ĳL�є�S���n�wX�'\�;2)l�ܝ�V�00�A0!B F1��Ǎ��яUU�lu���|ci��h�J�lR��1�clOҪ��xǌi��ƛl�ک���Jz��^1�W������x���1���<+M��x�X���Əb��cUa�++h�b��M����m֘�׌0۬m�z�=VՌa���cj�iZi�+EV<x�M4����b�[UV�m�6Ҵ�ƕ��4i�Lcm��+f�4cM�UU���lUi�ƛJ��⴬V��R�Ѷca��mX�i��f�S6�LM4uZM���F<6�h�W�c��M1�O[aJ�M�cM���x٦<J�4V�V+lSJۭ�ٍ�T�m�Sf1�1�+lh�ja�u���x��V�m��ƕ�4�i���i<c�iR���M4���cm6�M=z��į��|cMۭ4�h����I�<i�xǆ޾6���J�m�7U��k�&[m��%L*FAI&�P�"�Dc	�6T��8�a��6��4����p$0����uB"�@�)�4���
��b���Ć Ρ�<�[� ف�!ƿO�
����S0�oL�$$,p��P��H(�T�DJA?��QU�a����`l0�%�O0�(U��L$#�9�4N!�E	L�`��U*�UHY��Tl*aNB�3QL�Ʌ+%��G��f~A��3	!����(�-��2�@�L�D&0�	4\�%�"�p��j1.#)�"@��
���A���1��QUB?�$HD'��9����~�����#��O�?�$��VD��?o����}��Ǘ<�;������;%^������5�dU��cN�钷�tB�O,��˥\b7����9��2�,�U1��]�k����t5���Sn��N�\)�G����E�W>�K�s�B����5,u�B��R����a��[�{�	%��7��[���n)s��u8Aى��Z�#jvS �u�^>���:Ǯ�R�M��ݗmo�)�}o���n���S����wqw��j����N=�Y�]��LJ�@��K�R���J�ܓ�����[�ǒ���Z��$�*2��F��g_J�ߑE��Ri1	1����+F�j�G���3��λ��^U�<s#'9�m�C��
-�|��öӼ��ʺ�G��7}˚�AN��p�[F!qxf�he��C��P�yR<�@�!7vڌݙdF�P�R֝�N��o�s����'nӵ+��%�/�
��3����R��Tm�ʢW����޼�)�9'[V�V���6����%�4v@৴���G�(ln��/3����̎�_��uNJ��\�dhL.�5!/�c8�ϱu��.�E�vpw���K��t�w�T.��=�aj��q��0%( ��� ӇN��ӧN�:t��ӧN�:t�ӧGN�:t�ӧN)ӧN�:xt�ӦΝ:t�ӧ�N�4t�Ӧ��:t��ӧN�a�n��<�ۃf'A91^Mk�,�;�&	(f�J�S��1q��cQ�ьW��OG3���Ә��1S�Z�	��ǽ�ju&���%����p�X�;�if��cy��n�!h�r����)��J�z�/{*v�jf��0�M�w�������6"�n��t�b��&���a�U��v	�4b�^%�]�������V�1�//:R�|�(S8�S<��mi��ʫ��.o��9��Mܬ�!w��:�k�j���]e>9ź�-ͅ��à�9p�i4��j�_a�+��S���ws����o��Jй,cɓ�R۵��;iЮ�fV[�gp[��niJ���n�Ʀ��S��<U��֮�uG�.��&�m��!LNl�/�I�ס˾�)��Fżx�*�;^%wJ�����%LM�
\r��`����i��Tj�����t�ΞԪz�4�ܚ����`}��xXkT����\JP��4��H.p~���\i2�7ڱ%�	P븳%Egj=R��Va���he1}��bdf��n!�cy7s�m�{�Hu�Mˌ�2�:�a�C���M*Րڗ6�	B��E�J(]sÓ�i��9kQmx\}�Kv.�!���Ms�W<�X� �`#V�E ��Ԁ}{����r�P
�;�/~OkY���>:t���Ӧ:t�ӧO�N��ӧN�:t��ӧN�:t�ӧGN�:t��ӧN�:t�ӧN�>:aӧN�6t�ӧO�:a~|�7�I���[�Q��ohR�6�B�P��whG�g�#М��P��8�l�Cɫ�P�9vYނ�(`�7�Y@�%�y�R��%��������\�H�W>�Ms^/�B�v��ں<z�c�r�b���@�n���~ûC;�Y�;h���>;۹������d{y����n�r�[5��b���@vP��k���'t?\B������ �"
d�����,�e����)1`�0)^j)1o�Vh�aQ �X�bD=�o0[yC�.�}�;��+�G��d�걊ǼH�b!�]�$�`xy:	����x���EWT(j�<�J� ]�#���+�K��b���u*���G����6c��G�*��������e4c�v/����wn�.5d
�\� ����n��*����I$�Puv �f`v�%�a�Å�l���B���@����Dsͪ�@+�b�Xz����J�
LU�����c�z�/ƕ�#�����3���=��ଗƻ�:����tͷ� ��(��3��z[�%��c����w���ϝG`�m��)���r%�|���	��P�=����([Q��B�H*S��tJY��)/��3Mt�g��~�Ae��J��{�Yt�݁�eص��Z��K.�$�sf�Q��픣o1���+�D��\���/z[�*�6m	��B9�C�o���$� z�iB����O�Pj���A�e�LRa�� 7KE��Q�Үq/���i޳h�4�)+@3����QN+�*�:�:'��<֧��g��=����G�çN�=:t��GN�:t��ӧL:t�ӧN��)ӧN�:t�ã�N�:t���Ӧ:t�ӧN�8t�N�:t��ӧN�:t���|�5�
�:�]#R_�}ӭ����Qv��M"�#�1��iVk,�3����]��ٮG�b�	����>�uhǩsz�Vvs �v���^�̭ ��@{���Д�� �uD֛f*��^�n��j�R!�UDB�[T�Qǔ�PL�D#�m�*�^y,�ú����z��W<����Ӷܶ3�]�3q.̫��I`�@���1:'�,h^bg�ºL��VT��<��`�W1�gR�0��`&{.�k�V��6�����Wu��x��y`���� {�d���gFt䳿h��^�^��v8�5e��ت��w����O9�i��ž���D�M	Z�g�«3£�a�aX��Q1���Z(��@�ZI�̬��C�`Gzp�¸x=�K���}R95���~�U�F�ܒv�pZ�or�E��Z����3!r�i�1ćέ.x =��f�w�K��T���n�:`�W����:N�'s����f
��tV�c��3L�ʮ�a,�H��6;��ٗ��N6kF�L�f$��;���g��}E���)q��p��)�����8#7��ݎ!�@LUG�k88Rw2��e�0�p�Aл	�3��62�
k��^e��º���3De�w����7ѝ�S�;�|t�-1�����k�=�A���gO��:t��çN�:l�ӧN�:t飧N�:t��Ӧ:t�ӧO�N��ӧN�:t��ӧN�:t�ӧGN�:t��ӧN��p�7�b��G����NDe��)�xU�� ���}h`���-N���Jm*2=�b�),\79������|�6�H�}�I5Go.�NuWf�1.*���ͫDйX�|p�Q�&Bq�#q�2�=�4GP�eM�)��T�uy��i�(fv<V��ih�]W_[�THl5�;#�x�Ǌ��i�|�@#Y,��i��Ѕ�K�a�z�D��6n�]ܵ ���}o�%�;N1U�fk��on�5:A�����v퍶j��Nжj��stp�]��()�������C�M�e47j��c�p�W{������ә�p��r�n���9����!`����Y�ΡȘ���m����U�R��(��*�?.'�iT�_vZ�F��$� ����(Ժ�4(0���\�uwV=����f�Ik����L{>����5��$��g_R��t���,�[˭���d��6@���R�Kn�ʸރr�)��P��{��0�]���u�5�,*�x;(c�Du��N�-O>A��V�rsA9w��%��Ѷ���]�Y9u���I�+��uPg�c�ż��}B4�_¸��kD�����2�2Jq�ۡ�b��U�L��6h��Ӈ��:l�ӧN�<:t��gN�:t�ӧN�<:t��GN�:t��ӧL:t�ӧN���:t�ӧN�::t�ӧN�>8
��8
 �$&�7�����k2���n�Ty���$���}�����F�}ΐ�1�2�8�k�B�[2��xw�^-�R�!޲-·v�\w)�=
	�9�v��ޭ�<G c�u�g!}	c����Γ�ugZ���es-����~ީ���<8*U��;)�u$�]m]�Y�+ȷ)^���㹩7�P�)Q��U�n�3µ[�M�rʺ�Z��#wZ��-�,*�u�T� \������w5c�	��z��zS$b�\h�C�Wۇ�M�kGl&�'d��]Wkw�䶰 ��b�0K�t��e�Yk�T��a�����+��A]P�tzT�qk�{hW'��T`D(�J/U]�h�c/m�R�歉ΩN�#��j-�܇�����[Nl��x����iV���G��b��¯!�_r��.��.����#�T)�LW7u�!n%B�ˌ,8֠�sx��y�/�ata)V�����,�Ԍ�6DL�u��a�&̺�/�t|\�L���a	�+r(�]Օws�T�ybwE�bU�>�b�*ټ�L5{~����^Ȳ>����ʾ�F���^u�g�X�|��+j�av,��c���͍u�G�������4t�ӧN�=:t飧N�:t��ӧM�:t��gN�:t��ӧM:t�ӧ�GN�:t�ӧN�:S�N�:t�Ӏ�� �5�62�>wT����Q�����g)UPV���ܺzl:I�����4=�y�{ιWn��ǻ����.!H�G�CV�.�mp�r'M���T�l���!�����ڊ���ʼ��;Y+.�bO���(-o���r�ݱ-�B^ګ	q� F���c���O9 ���>-�%���஄.n.���X�Vu��S�!���v����8��.�k��ػ��H\A���2�Y!�U�֌��NR��ON�<��3�5ò�p��r'-÷u�`�x��
W�����J>u}�r�G0��R�'�;.�zЬ�q�ͻn�&���~`<��ʻ�5$G*^-ͧ��T���/��/*�N|���ǖ��V��Y�(��"���7�՘m�/�����+ew��#�]G.�s5Uҹ!:���Z'��A�-in�P��XQ�&�B�]�^
C���G���OJ�f�f\+)b'L�*�����6��7�X�aֱ��m��9~��ybD�P}�����̊9�3M�����Ƅ�<�/��HР�\qes���YX�s��{��k6�1L�Eۖ�5�M�=Rt��u݂���˛��.��<���s��` ��iӇJt�ӧN�:|:tçN�:t��ӧM:t��gN�:t��ӧN�:t�ӧ�N�0�ӧN�:|:t�N�:t����ӧL<��;�2�޹D�:��V���a���6�m���9*u�u5��o�ߴc�{vK�S��Y���!
�f^&��Kt>w�k6�;4D�G:faf%�b)�6�։�Ѽ�x!�������эd�@��h���G/)�2�Μ��WC뺹]��uhGz;vt=�,�݀ʫǫr�h�NRa�3n#.��+�2�d7$ܬ�F�.������Y�U+���tL���s�]&{^�%ѭ��^�Ks�������s�7�u]h�q",���/�f�GfQA��O�#��V���e�4�1X�Y�tJ�W,L��*��2us$��`U���̮t}�Ux���J�����
�q�A��=)e^K��/V=�F�C\k���q����J33]�UlyW�l�7;m����;�q��x�"5	y�7s`�Q��ݍ��Ҳ,�*[�J�XS@�5ǖ��LX�neV �]�z6gs�Ջe�r���s�x�������M�����KTV)Wb�-<ē��OuuY�5E13\3^֨s-���a�����vB%Ԙg+'i[�df�Ja
\	N��s�2�"��G���a�tZ�:I���SK��h�;n��5�Yo�B��!�:|:t��ӧN�:t�ӇJt�ӧN�:t�ҝ:t�ӧON�:h�ӧN�<:t��gN�:h�ӧN�=:t��GN�:t��ӡ��8�l�\��Ͱ�.�ꆻ�quaYuU�
"f:k����ػ����PΪ�-j�m�,T�y����BlapKU�,�"�\��\��ʬ*�e\V�w��)��nծNgYH�w�xM۸vG1B��P�r�ڬgonצ(�h�i��׽G�$��T+�帤���q(Z"��b��lXz�X��L�@�n�2��QC����jn�٩c��WC|5�������r�G/ ��5��d�zi�+r�T�{g�m<�駜�6팖����P��f��z?t�
DU�^Ĩ��{!\N�����Oq������ʜXSld���A>�
R�����+S{��	�$`�Z�aH�'b���!��G�nN���Ү�Z�pk�5T�^f���d�-uE�C���i�R�u�P�[Y��.P�@�-K��2t�R/�jRBHrR�{��)�O��eq;#�;/�|_���X��X�cvۂ�:�Mֲ<�W��vr��_k8�L�4�O��VsoecܺBػ��!XC���s6��k4De��kV7eǖ�jY�2�����ro>ic�0��[m���,G��X���T��
�E���y����WX��u�;�n6R��8d0��m�j��BʋO"�&<�T�CU'V��;�X��zs�}U�1�W���}EY���H�w9�j�U�Ŋ	�����ݧ����c������u)���ni�eŕ��S�丫�iIs�B�r�/�a{!o��M���M޲.F]�� ܲ��{���K��}��Iu>�z.9\h,���M�HR��0"T��㉹�7#��r�e�%��L���KK�"�G�0Z*���1�mI��i����3���5��$J��[gk�(n����VB��}V�7fuEf���w�u���O&��be�W[&kӴqQ�D��|�c�L`��:�3wy��,$`{iwa�޹����Z�)`P����(�ͬ���U���Ut�^�v�6m�&��̣�=]�r2�YC��Sv���1ʙ��Zk-f�ٵ���3u��dVm��6���)c:ũ��X<�Y�/*j�Q�Xɒ��p�QsEKK��Ys��G7�̺n�S�E���}G(Z�MU�K�)�9fe�}��A��u��cdƛ��6i8uV��G�+I�����JJ:������f���k������x{�����������>�����^I������o��_<]Z��xn3"0ʅ"IH!E�m$�0�IFO�'?��e�O���*�Q7K|5��6(��!�M�nfD��((�͆�pq��of>0u7\ͳQww��!#��������ubwn���G���ˇ�����mɥ3s*�oђ�JcWY=�2+������f2��g_:�����y�S˗���\���p.�ۛϨ��W�b#jb� y���M.��w����{�rVS���,����O�P��6�n�Ɛ.N��2�W�K����wj�(q�6��\�Z"rwV&8xb�)'�HB�1�[���}�k�����{^L��!;[��C�󆘓��u
��qŢ���rk7Ff[|c(�w[���̜�B�$uTX�Cf���|i�m����Y��{�a�U�lǵ9Pk�6�GG�����6�+���0.��qc"�l�I������K,.Th��Q�86̂��v��������)P�bӨK"��$�Ux�E*�/��*�"9Z�'مm\f�Z�d�ON'�S5��E����M��u�m'�^f�X�o`���e�}�f�l�8����2�S&m>Ed�|-wq�{w�f����P}s:��wz��6N���I� a4p@��cM+f��SjV�i���Jm�i�4h��M+m�Vجx����iLM�M��l1[h���1X�V�cJ4Ɓ1���A�c��a��i�f\D;l0R�5HA!L��$T���Fm��%�)�0)&X>w$=�j���Չ��ضe��j�o3vZ��<>8p��ll�5Mؚ��O�㴍)R՝�yp{�i�V!h��*����ֹx���b"�>�l���ÇN���---KV�Y$�"�U�W,Z"�(�DZ��fQS^�Ւ�j,[d�%�E���ku��-X�?:�5�S�I��KRV�2�0�E�r�-�r�%�-�QU�����L����d�^wIRT[ڹIj{�%�UR׹�i采���ÇNu�I�[�\j��1R���2"K]�<�D[�t��Չ�yדx�DR*�#�b��1h�J���4$�<WI%뮤�6�^�l���ӧM�뱋]��2UՌYV�KSL�锦��,��&��,�OK�%%��ч�1a��2G�7�M����ӧO���Z���ygj�Ǖ0��1j����L#V]�y��U�&���VF�l�ӧN�w#�Ҋ��d���������-0�>W�Go�׌��Ս��J|=6t�}>��G�',���O�X�[5ܑ���"Z�U)���ӧN��؏lCԹ̑���VQj���7S*KM�'˵7b�5��Q)<��n������[�4�kz̛���/����hƢ��>�z�sA+ﳺ�Siq���?9;��;B\�N�� �ѧ6�i�ʲ�k+Y�o{m���������3�z�4�ӟ����.�n�
�(�	��O��j����~�;W*뻎(:�]�*�+��Q��$�CA��/�l�ᾞ�����g�O����]�8nFG����}�.L�ʾ��)i��}��a���	�c�ϫ�@\�%�=o�tzx��ǈlÇ�	��ş	��ʚg��D ��u���>�}�>Θ>c����T��`�Q�f��G)�����W�'�� �{�X.���`��͉Gq��iC�O��?|��r�w��'�NVqv�2oj�����G}��a�%��n��=����y��bI}�\	���wds��r�oc������"�P�>QK�w�(Q�����wO5̜�>�wN[�",G�fy�a�d;�:���(�$8l�rzb7g�.�[zf�}�����{�=�k����������jG�N#��g��8c>ͣK�ڏkҥ�"���N����,$�ln�UF3�k�J�w���ۗz��W�T�1[�mf�\n���G��׻tc�z+����IX[��/l���������Ž;��;n��K��wN��G�}Z�_�ꍁ�[�Ia�st"�qqP �{3}ļ��׫��Lo鿭H7t�� �&�5���r	����������>~���:+�P���K�Dp�F�q�<��;��u�8�"�ݰ+=��jc�o�{!���\`]���B/�+z �|	6L�wK����I)�O�w�pf�'�kܛ���	���@��I�11�31�i�uv���p"�!CB,9	K?�, \�k�R¾;��
�V���g��~�1�c7�fdgn��,�ds�݄
݋wȏ��+�>熹|�fo?�T�y�e�Fb���v4���g�����7u`Y8ׇ݇6U.��xrx�J�j��7/��9Io��vA;����7rf�|���T2~�y�Te:�4TiJ�#Mt�oc,7f������E��vV��i��=fIҦܱQ�Te�p��#��E�z�C���sj��օ�=�u-!�:&����U�c\.;ݺ�XM�T�r
D�f�<y�G��;uwddr�nw('�����@�왾����ppw�`
��'�B�h�>��T��/�}�D�p�?�g�^��.���f�w�vZ�[����\�]�QJ���G�:��Tdm�L�Tf�Ƀ���}a��q9-矜X�o����.m�a��`G�7�r���]ٮ�@�Ł�H�}���1�"r�ϧ`��a=#�+�����ko����'x�.��KϪ+ޟj�2=��nux����6��M��|�&��{����lhaYdQ�9a����79�}Ņ�+�ΨdUi�2N�8��R8����x�z�ߠ��"�_O�C^��&zg���\�5�9�ٍ������ňߒ��u��B�k�h�z�;n(�;��0���'��{/r��}�Ng�O��[�U�L�\K�Y�r-]�_�l-�gkXtֻAm���v�EP��,Y�h���׹:zt���JW��I� �^*O�Um�p�[�R�s���-��Ȍ�r���~N��53��b��&�Eүʑ.�:��le���b,�f���+˨��]=�k���4���&!���~�Fĳ�tw��r�c�Y4@vsf�8�ɫ�{�f+��ٚ��2VB
��_q�a�*W=H'!g�`���v�՝���34{+X'E��j���h�l �����]����0E�ǜ��4�m�CwW�x�ѫ����>��\���?�������>�P׼��v��+~~�Ϥ�o.����!����<A�V�m=��@j��eƎ�>]�C8���9��i���0]�X��i�<U,����6�P��U��9���ƀ��~�<�K��X�>�oX�Q���W����<[����R�qs��w��N��GGfFv��7��[{8����;�o��VU�?���/'~��o�^��z��V���]gV��[�X�V�c�����L��im>:�u�=�&==��*��r�>�����W��A[J`���y-�F~�t �X+���!@��p�+���*k�O��F|�WϮa.{�R�fsj�]�A�ZͶ�o,��œ�tV;�σB��h"�P��0���RPT��(J���W�:���&��������㞅Cy���z�5�"t���=A욌���ޓ�;�*f�?X��C�e������<�^�*�[�����Y��L���X�
�itO�/W[���j3y^��zvh���|E��J>�lp���_t@�� ���f��2�|&�ׅeJG~&f\�\��%,U@q�o�v��+�{^�]�xSCF��<R��d�ܹ��^
u��93���e��j{�V^���N�[E�ȳ�qþs��؏3�h�-���� �B�@�V� 3�[$׉�ޒO0��g�x�e����Hj���=��A���!�[����Z�w^䶎܍W� \�۷���l�7�X�0�:s�zg�U�J|^���� *~yn�)����}�U#���U��gL�g7lq��F���4sT���ᣇ����7	�g�˳A�Z8T�AT+�YkL�oU\\��.����!�n��W���Kނ�	X��6�F�2��@��7��S,׀V��X ]�5Ё�t�������'�����:�U$2f�n��:Թ���_L���;���:�3VI|�U�s�nw-�;����/��p�ΟoH瓔N�sj?�fv�w�c}�]>��<�|A�9��I�����9�9�y�.I���x���M�Ve�ӽ�*�O���p`7m�f2+�$��7��@n{��M�s��H�37��.Eu����p�X�{L�d=�2,���g��Gj+:&��O�vpŜ� �~��w}���,&��� �x���u�Z˪�zw�k^�ή����%Sg��T�2�՚���h�_��5~�=}��Gw0�� �t�G@X��l�����r 9[�=`�`�i���=z��z�ٛ��+��<�-�fś��r�M���I����ca�_D�F�5�''���_������i�u[�(+{��x7�ǽH�����
�(
�r�l�������+
�,� 
����N{(O4�xD*���3p>�9E���y��<�����խw ��U������#k��l�pY�U[˺a%{.���Ƞ���V�|ؕ��GOk����ϋ��k�We��;�j*�ZJNVw+�7;]Ǳ���vp��gM�柭�}5�	����#>��,��;=U%�M}��9,�ujT�U�Gnoce�"Ɛ;l	�aě��q�m����`�z�-rx��I�u����~���sR8�Q�:ˁ��nꉳ�K��Q#}+���w��5}��g���x���8썎9^�{�Y��w��'}.�#SyZ���<�[�_�am�f�!Ȉ�DV$��8�4�o���f�CL���{�=���MK�_-�2����TA�?T�'�Ã`�|���Cvv6g�E�u`�Z��q5$gіO�AnΫ����v��dp�6�(��q�F^wk�4G]i�6@p�g�'<&��U��kscg��z@4Ǹ�:t`"���Q��^�r�b�gkS��X~t#��}�Cg�W���v����>vSΈw���]���ٶ;���
���3������e\����r�C��5���z#~JQ^�Y:m��ýS��gxݥ�P�Vi�p�� �~aC���(X�g=��*�=��F|��+)�e79��:v�p�K�e�ɦ�GM9���m��yΒeLx�m�� ��C(�H5��s���e��n/��>�t��sb���:�Wcw$���[5g{�u�7H~<OWS�B�������S!�S1Kp�͓3==#�;��E�h�_��[���:�|�R]�Ó���P��ju��؃_Uu���B����ed�U�H�o�`�Y�.�'|F�bןR���Ǉ2�o�L�p{m;���e�;5C�|k �.u����[�Y�KW*���������S��7鶾ʭ 53M���[�ޯ3Xܻ�?y�h׉����`&�d��6jߋ��x�b^��}̏mr6ޞ{}��+߄q��h���!��p%�q�w}�?[{�����v�}�熯��x������T2�����(�⩳�"�}�χf>�5�Ӳf�ŷ� m_�P���LtϾ��mS�Ͼ��To��mU_�n�bK�tv�n58顕W|��7cM��L��^-��Nx�I]E�1������'���ǎ�y�v��Λ"���dDCA$��o.��-{�'dv�����Wmk����0��^�t6e��Nv�R\߉���=��ǭ=cLiU�cJѦ�i�A/�l�
$�ƿ�!/sn�9"Dx;>3z����=gn	7/���r~:�^���Yٺ:A퇝���~�o�Nɟ<���=�L��x�S��inDl78�{�m��U5/�]ُ��W#�x������9#����:��������}�멣ń{R�ߚ� 1~�-��p���q������u+>��c�,Ϯ�[�:��e�ӭˉ���K�t��)*i�~C1��/�G�`,�C�t+]z�eo�
�;���k|cћ�?	�G��`�|r��x#�W��(s�~�gLwú���_�8���X5�/�C���,�w
�9"��|��C��E���@�/�$M~s.�r���X�:����#n��QӰe�4�h�"��Az:��g`�m����&��x��C����=����y_-DY����X��c�V�'��~��qk�����g�~�mhă#�C�k�(���U���Q�d��`��
�������}ٹ�<D��C��U.Ŵ���Wkӏ�e���rd؄�P�}+T�יU���b��;B� ��<�j;��ۏ�N����y%VUK�*��q�/�����Y�(�ɂ�5�>O�<�=�\K`��s��j�z0�y�^j\�`n����w?Vf���#��ŀhO� �~�_cc�o,=}�M+l�hg�=�8;��>��Ω.ⷾ��`�0Zo�_�'�;s�מ<^i�uuzM�}Sq5"���W0~�n}׋�R��5����ƶ!�}�̓���Ӈ���a~$���Ԁj��x��k2��^ͣ��=��sSM��=�o�]�9��	���2��u�Ϫ�{q��hψ`�S�<J�2��r��|fvX�4���W� sK�{ހ=��=��.E��[��\��d>�zeG(?������>�{@���?��P��oz�u_����d�!F�3#:��϶s�]UGR�c�;ȕ#�4=�=.�y�(�!V��P�7��k�A<I�\W�3ˬt7��k(s|��\9�h�E��6��5#!������9�{K�)�VWc�t^,��o�m��ܩ��_\�mf�f@�@�a=�=�m3e�i	R>�ŋ�/M�3�������w�[Gm��\��M䛕i����V�_`�zE�4����f�h8�o�wv&�;݈���$�cF,�������O��WK�g+�\��Z�U�x��&\p�QN��B��T���"Sw�ؒb���:"F�%&"�]Q闊��W��Mb�H'���V�	�^mYmi75.7�A�ŧF�n���ۏ���ı�t��gz�%m�*�ج*�9ν���=���Mvwr��ݚq��U}���ȭG�-���\�%1�N�{o.��j�fb=��9�L��Q	Dg��s�X-�\v�u�Zo�J7�(#P��o`2��j�]�W*���98�<��+۵�:��͖^�n��B��4L͂�1Vf��C��:��FxseT��:�C�֝�Q=�{ݹ..t^�����s�5D+�Ԋ�l��\QSޣ����%t�@��5<ܷ�'V.��Ͱ��:��]\�z�̈^�����v�-]^����R���F�y;֓"��c����Ϟ*�Ǯ|_�6��#�C}�Of��x`��ʡ�\u��S�Z�ɣloj�Y����^�lm�"�Oď@>C�g/��J	]�{A]��61�#z�e�1���!�·Su��&aF#fdJ��5l����e�^+ބ���36ɋ���.굈U�-�;n�>|8�:����]s����N}�nk]�uC�ݗ]%���l��X��C�0����v�=WT]Ŧv���t�!�����"ښ;��㴯N7͐�V[���M�v�G�ؕ�դ#9e�+z'N��g/�DlL��ˡpѥ�;�3���ßr�+�-�P���8b����Hf�!�.�J���Žy͸�3�qL��\�����y��E3 :���AwM6�5}UZ6J�6l���&E5ѝ���[}�y��Z���f8�]L��3�z5�uV��uv6�گT��.��Y)�Յ�Yk��6�Oj��I��gb�O����I����R٠2� ��yr.F��bZ��*���Ùz[�&Ku+n)�s=��N>B;�X�����vI�Ugf��7eˇ���ж�3�w��V��]k%���Ç�mb���[��D�m���\����ښ_X�Ln!�>�mܾ��Z]�6𹈺�ί��a���o.����������㏓Y�������Q�FYDj\�B�31>S6xxt�p�|�,�����(��v6|���;�(]bKR)��F�O�N�>�ϜX���b�Z���_���DnX��nV�s�+�h���ӇO�)j-�-폐�_~�{�r�Ahر���4i��:xzt����q*���j{����oMp�V�$��Օ�0�����ӧ�{{Qj��d�sZB�eG�F���a��������'��gŃ�-nɖ%�>+V7b-��xt���ӧy/��|nk�U˛wuưŖ}R5cG���O����'�݃�I-�|W���Ô�����\�5ȫp׷��`����
��yn����<ImpcE泃�V�t7�pNR�y)u��Ys�3������ŋ1�J�|�fb�a��;��K�S��L?1�J~1����`�	�f��C����ے��:n�24jp��\7�S���Ӏ���I���Ͱ��g�;X��z��w�~�˒�%�_F36}w>ц�e3���ց����s��._#]��	�!�0l��77$��#���4�qK��x�����O�]�;@�����U�Y�2tl�Vu?{�>_�e��CQ;�	��+b�v��A"�b�D���Ϩ���k�1@ƴ��ٟ��0|M|>�D|�����V�<�q,{�|��[J�V_�L ��CheF7�Z����]�|׵oY)/;�XN<^����64�d�w �Dd�m�P�Ϧ4ɯ�_��hJ�,�!Tq�[Zq$��+d���`w���[ױ�{O%�b�Mì�	�u�T[��we��!�!����F��َeM,�d��9�w��>��b��
>�	��#��z����W9.�ߔ[�c�6�V���XE��O�C6S�4�b�cq��a��p�4�~�*�i�]p@�d���٘@�7B{�_��%����7�g���}�
k�Wp�4��\n�N�Q%�pr���܋��׉���!�e�l�җ7�OW���d��5s�:�����|�̂4�'��>�O_���t�7�'��p9
�1/����Lnٛq�	�(�O5����<�3y���������Y=�*)c,qtQK��?=���ߪR��QP`�w\�ao`G�Lk?=>��O�6�� Asj��Xu�*�Bo��%N�Gúd=�w���^�߁8?`����y���ǟ�i�ΊT]�ޡ��g�*����YW"�䦰@�&#ߩ�{{����eW�
&X���3�	a�+�-�(��m�x|e.4�PǤ�#L���%8�=#�Ӗ\	h�i�ŋ0md��YR����"��=��3r�=k�6(h�Əd��� >�X�uNK�m��κ���Y�pZ8�������юs�x������u�(�N���0���f����oE�����s��p�j�?A�,�|��KKK>�Ɩt��)N����b~�<{m��V'��lu&D��~,q�̟/vG34��L�M�m�s�m10�/fD�G�OR��qm�F�B۶��]�6k^�b�/#Y�1szD=^�/y�B��'��z�@?���]�Y�u4]7��f�ޮ41�J��]��	��u}+���ʇ�߹��Q����/E*L^)�=f���5��a����!F����ۮ�D<�+iB��v��&�܉�y�W&Z�λUY�U���$ZS��S#80�dA�&����i{�c�I_)H�̺����{���jJJY��<S��U�.���7�Mb|�AZ�vO!`P���*��F��1T˦[��Z��Ǜ�7�V�����X�X����R�T¡J��Dz�,����'��Xax��T/��� ��9������6�~���_����둚
�����iq�=G6>U^�#��i� 3aۺ�-�Qm0�LY�m7���g�S�`5��J�=�S^4�E?p�������B����Nz�1��1�4���F�3����p9�f���<�櫇7w\�b��׶����s���\�7�)�%�b�'�+�Т�c�v���%�cH���^���Aѭ9Q��Ōk��O4 �:����EJecL�m�����ř�Pڠ��?�-�������%�_G<�V#��M��q��+<�0�Qm�G ���5��G)j�R�Vڈ�'U6��M����*�~o3�A�X?���V��� �)��YQ��)��jV^)iO��T���R�Ю�c;�f�s�Sȗ�Oq��IH��7f=9Kz2��Gu�u���ޫ>?~�A�D��a���������}^��-0�C�r� LPv��@�;��e�r1���O@�hP����_��'��_��
^rd���tA�Sg��s�]ˆ��nh�HNIz�roӹ�yvVZ���bh;ï}�6k�P�.o��t�`>	�mէ���@x���m���4��^��Wy��f��l,���t�%>���0o	Y-t�Ϛ��w������'�?E��y,�aAJ%,'�R�n�
� ��ӌ�	mo��6c8��Ù�G�g�w,���"=�ˤD�S��%M��|�>�wg8y��a>C��VB�DgDK�_�����r1��,�;��C�Z���˯u��,��"����U�^�~`�!�t`uq�b�5�E܏;E�(���>��A� Kh/z�!h����"�u�ɳy-�v�O�Z����q�SQMҔ��C��wH,k�(V>m�����U{+J��/!zz�!�^��m!���E�K�boY�C^(lSO�G�D�nz��fʩ|2w4'bm���[�?���+}�_�jD����(�05�+��Z�{�����<t�~�v��ဆ�ך����rٗ�,K�ykEec�<����
��+ݏ~0��v��T�;	-�rJ�9"G<�9�:aEW�ǻ=�Y�aY�y�Vs� l�6of�ǣ��Wg	Kc#�^}2@����y�+�P�^��'�I������s�p�+��:�,���ﺼ)��/߫��G��-@A�ה��J9���Њ�:^�b5����n)�����x�9?7�d��S�o�����'�A1Q��u��(v��lj�R�c���������R�[���.ݎ���oX=�{�o�����D�pJ��y[���du�M'7����Z��!�*
YTZ����2��B�!J$�$�r���R�xio����#`hla����@+2�h����k���B�N�p�T�-z������s������9�����Pg N��A���}�B)��QC�<�E����8����g��4Q��"�Y|���8��h�]��1�i�@4 'I�K�Ar�2�M������cIt"�c2rr/_�pdx:׹/z�','�
 �LU����CΨ��B�Yy(Hqa��#���sϢ��S���-B��K�����O#8<�Cˑ��Η�2;�y���*b�Lh��M@K�LV;7�Q̯a����8#
��c36iآ��inK�}��ÔK�,%?&_���O4�k����6ty�7��}QJӫ����V˯��Q��V�~��5K�ڑ_o�BҘ��H��_�?�E6�� #>� ��d�J냜�k�:�N'�[�OX�D����*J�����9R*�7�Z��K��Z9v0rN�S�O,�pd�uɍ���
m���b��g;X_7)YN�`�l�?rm4�S�}=����w�wOu;���7�7ΩpU�cZ��o^�i)�S1�ڢ#%tx��.�obd+{aAc�@�t�e���٥7��9��}ם���x�T��k����kYą�͋x�^�4�T�V�.�Y0��9. ?����� =�xPIJ$�0�$��%,�J�R�$��}s����5�����;Y�=���^����Xe��SjQv��[;U�㬭��ʙ�K�A�̋Y�#��^Y�M�Q�D�� �Ml$���It��%Bbo�*k�0���L�L|o4�jZ����G����L=��V<a�`��xzN�-@K���G�8��E'�3��<O��ڈO)�+n�GT��t��F0�&5��znjOM]�&���&���f�o.�YU���م؊��ݭ���� 2h\��M���nD󕮮q���m��\���Ж[�^�-Æf�ɬq��)��փ���5��d~�����)�׸��LOm�?u:/,|Z�Z��e�{ߩp��>��<�Q��L�`���<�*'b9eS����o�߅b�	U-5��u��P=�n�|�_oYc�t�jKn�-g��X���A)��[�F~]�2�Q0����o���g�7WK@�P�R&��8�:is�E����r��b����#��Ȝ����0�x���D�{/��^� �����疄=#:QE,ڼ��zwW��x�꒍u�ZQ�[�ݏ&��k:��̪K���U�\P�d��
�m�?��/�F��<(�����r��<�˺��7��^X�6is���s��wG���jQt���5����q��cM)�h�.ks4��cZ���D~�	J�E(%**"%(IJ�L�(�Rv��H�~�\���}���u����Ld�~�S�����|]��_L�@��ɥZ�Y�~Lik:?O���ܟ�V_��T����*�5����̽��č�����Ѻ�sx���y�S��� �W�^��3��Z5�q_5l%�k��e��P��c� f(1���z.��ͻ���5�fq�u�z��-ˣ�b9��/LJ��/t��QM"߃xy�t4	����jkW�}�����7*^.�h3��g�_���?�Ahs��2��b����eMFH�!��#;xWn�¯^��#�N��yǃ�z�� M��`O��%���>�kLx�6�5����<]�s�.�]b������|w�n 
9W�5C���W8fΙ<��[�ά��xG_!�:�1L��
�t�f�ly�ǜ�҉~\\�M~k��^y�:�*FoK4*Ȭ���G�!vB��y�)���M����0ͩB������z�q�V���)��R� &�~hO��F���}ԧP���0,s���~���>����
֥M��G�:�;��ܧڗ_C�����m���1>�pJ��4P��q����J5m�= ���f���3%���.��ǀdxA#A���ێA��2�h�.�/��wJa�*��Vm^BS㜕�5�5���]Cj'��(;�5��۞s��ײ��>P?E")d"�A)P��$�$��$�!2�y��}�����Ϟ�;o�t�x���'�<�_ەhػQ�Ċ��TxX��0�,�Wg=Ae�ε�맲�W���n�܉���%~p�
�ן[�>���S<�����taț8�����O���4b�%��*��L� ��
���=�yY��}B������)L��ۭ<�c޸,\�7���By��}��E`��4q1a��
�<�B#��'�g���Ӫs�Ƈ����$C�W��ܩf��8���K0/HR�����/���\~3��� PgD��c�;���S��ۼ�[48���=Ӡ[�{���qXsq(ˢ�oC��0;�$@�����Rm��D>���E�������;F(����< ���p�\^5t-ju�;�O����ѣ�PY(���6}��j�=���3�<wH,j��|mЭ���}'�0W�O����̮*���:s�g���_%�6O��.}��D�J�����R�7q4�s������@��an���֨��9��K��~
�1�>�C�7u4>^s�}Tu��P���X�LUz9�y�Ա�G��z�k�Y�gg����Ct�ĕ1����ƞ�M��IF[�����j���2���\��Q�7C����gq��}����I;�9�i��K�4MR5��������>���I>�%�#$B�R�B�$�)�B2ȓ
H�v��������q���O� ��j���QM�Ͱ�`Kt� ב�+��<�G+���9ۅ�s�!�]aL�^L)��5�2�nH�as��p$�a8U�buM6O�M�wE���q6�e�7����ܞX��u��:6}Q�7�5�@|�+�q~/�zm?6'�~t�c�I�K�,��}��S�|�U�aO�$p�����}Jx���gR�� �it�洚�!�u8�ݗy��Ã1�q���t X~G�\��
�'��%/|.��̷H̙��lt ����@P ���vi�0���Y���!@�B�g8f�shP,/��}A��/��㣈�i��D�ܓ�^˺H�܎O��<L�;����#^��[�A� +�т���t�E����bY�˯k�=�p�E��곏�]h��D	b��^�9a<P�GI�wQ̢,��W�o|~��|��4
�Ň�g�lX�����m�\�f/���3�f�m��W.�v��ɶu�[�k�C���/���̯�^zn�����`��L;�9V�N�&5�6I؜�++-_�B{�H7�dVnAܜ��[�wmɝ��ϩ�\:�}<u��d?ЀGF��Z��艼N9���g:��Mٶ�p]���mf5��p��]V�>��44�I��#�+��?E�J�yb&'ڄ�XHRȂ�,�Y P�� ����M�^�z�so�ח}he����y�	��g�������_D�7]�]�z��Bv����y
u��p
'|Pp~@iJآ�}�ɨ�H���e�5����ukmFn�s��b��	o�� A(~|�N�|L�|��e"'��7?r�+�o<�Ê���.E3�h���&i;e��6�i�R���u=� S� ���b\�'%��Ҳ@	���a�|���J�:��qtљ7RT''�"8�Ȑ�b�B�~��������/9M������J�.�[%6�ݬ�7�숂�q5i4��]�=�-�e�ڄ0�"ۃT�]��6ÊͣF��Jx� k|y�ח&�Y����c��U����Ǩ5���#@g.͸.<s��4��8'���ь�P�����B]%�o��$;���l���r�5�¸������~�3�����J�Zr;��}�n��H�_Cya�z��w��@��ԑ���4�6|��x鸸��xy��*�0�q�@4ۯP%����.�4������B)��P�A�t� ���(sT�O�|&l!d+j���s,�r��o=uk�������ݶ����C�-*ʊk�����M�˙�Ԛ��-ud<�/v.���S���n޼���Է�YL��Ā�<	�P�z:oe�-�|ohY{z���6�UU �����3�*���{$�Ep������`�5�(��_�ᡸ.e!�փ� 7�����ܵ����Fd��cpʱz`�%
z�l��,�޽�;z;�7�Ԧ�
#Z:%�[ͦ�0�o]�Q�����sy�����9Dh�yۢCh��k�g^�誄6���+jX���z��d�j����FJ'c9m�Y�8�-�"T�ڴZ���:�j��S�.ή�G^��M.���w4�3u��'m��V� �.���r�=Ҍ��xj����t���=���u{F��H��d>E�:�{�����'pW�H�0�e��L}dB�Jlw_;���mqW��:�!"�x�����I��.���wQm��E�M���ksgt��L�V��mA���Gj~�*I[���%=�Ġ��v󯰓YK+s����^V;���e�؟7�u�3nT�8t��e
��(pomP4��gw��ŕ6l9�pvD�6��-�̾�G��m��QWv�X_[Pڋ��VmmN��3�Bϕ{נؿH0X�ru�(XdH�m!$Q`�O��aB��P!5
t+DP�����p �?Pb�₈��H��A��b@�`��tՅA���P`�^��Ac�ǆ�|��G�!�Z�s�K�Tc�h4�]m����ŋ�A�B�"a���\5�XA���I�Ea��j9�� Ԍf%�	���9����X�h��md�j���G`�G*��.p���}4!��H�W�d���u��&�W["���L_;�.��6��<D�z�=�f�km���.��W�a�Ǹ��y� 3�6�{��/�Q��l�W!ś�w��ĽZ�����v�8I]igG}����o)�����S0�wb���mHj��@]��ʽ�η`Ĳ��-��WʅGbm����7��Je���ER^2c�]��۵\�U��ns�TŻ�\���Ўnڪ�޴b�4𺤹꩝�W��:�._og2�Q���D�N���\o{�Yv,��BnL}��v捲�U�J^�cE��Q���o{b��2*�#��y�j��vi~�>����ʎYf^������uenv8b��Y��l$�v�N�y�(t�vv�/�#&��x����
� /*]�m��L�/��wUl���M�BA�˽%���y���wz�:t�u�)����T��3�����ӽ�m�X�v���ɷ{�S^Ʒx<^l�O.��30M�o��7����9wf����<)";*Qr��Q��׋,⬭D_s{UL�m���y@�{��LF�Ҷ�ھ�!�[�ҹHn\�J�s�d�Ê=�}9�<�j�H]VV5�Op���` ,6ޕ�R�|l�i�m�M<cf+Li�V+m��M�Ƙڶ�6�4Ҷ��ѥq��<<cV4m��m��c��ڪ��6�LV��l�ccl`@1��?@�)#-کK$��m'�3)m�I�Q�6�p��Ċ�e0iĠQ	�Bb�(�H�����oS[�\���Ԟ�d��[lOn�J�9�Q^.m��^��^�_���:|N,�R[7�j[���m}��m��x�?7o2�u��4|>�:|rdO,�ci4��U�<�}ur���,w1Jt��zt���+�V^�4��cb��s+���zt�R�W��8p���Ք�*���+)�龛�
�;W�o2�����ܔ��������J��9E[ez�u�ƓF�K�sk��8h����ÜZ�fY�X���77����k�x(��d�d���Fχ����r�e�{r�gtl^-�x�-_mr��&\�ɗ,R�4t�zt��9e������kɱ�����i�J/wv�Q���F���EN�c�i*�$Ki������{��+Z�(�`�b�w'Y�5�_[�v]�BU&b#k��`�u���ֵБZ1�O=���<1\uXƌ6ښm��ê�q������Mow+w.�޿h���XAJ�)Q$��Y	���)Q(  %���h�00�E�V�x�?��{��|�3����L2�q�����]q�k.�������;K�h�d��3y�',�\0lO�r����!�ϽdH�
����s��m+6��2�ǚ��b���7���MP�~�A��W��#_�y�Z[�q�db��������ա��U7j�a^<�%��P�4�<�"�Nz����"�<N�p�ٌ�
��^ϦzF�[�u��[�N�O&����k�!�PZ|�%�;��W�����X�6	��+V{��y�*3�wՑ��K�x��zB�;@���u��3C�`��@���>���󟚚�c�i��R�!0��S�'��ٯ��|�Pe?��9�X�/���8�ͷ�!��m��#A$VÈ��5��Y]a2����T�@�"��7�er)�%�1A�B@��b���b���O����x��o�c#
Y��L��|E�����ww�`�[K����0OUR^5�>g�{3�?�<4҂�td�x��r���@4��K�8�7�����.����b{�H�ď�K���;1�N%0�������i����bgr�(��UV�T��:�\�5�
_XlU�}��k��Q[1ח~4=x��ϧ^�e�#�%�;��F4vP��C���P��hK����.�жw�l���8�#L]m�۝��m��A��u:Z��J�k��S�v�U�ޛ�;'���� T�rȓ	%)$݈�T�	)d#%,!�Q�=�+7h�Ľ��z�L��kl^�ʹ~y2�u*��(<�����w���%����nD�,��n^.�^A��\ީ)��E6s�x��J�wA�L^LgP�PU3c�_��9�HG����W���(spj�I��Y2}�S@;P[y��.Ԡz�w�un.sC><��*ޜ�n����ލ�w|����x����l��Øx<��ZS#@�มԧXq�o9H��	TSsM���MUQ���P����4!/�ZX |��!?&@��������
�_�f������Ƶ�|L�[m�3�#5nq�@V�ìLC�ÿ��(3��G�|���(~����g���,�sgg�3Z6��>�w��h`"�?Z������S =����<H=�&4���(u�D-7����ߖr��F!���7͔��%�`�	8�M8zi� ~o���\�8����#��)��M̅;��I��������}L0$(�E� ���q��vPs2������ت�ê�P���=��v��a��x6?�c8��G�v��§�61��,�=Ҋ�����Ո�0o�W3�g���:q\��YQ�f�PSt.���Aڍ����p5@լ�vL:li`.��g6P�N�!�Ly�E�EMR�\]G��L��6�ՠ���d��2�Ѹ���gV&!#�VUU&�k������HJT�r�rB��,�R�J$R�R�%*!� {�ʖn-u+��}��5~`쒁�Sь"+;�M�)߇���� Q�$H,ү��^B�8n:5?�(�_]�"��@p�>4h;|���5H�6�<(�|C��g̨z+p/� 6�x�v�`-�hq���mAj�"�[�f�4#�y3ԿiC����]j+�K��+�⚙���hn�3��|����uU�$��%*�T3b�K��6�u�Q�Z�2n�d��������=rXO����j��*:T@�q��(G���c�`����v���v����k�$"5����ܙ�<��&D&��@f�v&��m9�$ͷK��ȵ���Ck~���������
�A,=0�@lx\ջʅ�;�����!M��ZQ��Ɓ2���,bUٽ�Y$u�ۖ��w��yf��v��$�bL�z�ty��N����<�&�t���9t�O�HX轷1mw��=,h|����_�G�a*b�	j��Gf�y���N^�-(	��d\$b�Q��p	��=hT��f��6��CdO�~.�6	���4B���;�sy�)�Sn?�r�u�oi~̵2�n�/k�n�[U:��[�+�3�8�c�u�s�'�n�`T��CH��"7WCٯc6,S_��I��b~�gu��->+{��8u��U��&ćs�w�3zן;�w����A���Ol�a`JT"���H(��0���գ��+^��K�:��C=�W0���_�TO����pAȡ���X�w�_o�a���7o�],�9)�"]1�c�z��m{�OC����i��xvr^��J�p���~S��Q�7/'�^�`p� @)|G��"�X \2�,$8^�O��l��Č����; �,�N���k�O�{}��}�dPE��oɓ�a ��a.Q�sx�1��ʏB1ۑ��ms���Y��A�z�%1�[,�B��	x�����P�`I&r����� ��Kcy>-~�1��;a����͝{��܁܀���{��v�N<�-{�K�\\@�A�8�9������8Q�t�V�
~�)��-�F�7/�,
�����d�fOD�O��i���d�����}�������A1�x�޹讍�� N�km�Lp���i�kca��t@�,d�����Κf��2��Ow\�
��@"2L���Rzm����P09�������N E��M�E��H4c�uZ���f��I���;+�6|"�~�h�QL@׹N���{az��3d�װ�H	�\E�_��c�6{^�2z���C��J��=��R�k�StF8��f죽���; |k�b;b�k�M�ǘ��µX��h�kle-Z�a�!@�(z�0(HՂ�4So�L�S���b���Ι�R�-k�u3!{K�m�n����,�S�F6>��U�1���m�0 C�0�J�޴m��Y��G�~�R�$��e5YJ�SV���i���&D��uQ:��À�;�/D�@��!�㕌$pM�c���͌2%ĕ�?��,KI��9���^㫠Js<�O%�T7�5�/tEs��_�5��U�ٞ�����b?�"|��\��?�u��E�J��]y�ݗ��}oL�s��@�~��Q��]� h5��T�'��٩����z6�_K�b^v�6��/3m�"���?��Idܮ9�
Ng�-���q�d@�T��7^ޗO
�d�m�m����UB�y.��s`�ExV��Ǳ�c�{7��q`'�|����v���{O_�p&��D�6(y��;���
�h�����@7���)��d���$CΧ[�wط��{Տ�|3��$XXI&ـ=������x���#NH�SyGe�hSP���z�E�xSt=���Izv��ج~i�~a�? �G�?��0|~�l��y�N���kDf�FTuX�O��z�������ĳ��/b��V�=��$D�	S�!�l�7a����W����31}����T��>��"`�>%���`��Ҝ���~����+�=�p�����X_��ӯfd�C����.�ջʯ1+�d����\�����lO�V��e�Z�r7�߻�ov���\#�I$��|�"�	ڴ��gU<���F5,Q��v��F��F�S��t���X&0���{~� ��� ��)RL�RL*%,IJ�R�RęR{�}�~��:w�?Kf���1�hQ�V�_�3w��}���5�NC�1N�VP�b��׶��p��m 6����o��n��7p�B�N��BQM!ǽ�\P ��X���
��vg���N$.j�p�^�:�e�;>�P�E���w�{����B�F�9����co���<��y��Y~������}��,{I�B��k�� u�1�b����b�� �^��^7�9����r�>�����0�\�z|���X{H~� ��ɔ�J�
2�~$�cO�6��~�,��3����Y����  ��^�������wƂb�s�>�>�]��=-��)�������pX�≜���������◀	����? f��ML���M�!��0[y�tT�V5O6�
�@f�(憡�lC���K��"K������ٮ�((Z2= h�`��N\t��v5�#`s�������������i?���@� t�V<��
�V'����dNj�N.�AO6��L��|�U��\%zy� �& �,+<��|I�ƆW
)|�ʤ{�?,|{���3�>��LB�
xs���#.<��O���?'�zˇ��o��t��ȅ��2�w1����A՛��<��噙×eAԞTZo��_&վ�RS���k�:���Ыj�w���R�f)���SWS����r�����'�
T�JX��
Tybaa)d�����?>�_���7�"�PNpx`5Ϩ����o@C��A1D��V?�����B��{�z�6������N�[����K饀����yN0"A��������H��̯��#��i�釞u.�兆�9L/C  A,����"r���>���#����@��y�8Y�{.1��!-~��M��e�BkՒS���H �X�jw�-٭�������g���^[�K�������CB�_��f���1�P$�Co�#_}�+��#�]�*�oh�Y��=�3�x���Yd�����t�_ۤDcKG<S9��у�ސ ey����O�i�BR,�匋�ɍ�:݉y�8|��:�M������MNT�vI�f�K?�~hC�T�����M5�$g�k+�>_
#�x�n`����^ĸrl�m�Vxe���O���>�� 񁎒���0��#>C��lgk)zC�sEd#^	X��b��E6�YXQy0=x�)䧚c"�}�������uC��z44٩��\�]0*c�y�0R�i�jnG��lw��p�7����,��u&
W�w&ԧӦ<缪2T��{7�ffu�+�/Bus���\۠,X�~aeܷ��H&wJ�n��d̗v�I��xj���s�:��釷VD����G�T�eG�_��I��
�J�K	J��3��a�L<�7�=k;y��^�{i����=���oH$^{!�U���C�+����8����(�N�q�t�9i�>/�b�a���Zluz_!:����q�F�c����%��r���9G]�� 	E��|�3����OD(0@-��ހ6o�lχ5�6�R���W�cP�
�:~'�$�;�!+��t�E�x��w篱��;�{��Kx.�R�N	Q`_�O5-�N7�ky�3]Pmn �h2�	�a|�����_���_��J�0Ҽ9���kj)�L_���k���g����z5�������6xe��[�%�)��� ;�4 %N�W�.[凤�#`cH|�8b�lz�=;�@�\��r�x�A��2O�-��8��{Ajvo�Na0�~]�!D,cc �-�["xDW�S���þ���ݫ��������]�'�;r2��ʱ�4�i���͆s+��`:�dJ�1���<(���F!a�ee�!��0?T^T�&G妒���?~p����$Dŷ+8�2c26��a���6��r��R=z�6oC5 �Դ�PzR������0j'a
6{����|���>Ȫ��Q��(���ç�-Jھy�أ�\��y(�WP�a�M����5n6��`���u:ސ�2vE��~�ʨ�IUBM'��<wlܜ�ipz���vfV�R�I8����rL�7���k�^�=�E��u�``A�����Vj�H�*nTaGl��K
X�.�¢�!�������ޯ�18X'.�~������ȶNȐ���fx���bZ�|�SayZnT��SV|�戮�ߎ�*��}y*��B2E5צ��.�AQMlCsg��X��NU6�[D5ߵNC�u�-�سa��նbpx��`�P��|kL��@�!py���c��֫��_�K�Un�}t
�c��f_4��/t�G=�+�V�x߅ c�L��Ϡ���_�y֡Cg��|�9x�j*���3.�$ƶb"�z��cPn~(3�� E�R����/2r���Bv�E)���|��~�R>�m�e�	4/���w(�z�Y�B{�����9
���V���8�[̕o]zV��2 �;@��2k��i�@�+������}��CcЖ�~X���I����$W�uw��QW�3��C$Jy� `%��7��u	�q��)�=D<��tc���Yԟ�y�P�"�I��n�Xïv���gp�,#�ГԼ������zdV����9���3��X���*�+r%�7J�۴8Lt"|��#��W|�hD4����� MY�P0nAN2�dz��JK��W�m�ot]�:w��[v��Hw_r�&�5v��CS���[ׅ^����sB�I�w�R�vQw;�<���(W1|EUH	������Uݽ�����!�����iX��fCK{M�yM��9p8E��qnD)CU�w����� @"���F
Rp��Jk{�v�<e�w��η��m 'pQK(_���Hڿ��/�uo���H�EQ��sW��_��U�I�<�Q1� M;�>�����0g�>P|����gǾ{�,�]�ޡhK����eT�r�ZХ>�007��4��4��gO�\�7�
��f fV��b��O�?oc\�^wy`bb�T!'�ޚ�v�O���9fh���	�i�P���'�npi{�a�K�B���E���fZ�����p��8Q߰�}߻�C�Li}���!7�S���xŉx�SZ������U7~�*.�FC�-p>j
��^���}��n�T�0|�k�|�@B0 ��"p�~� ���ip�D>uC�}ms�~D�A�kN��א8 ���g�W*��&W�����<�4�K��om�u��2}�l��[��4b��QvX ��v`k�����~9yR��<�v�}�����[��J�~§�M�-�z�ʸ3���YĄ&���3�0J���2�dC��{���L<�������#�p��k��Z���Vn��Ѭً�O� ��亘��Κ|,�����M�oM���q�LQ\鄝�q�q�w�VX�rUuI�frQ_Q��9�+x�:AF
�#3�,��E�1՞��he�Q��;XS�[�A��b�IԻv�n����HS�����%��"������hګ�Xu�2ޮ�η��!P�-b�!�F�)��a�$,�ה���I�򕛢�7��I��"Z��]{<��5ٳM�d�����9wɺOZ��{l\�̬6Z��g�E;4����G�Z*1��ԭsUԼN㗏�M엘Ƀ��ƻ`N�2�0M�(+;�����UN�{�zjS�5ӲgM&���u��{Wa=��<���s����4+H/r.O�33���.�1po�[�I9՗�m�ЊŌ_7�¤�Y�"����{r�U
�s��KV�9��mU��zV)����ٗ����9Ⱥ΢���*��P��Mݹ�ZvE]��ڥ�Tn�jr�t��h���.��B:����:n5Du
%Ns�v�6�����	ҟ9]o����J}Þ�Y��u���`�ZS��	��;v�R{N�39j4G�N�/��˰��R0-,=!��vs�cM���׷����S�N�+Om���y2���8�,�w��Ε����z�Yu�2�L�pݔ6-�/�аi�

~AD+6f��hi���dƄ� �W��u�`��\��U1 B�q{��0`��Ƌ�pA0	騂wԤ�Z�p^�1PjVj[�nh��2=q�5�Vn];f]�Z|��JJ�T2���������ܼ���opBJ��,�/4�L�dȯ��{�q'���*�9ķ���T[Puy��C9���ѕ�t=Ս2���mK��eT�\	�C�Ķ;2�78�!m�Β�M|���v�]�S�N|"6�t�r.�D�idL�K=/$Δe�,��^��]�vg>����{����ŧrC Ëe$Ed%*}R��u&�T����Q��b9v�m�8D2g6g��S���5�-��B�k}��TN��lkH��r�Z��+��MS9X���cYy�����/jH1�٫B��U�>��.�ڡޱ|x/LEہ��q>��V*ާ����U�ʤ�M���P�V3:�+�Φyjʺu���GFe��%TX�D�b�W��:�����}�u-ۤ���1����*u��M���bk3����7"k�s4��*�}�r�콸�L�M�^8O�<��Y1�w(��0���l�خ%!�ݷ�o:UK�_[P��1��<F���<��:�����U�Ÿ5M	����cM~�� M�vQ"�����n[߾�Fץp����0������㊲���{��ۗ�����ci�ɺk����0��ӇN�',[b��ά�o��s_]֌S4���3�YU)i�N����_��hϝ^<c>�nQ�*7�J�Q��"Ĳ��8xzp��r��-�Cb����k�9AB���SGN��:t��Wn,�����`���^�F�m�k�im������g�N������I��˟]��r�x���wF��i_+�{�u�_+�}�/n�.F�#�nXH�"*(�ۢ�Y��U)���>+�� ���N�K&�d(5����&�2��D�צ涨�H$�A�<׍�x� �����ٳ$�9�ާS�z+3�q��S�H�v�/�Ҹ�c����&Ǘ�4�snZ�}�U�!7t�\}װ{�=���@ �[c;uM)uXY�L,�+/u<�� ?���@z�� �:O~��M�C�٤9m�tT�W���m�+s�0�/x�8�e��V����o���+ w
Y�P���^O%��dO���qr�Xq��J�^�n"H��2s�.�?Y��̤�!���	���Ԗ��o��X�e�B�i�.*�F�4\��+H^�}�8�\_�؅ε<��h�WI�iŵ�-��ủ|�א�f�(Pvr��C0`�݉P�ec՘jMi����a�鷁���p��9ٖ2�D�8���w�����1�sLY�Bq �
�U�j��:�^���_�6vlul_����0�
;FhD ��$aYP���k|a6ؼ��X`HY��?o)�u�&�<g��
^�hv5�Cr�e��=�ϾY\���[�@���D���n�=p����M;�ݥ].�㗛f�U0e�4ϊ��"Tk ���|Ê�o?b�.� hlb��%��\;s��'��~*���
�]" ���=��~?�*�!�)C���<���)��D�*�WWnWЬr�b�� _�F[���w+l��o�6i�T+�:ߟ&/2�ʪa�ެ��X�bs�7ø�4�oM������w ��:�`/y���#>�ۗ��g�U�\���o���p�}���J��֋5�I�3yGX�v�� �׶.�o���5P���������-Y���Q҈��mУR�d���1̏Kc�2�(ny�lK#d�d��l�c�~[�����r&�M�j��
q? ���{'���$"�͟��
�}�(kX�c�+� l�Lk�U`S���X�����5l�`��D.�>��ԏJ��|�N��Y��ce��gqG$qo(E������Sw`*���_���oT��\��S፲���ڃ[W�T��8� �z�g�))E����O`�����׹*il�k�/g)Lo����5��5�*>�:�����笐4�Xz�O�7����]˫�Z{z,�oH�i��^1�[��IF75��"g�pmaa0�=��xx�\�PyY���[q�JZ�� ����Jk`���Q��(��KH���Bk�L�K�`5��0vn|�$���Q�e�"a����yO���gM50�*�]���^��;���A�� ��^��L��_nt��G�>
\
~��&|s�]/����]������r��?������{���,d5|�v��P��m�f.y޾`�4�N���4��VAU�\г��0�W�{�9悹}�n��ly�H$��
"�$&i�,!p� ˫��#�����V�vV
�*ꇖ���c��9��f���`ޏ��x{v�"���[�[�nT4�b�2�[�a`A@� ��0C�b`����L�G��XYJR�O�j貚�fג�J����@� D4)�XL���h
Б8�? �[��0��|�b��Qa�k�ljw��"�e'��O:�vs;���_1>O����C[F��r��F�ۤX�M0?�C�����q߾�<[&Ks��/��p9A�`r�O�6`p���B�T��Q-$������y�dDŷ-�����ʟ6�:mm9��^�K�E���� �W�3����#����=�N_���N��N����s��m�bxDw�̌��x��@uw6�w<��D�s�y{��߷�2���_���Z�L�{vO���^\�;A#��NC�s�l2z�iM�!��z%���m��ЩyxgS3�v��f�i� �?�Vn7#��Ip�m��q'8�)EA����z]�7�Oiq�QN8{C�����?���<�*Tp���,�7/lY��3ZO��o��twnՈ�/7K��6O[��,��V3o&�{Zy\�z;�O�Eg ��>��T��)�7�ݵ����K��ƽ��P.�^��L@ ̧�p0���(uħ�ؖ kv	k���� 3��c��0g�櫤'�<�����W�0^-��m�(w�<��]���QP�C/"���Wy3uv]������BlR�´?ץF	�տ!�5˔��j}�燨[谽��Ɍ������9q�5�����۹��qEFU�<��'��@���@� Q��rgĽ���	Ṧ��i���:������tke�ء5� ��ت��J���Y���jP�O��� ���O"�	j�7�}����i��+ϢЊlx5p��p� ���tIf�n���5�0^A�<�&{����9�������hk�9ؘc1��+�߷���3��/�	0~�@)�0Y^��Qr��_���9���V�6t���Afgr�/sHkn�~^�ibۍW��:b!#���F-��֐`��~���(�>R��p��O�P����������@<��Uy������@#bc�Q��X��B��m���,P�#����elP�fM�/�٠�֒�z0x2E哘�t��.���kn)�.�N��tj��"��H��nOc��;3��8�ɽ�V��*�pT�9�Lc�W6�]�dͷGn��oB��y���@4&���*�,л|	��E�����1ށr֜V����J7t�)�}��p�� CF:��`J�٨�0��m趦
^X��PR�h���<
 �ܵ)"R����Y�c�/)~G%f~��k��F~�ԓirL꽢�6߮�5VTNV΅ɷF�gܫ��p�dq^�-�/�v�^�io�{̜o��1F�ZG�V��[��u0�+�݆�Y�k��_<�����@�� q8��%ӱ5���$#ۣ��˰��~B��� �vW|�D�
����|���孰�8��+/�{w�+�>	>;�~�.Xò6���kv���C��h��{j-���\;�[�j�����עr�(f^��李���-yX,r�g�\8ؾT7/(w��X-bB�$���+L)�QV|}��/~��Pc�b��X��O=��'�ɀ�� 7��ݍ�	2�9�4E>ΰ�c������(a�����G_�>h�?��x��9h�d>��L3Ԗ�{�L�G6��[_�lUF,]��2�|�
:4k�P���I`D�F��5Uv|���ȯ~�y�+7�-G�%n��ޞ�~�[w�9�����0JY�|��?<%<�G����{��+s"�(�3�o��-\N^#�\"��*����3Os�ĥ0�g�j �7@��70f�Q��LƧ�jjܘ�!r4��oH���#�n(�
�dk`��-@���=�^~2I�f0���Υ앙�0x���N\^OFf��>2����S�?�� ���_��P�[�E�ׇ���֙|���Wr�5�������Z���%������`v����v����[x��x �1���c}�,�_~9Ls�c����AT�`@�B����ԣ�[�'���[S�$�V��J��W�D���{�?�i� �@��΋j���/�R��s��q-"v���J2���7���3.�l��h��,��#+������xy~�&W+��a ��:�A���ɴ4]\f��O����߯��b�S�y�# � RmQ@�G�{&w�+坵�F������ 3�^Ϙ�O=��!�w!�WuW�c��޺���ɚ�۵�@�?=������
{�H��9�G�x����BG�&l�O�T����9_�g)2�{�X��}x@���X�\�M�o�� ׷"k�SL�E��_�.�u>��������1�t���?svft7?�s���3��*�g��?�=�6�gf�B��NU�1��۠�M�>�<��x�Ȑ�Z��&��2�9��h��a��')�A���2��f��wP3]�<���>,Y G�˵� ����/b�P�`T�n��f�<���Q�v���5!�m �Ҝ��y�
50�Ĭ�S����@-�;!�%+�D��ʃ<���g?eO&�r�:�ˌsu�k�_�@v��s
�h�SC6�����!ሣ��h��o﷠�v�kj���GsF�\�U�6��3;w#��{FX��+�iM]��/kа�n4��5acb���F�P| c5��H�j�8@�PDbCh��C����'���ׄƶc"�#��pY}��s��"��j�d��BJ�tiV����������@�0@ a0~����	��EB�	�����"`  0� ��W�ڶ�'p(W�?xQ����J��<gK�1ܭҡ������뿄F@�g�)� e��bt��9���Go+kوb���Gg�����n[%Sy��$Z"�3l��5?0��9�(l��յBQ|�%�hhmk�馡�e�oTr��Dƶ-r@e� �6$[��5k����2�S6x�(I�_�<�Ǥ��V@�_�bnA��A�ĝY��������,'�C�D��e� O�@�
<0���db��`[e��l�`���LB��w� ��-&"CC5�o�;,���?�� 2a�C��׆;6Q��5���'����[�����(X�:F0-`�@"G&o�S�K���y��*�,�w������MG�C!S����D��,y�s@������PCN�3bi�y����;6�x���0Fgg�׾��U�HA�%h�`g��k������>�>�>Ζg��`b�5ޜ�"{����{�\:�/�9|���+ԍ-R*�"�@p"��.�@^�i�7\����r�}��l~	9�y�ִ?c�J�$�_����������&{1}����v*=�t���]�Ee�c3^H�LC��PC`Y�Z��:�A袽LP��2.��v�gS�|+5�V��7��9�+�c�h.�:�u�����-�i��$�:�ϟ���w���o��}-�t�����2~?\.�U}4z)��=��x8�ō�Sw�A4��.����K��r�M������ڳ��o!���	}~���!)-߃׃[+waC�1Pz���ص�f*��p�NIײa16�������r��2���p3շ�b4{�6�T��V��Y�7�i��R����óĴ���\���'�*F�{���M�}�� �P\Ͳ+C�bN��=���8�k�1�2j�����������h
N&^��=��*3���!#�(���0�w�����ڶQ�J�H<�`�����\{Ր~�������=K�M�cY$�|�Ќ�j���}T߽��	����S�>�=I�������cL�<4'E��.�лe���;ƪ�*)��KE��;Nfuׯ��0��m��e�	uc�	+X+��~O�~���#���Er�/�W��,��`[W��l�~7V��-�P.��io��tTAg� `��w�PL+y�dov^����dO�Լ�G`y��#m�*����c��<�7Z��(�i� �B�KS7�d4��� �3�n��N>:����}�b��^�6b*���{��=^'l�N�Q X���V��)��,TeW�˲s�O��+�*ƋN�4Jf��(2�ܷ��n\��%1l�{�� $@�k,g�q�U��;��!����� Z�g=���ܾk������gO^�|K�ĳ�fCa���e��<�%����� q� �,�)�Z�q�ś��f�,�M�k`[;Z�mq.��2��OD���~s�GMIg��	`p=�gu
;h#e��x����@��ߥI
2��^b엒1���b Xެt+�_���o�?�~���S�Ԩ��j�:�b�f]6��y��k�:X��҈/��E��i����/�ZE�bz��C[x]��a��t�PS�&����Y#uq~�C-�C*~c�[�E��N�|?ywPl8�����z}�0�2���4\��c�qW�ߜCN�?cR$dt������m
א����\�>��l-E���k��XFmF��oBn� !�Eж�����&m� X�j��hl�lLϙ���v���[ک��.����lgm��&t�d�ye0���]Cq���E�T\�Aw|�Y���C��rT�a!�&1!㚰'��-_���Wy4��j�%�m_{o�jW�L�C�4k&w7�Yf�̕v�T���.�f7��[���ѹJ�U�jc̏ �=���o:�//�<וnoy�㱹�*��:��q�i�����Ӣ�[A2>���^g{�퟇��hkLS)�n�τٴDMF0�Β�`1<�qE6�|�hi,�?�A��	/|�?S ��+pC<�V%�ϏD�։��8c6�����;CjQ,;؅ε��t%ł�_=��I����2�3�2���`�?$����C��S+� DDo��e�\q�p�RMn/M ��x�ސ�5����{�o�����7�8�L.��^ɦM0�_ �ނϽ�^�0 jK�i��b���]óf�wf�N���Fsȏ�� -v|��B��?g+�9��J�p �����
��k5�3�\މh�V"=�ܧ i�]:\P�������]õ�x�͝N��	�L8��tú���1���wU��F�D�X-x���(�	�l�^8����)���P�uF���WЃ2O,�Ѓn��k������Rp�?U��b���>���"yb	����ݟ@� :%�!2��	����>ݳ�8�r��ľ�H/���b�3ӛUӯ�X�	�Mt2t���G�̡���o�e��2%�����Vl[�ʈt<8x{��'�0:2�y�Eb���z���p�����2���6�0G�U��	�*�e�ams
����!M���ʑhC��n���2ޑ.�܄ƥ�0��g7*��J�a�,�8���l��͠��\�ŋ��K㜟9���V�ړU���\�[��=H�;�(�oPz����1����ط��H�垆�*���ʃ�6�#N��ts������u�ˆ�G��\�ڙgT��֪+�]���Ƨ�N.ev]�RB��Ҵ�]e�o��y�]�����0�=]6-�I�_f�"�d<*����#��|�Sʴ���T���B[{�B��^��n�+�^�j�&��]�0u���.[|gl6K�)>��9K(Vb�����{2t�Ԣ�Z�em�yj����0���\���x/N�(F�˥qSc��>P���̪�9:�el�ك�8b�<��˸�{f�tؕ���*����nu��6P�qK�����5XY{+�tz;��Δ���î�^�c
ʜև�ܑZ�V/��E�ơ(�Z�5�������=��N���]�2,�u�[I�q�8+o�"2V�)�pYƜ��qu���j��t�^1>�Wne��XP��ZS��i,�3�vevBU�;Q����;���T���	�Q�z
��B@� ���_Uu��9f�#��y�T�*;a�G՞�2�^>�E��1�w��}jϨ�dN�l����t4m�wr�K���Q����QB�AT1ؚ�h����.��l���Hb��D�2��t!��/x߻�h�,2���U��L�tC:� ��z���\]�!��!��uk�04A�i5��Tk��pC)�V�pu�݋t*��U��[o�:�$f�ᗗ�t���_�we���"f�ƹ%s�ռEkܕ����W<���
jFf��>/�Sw0�:���q��y�0ʎ�Yg�X��([&�Z�ԋ���=�V���e�����d�@�N���|F�
�9��M��7l�.,w�V�Yy~%T�œ9K����}w�kC/sT�홳#+8�7���Lz�q���T�j�2�*�U$t�|v�elA�J�s#��8
�U�'v%Dr������G���u��4�gEú�����`|����b\V�`ݱ8WD����Ykz��iI+(�(��0�|���l|��b���k�Uf��v�2wQ�X~��h0��3��u�&~}Π��v���vz�ǁt��2򶫪�z���q��
����6������A���g"����j��tަ�zhs
���<�2tl�p�]�ua��H�`�Һ�ox˲���De7syY�7��4���M�噊�(��Xh�c[cLhڶڱ��V�hǊ�ZW��1�x�lm����m�U�&���M*���lmM��񤭶i�m�1�J�c @@0�u$)�,�Z���AF�B%%Q��8`�@X0%���l4a
2�LF� HA"��?�>��z�F��b>�qz��a��J�_Ư����}99^fT[���e�S�I�PW����� ���Ų�0����ӧ�J�g�����$O��wb`Kn\���nS8xp���)�!K�	I���"�0D���=z��P飧O�N�7��{m[�2�d����$�;����ϝw��u�iiL4t�z|:|��a��'�tf^��z�|��1>�-YlX�:xt��Æ�G*�=�y�y�#$��ߝ{��Rի-�l�������>VOU��r�g��_n���.����W����Î-����L�Úb�mZ��۰��^g�YB#$L���������A$���l�,a�m��e-��}mJ��ۮW�q!,l�jbLS�T�x�0�z[�V���v�v�+�G�UX���R�rl�E���[+J�M���+r�7������a&G���Z���"@@ ��ǻϞx`PA�Z �����&��X����`�ɐ�xsȂǯ��b��E6�ƹ|��P׌;��#�*��d3��XBN.����+����BY�h-~��*����oBaS��4��Rͮ�$Ӿ�ּ=4؁ɶ�&m�_�a�S�j�$���@٨�[�X��M����%ڙG\ \����Ɵ[J��ᬄ�]t�_�T�����sg�|�J\"LQ���*k^��oH�<lE��/ �c$:6۔��s���<����!?0Q��R�Kc�%�0Q�]1r̉��t�xU�%E!�lO�A�?���ӳ_�q_:�P�Q�띵W-�`6�>{�
=	yNZ�E83�&Qҷ�?�}�?�xc��O���������U��[�f�ь�/k�``fHf�!�{nl/"ޖ���ͯ��:=Eg�Qkf�_�VT���UP� �m�V�w���*�~hwU��#��M���غ�^�ؑ�F��c�j����̠���h Aܗ�ǦCx'�X��fEkhߪ���S*�a�ad{�<FooĒ�<�>���bU/���]�u5Yz#}��T�g���x�lř�T�i0eQ1��|D���S�i����Ng����Wb3#ƪnv]3;x:Z�LJ����]ާn��9κ�B��)�ASw�g4��D 4Vި3�'�bf��Z�F����o� ��*�`>�������Q��͑;�}��l�-��3m�8����xzn+���v�� �^G���|���]/�P��"������xO����z�L���&��O,;�ϟ:��mb��3\�MӴ �,�_����*6_�bo�ڿ`Mb��Y=�[�CKԸДSH�!��º%����Xy�[����}�{�
�3��fr�~G��E��Bh��ƱҽJ�/\����=�Ƴ��@�@b��0=-�T�=��z����1Ml�B�X����Q ��^h^�/�$����`�������iBbl-�lRɶ�9\���l0� 0{�,������f���	G3E)��5��.�b)?��*�5���nE����+yI���ȃ��UF��,�ض�����o��f�_<y�ؑ��[v�L@�ź��^P�r!�4�!�� 1��
�LUd�/i�5�F�к�ɫ�O'S�G��{?N��0w>��Ǐ;���,�xMl�s�#y.V^��/��2s�36¿*��bY����Լ���H!Ӕ^;���k��jd�5��9)S���N%��)�M֤��I9�xz��B����i1�w��.N�����	� �� ; j�K���o��~yp�o����Ҳ������/���Y�'��8��v�Ƈ�"��N�y6ۮ�=��L�K�4�O�<G�=%�<���Y���!�9`+ �E��2�X�s����C�oSj&Rq�vE�v�s��[����Z<��q�}.�"�b�Ѹ��O�L�$&;B}y>1�##:���ӕ 5{\���s0k��X��~�f�>x��$M����wP9��R��h`��C�DC
�ڴ4���%��2e�2��6�ڞ���PS�1	A`0r�Ν���ֳ1oVO��7���/WŖ�`rza��_���&�r$�h�'��	�.�h͗ż�2����6��D�sШ�e���p[�!^��s�ـ�F�~��N(����}�絆o����F*J缿V�1^ۍ�"��{�,�A��1Q@:����wu׉(��{��n�,�b-�WAeD�
��Xo0o6F]1~�v�2��W�a�^T�
�M�G��g�K��_b�4��c5�"ڙ6[�"��;#J3�����׶S���jv#y�F���@��{�{�@��ə7��\����b�z�nyrkP��?{7�XWZ'�O�/
;�{V|5�)غT;������2�t��W�.s%�yG�zuR�y��1�5rUz�����~{�댟��~S)+wfJϷ>1�bQ*��un$[�4L\L�1������G)�	v�F�Ӏ�Uɗ�3͝�M�����{"� �C��/��T:m��th*����LS.~�T��tm�O���-Vn5�R`X��y�!;M���?{�ks#����g�0�m��&��!��0͘-����s=pw��Ӫ)�ֵ�e6�*V8�
9��66�a�g���G;��_q�=�z��;.�;i<���1>�[���%��@.�yx	�x����C�ˀr!����'Pb�.�Jj�3N�E����M�b�+�T'|0f�oQN/6
�"�y ��zb���b:�]���O��36��P�ܩ�@�]���F��/	��|.���sz���mѧ"�<��cN��3�/�%�7a8ӪG4܈��s����(sl/�"�"5�}B��_�~������N/�Y}g�p06,�s&��C�Ů�/�_ !��=��ͥ����`W�[�7��q���g�_�	"��7�}H�����zܼKw��W��e��u���212�u�`������g��1��X�!v��?�r2����aUF���n���ܶ���}Y��.bN�UvP�ܲQ�B�V�r��y�rz��=쪉���
�3�7?2DA!�����I(���k����WO��k�m�.R�[�����T�k�L]��f�oX��8�3grX)��f��]?p���A0 USm���XcM�eo5�mb�{�4���]je�/��ZZU/��@�`�|�U�}]�/���+�驟�K��|'���"=Ҋ���j�l���l"i�-��X~����Ɩ:�Z����w�\�9�$d����?(;��F���\9?�\�3=��_B��i������	�P�Ͳ�T��0x����{����v��瞒�۳���޼�=�y�>�f]R�����런���^g��=�v}�]Ю����'����[E�R��b&�J�@���ƺ��c���9��MS��/;���{;��%[R���ψc�n兲���U� '�����CQ��秅�:�^Yݝ��p.5�9R[/�d�}�ɶU�K�׭����CSd�7�K�E����ȕ��=l�ͪ@h^ޞ�����)>�OͩA��^�����aݱ�l�q7�ξ*�^'}��0XB�4�7�k���«ד�m�DȎQ���krcq֨Ʊ�e��t�#/o��jO����� Ű�H�ꛤfM���[<��j��[}���`_ Ş���񒰷���ʑ�~�Θ�����7ݢQ���v����8#�h�m^&�*C.�d�/�ˑF�&lm�����,�&AR=��(�g�n�-��j�Tr��*�tU��S�7y�!���C��J�3KKK)w{�y����!3�>b�ag�G�~�/���Δk��[�\�]�q��utb�V�����Z�ʆ�C;Y��8N����_S�����;n����Y�Y��K���#��/l��oFO��	��v���a�i��Y�ђੵ�/�Pt:mi�����;KN��Y��F�A2q��E���An͡��^+u����v�2L2򽛐2CG�~8����C�ɪU�i�:Z��T��><T����=�{>�X~�v{�:��h�y����7�aM"ӑa�\������.�t[�� �E#����LLS���1�����5# j��a���'L3<r�̞��	�l&����ffB�MR��m=!;op���P��-�ʗv��ho���a���~[t4&9�]��巶y��Z�ւY^�|v�V)�xi��$C�\����&��&���ӫM��{s�F������t3&��6��@jl�T�=�Ju���v4{}&�_TCs���)�⻂�u3���L]t����O(3W��S���xߵ�Fj�2e����C��ʫf��n��� S��\����n��}��D��j@����U�47s;j�'UHݷc�!Њ<�����5u����3[�Y�e-�)�p@o6.Y�������p5�@q;��‹S�u�%	������l5�TE� |>�g�)�����8�y֥�f�}f��̒�kkF8�O�����uf�m�܋cS���Rē{�Z#~/�4�<����B���SÃuB�L[ͷ�EE�S͵gܐ�jH��@�t��yҥ��4)&Ց�m����E��c�|�;\��ys��^/��=wAZ\��ޮt��nv����������\���ւ�VC�����{�I3UXΦw��B�^����/�	AAb^���{��`5����i��'P�?D��>G.��y����N�q\[��8�*�H���;`�+�:�V��I�Cȃ����?�o�*����x<���_"�>ᢆ��x�6ޟ#^�CZC���i�oF�+�O�Ϛ�B�"w�TJG������}2��>y�����Ht�@�f��G�a�l�~/7[��ށiBj.I�-�)�����{hʖyt5��z�6?�/>��!yl��X�W��6��|x�w촘.�="��ߋ��5�-ؤf/��fާl��7Pn1ìɒ8�y����j\PՕ���'QUrĆ@��$>Z��Y^\0:YV�ǁNݾk�/���O�J�3��l��[3�;۵'j�ewb23&��Wv;�����+3kk��dx���~ ���0�5)�p��S]׼���������7A�y�p*���y�Gd�pK�+�-�>y�fZl�6茙�ٔ��ȫMR�4_V�������k<��t���Ѭ^��`��Jn�lPu)�ӑ�<��a�;/Ld��80����![8�4��e4`�&�M�a-�>�ڀu4vf�]��ً��o�o�Ǜ��Z2֮{.��05�KxH�-���\���T�8��.�H͗nK_����0z�j�C,�R��{c�ė,�= T�sS�w%��>(���K/(-����3�~����8��o/$(Ǒ���B��6��9n܀CEfZ�_6c��>L��W>Fh�h�X�p&�f&Y��Yߜ�w��/i�#@�d������k�t�d�|��\R�DKt��o׷|��*�m�d����JwR�1���Uj�/�?�����Z������Y�n���w[�z4�9�q Ҝa���W;�>@gҎ��婳���:H8z�B�[a4Mu�s��啚���*��Q� U���c����O��\Z1����c�����~�`�}I[9��׬��T�P_KJH��̺�㣼:�P|1v��V�bl���[<x�umH��<U.�$[�Z�"�����(Z"(�
����#p%�L6�Ŋ����sg7�ջ�W��p��v�lL����c�"V�9Wi6�F0tknX��� G�)�MLj����[s<�{�?B�˃3@��@����<~�W�B��(F���7�1��Lŧ�/�S����R,��9@z�hkO�,�e͢�6�������y�Ŗ��??���^���G�0�N��>��ţ7�X��[�^��Z6�3��8%����{m�W����C��>��4D�����Sb� ,G�w��j�s����@33F��P	�:�R��Z���c}��B�t�^�^�צR�{�����pGY3/k�}jw-����a�¼����Re�����F�J�g�L��断e0v������?f@�w��`�^`o2{����]*
�h�'�����ݖ�~�;�Q؋d��	�Z��q�SQM�'-0���z�r1�we0X��ZD���ç�u���g5��헝�'��K4D4ǘ�.�P���ї��Pē6��xb�ݍ���LV^F�� h��`���n�j�>�A,�T��!�=�	�V@�g�=~ɒ�3^�P[w��u�j��f�;�q-�迄���`Ryb8m~�.��������:_L�\,I��&7�bȿ9�>��"�Z��&����ȥW�n��囇CJ���W�`�e bzŋ*<��_cɡ=��W-�2QBw6T1q�A=2�����C���.�T�\��w6������wrz~�,�J30�pp"<�Uy��Ṿ�x|9�=0�7Z�Ц�$+�l=�.XSN��IP<@l�}�0�v(�qioLu��)���#�4����r�.��>�����	J�9�R��m��,�a�Y���N'ކR��!�`f���vX)O7�e�B+��r�Sni'��s�|ۚ��Kg3T̽�$_ �}ex��6�w���o�3@R��-�*
~nY�S����ʞ;�D���f+`hh0h�j0`����L����Δhg��-�rp9��j3���\�%��b���.�m�O�Dޱ����}�ȹ ��|�=c�|�|����kF��(X#BA��o�|1��j~��/�uW����|��H�k��#�s @|s˥b�l-�U��Y�ػK���p0���'�퐌0��� �4��W�m0��&N���J�fm��ߙ�q�؄K�!.4��͟f0'��d���	����^��r�xcMmlf�"�]v5*�Zм�X��8�<=�7�}���c l�>�}��C�@����s����]ݝP�Ǭ�F���7��EJ�}���Ԇ���L��z*��3,ꌵ�]wY�M;u����ʜ^KcV�_�=��]�-��Kal;��'���/9�]A\�a6��Vѧ0AZK
>�-e����*f�(�=K+�m��c֘gq�S&��)� ��6>��MN�p'8��՗]�sh��JR���lRs���V9��f��]��6���;��'/�q%�F��Ӹݽ�O]���G�<R�L�'Ys���3=Y�>��E��33��o
ԦW�J��l�"�i'v���I�.�W.�P�k��yzFp����	�ۭk�uaW��o�w:��n�^��d�Y���Nn�Kr�Vٱ��-=�duaL�:5��\tij��J�uks�2m�2�:�C����[u�B�\��N�e��P$��]n�����w:�����9�C\���3���5/r^dꝡLg.��9���o&"�&Tzw��{��_��ni��ZR^���@se��M��RUs+��قRD�uN't�泞s��ot[J����x�C:��ٮ;ҏ^�[�z����I����(�:@sMj��k�+��[Ž.��Vf%��Ox+�t�R�P.�ʛE$�<(H$������hv�wdí�[��a�4)���v�袨�T���s����Zyч���1��S+!hSϠzl5:���$�+����k�4�en��z�W��L�6߆{J�,�]�e
��Ba��2�V
]y���AA��䇆��z�
"�c@cTP;g����{�T��γ�Pf:ܙ��c���.�ۋ6��U���]Uz�a�>����VƓUv�Ե���ל�s�Pu���9˓���Xj���y��)�e�Ո��T�f�tܬU�,�9Ԏ�9���B�4�-�Ȼ�D�B�@��i�r���b�w����"��s�v�E�Յj7}����o/b{�eH�n��N*�%A�.�sGf�g�^q!,���-[���&):��=}Yu��[8�si�^�)A@鮾����g�Z �4XO����R��t.��N�3�<��b�(t���;ݝ�e�]$N��:ZqLI/<Gk���vqx/:���'3yKg��`���|�ŷ��sR���j��+{!qȄ�������qUϖ��~]\CPa�W|к�]ێs1��A�t�w���ɢ�m���+�!R_Y��􎀲�oL�Y�4"�'{;w��2gRݦ��7��L��0J29�(�]ݭ���Ua�5�mc������v�S�1!�6i|����q�y�1g+�����]����[�Y���������s������,�7c�n#�}Y��y7U,GM'J�01�� ��E<o%~A�A$��Uo9/����ۙ�#�nIH�y^����ç9UmZ�eZ�2�-�1�Di��r�]�dH�ܙjϔa鳧�O�Oxr�}k;;�A%4��W	H��Χ�h�]^W��_+�|����k��pC�!��7��c�+��w�^��l�ӧNNYl���m�-JU���e��*S��8p��|
<sFbE}wf\܈��t�[㑥y^W��_'Ç�խ�U����^f[��&"|u����Wi_U�=>�:}9]�-�����2���^�ǔ���4}7<i�>>9j�ն��lc"2D�}����ۤ_�~y�}�����]xԚ Z�_,2�d����Wy�u��3�������L;_�J���;n`й<�����}ɴk��ɕ�����h% ��_b�8�������o���8�����?�~�GA0}�����B\��>FP�O�x��F�_�_�J��_~#{)[��|bW�Y>��_�Ȧ��^V\�&�yRY��Q�\��ֵ�����F�5,�T��xj)tK����!ߥ�'	��j7������d���sz/,1T(V1�8��|�c;U��������,��3�fե�NA080�4�z������)A�����Jr��/)e[m�s����Duw��ʨ/0�{H��0��O��f���j�Uk_�r�״H3���N'��jXr�mr:(����w��s
P�^��y�!?WόP:g�?��WtFﾃaֿP�$�V�u:j�,F![R��b��⚘��X������T)x�+�Hkͨ��
�F����v���X�i���9��3��Sg>;��� �o?�K�t^[���5\$3�����kG0�w~����w٠u!>���Os�L�`��d�rȻ=i���w��lZ���qN��]��edk$�B6���}��P%:��=ob��Jpͭ"�'u�&L�ƅ 4>�u�?1�l[������\fez"%�]	��J��e����wk�N��==�
��du��-�RƵ��m�μ�����HB�$ �0�0I���v��l?�����{ù���q������1����B�k6ŭ�6�vk�}�J_$+i֚���]�̄����U@uo�p�F*��>����@���}`v��&9�vM�O¥,ϞzM����yĆ8`�	���~&�q}�Ya��H��[&�A@�W1�
 w��c��7*x;�D�*�Q�^|�g��k˽�x؉�Fz	�a}_�W��`�B�T�����Z��N��ٽϒ�ϸ����36� �ʮ���a�1��fG��'e'�K�8��p�*ܧ��ٙ��[]����1b��V�˜;^�p�$ͻ����!���Lo���~�ð�sL蓖��l�������ӎ�l=s�����[cik>�ڝM�A�p
�?h�
_0����ܭ�ޛ��/���j��}�
5�KS&�|�`"������V���v�u�L
ؚ6۳z���	�[�Omp���ZoAf��nm~�c# �ϲ��r���X�$p2jw^��������uo��tFH��εz7�ȸ5�@f�T�>��{�0^�y���]��mֱfm���B����;�߲���g�Lͫ4�o�(��~�/��<7�ɕo#�Z�����GΨ�M��ـ�ۦ)^0]E�V������탷�� y�2;z2k0WR��R���ΣqU�a���cݕt��]���B����`��0� �@��H���l�.�v����Kai�����o���kP�@����f�+[�����_z�u�������!5O�Yb/��_Cz	�@�d8ӊ{-��gmA����Y�6`�k�EJez�S�9JoT(��e��|��pb^��l�ԭ�R���ϵ���SO=p+�y��S�(q��H�s����]�ن3Hg��@��w�͚{����<'��o�^�/�����8M
�Ry��)�~`/��3��a#F�ܱfb���=�5�/�d��Cb��sϒ���9�x��e��8��aW���!}��v�^���	���>�+7K�
���b��C۞Ŧ=�o6B�T�qZ���![9�������J�zr���"A��ͅ���kQh����D~$IXE����:��褯����? � ��<��#Ǥ��&Y�Y�����G�t���@m��OSw�=62�yHSv�[ѯ|}��X"��Ә��~x��V�jϖV���ޖA��+�+˚Z�;�d���;�J9滫
j����\y/[Jy�w�)��b�3����o0�*�����TDX��.����Ǘ�t�}�ޓs�4o���j]l�ɮ�H��m#qݣ;;&��y'��MO�=d
g3ۗU�Y����T���Ⱥ3�bLg���U'W���ռKkq��7����Y�^nt��л,����������_}����߿y�[ZDZ�j�4���Y^�$hP�0,W"m�խ")�����T_4wWvg�X��A+<��ѰІ�1ޗ?qs�(��Y5��]p��i����>������� �otiƮ�	Z]b�,�`Ѳ�5�+�>v��q����>�Q���<h
U*�&��T�K���LS߻T�
���� p��Wƚ�v"lg���B_"�7j柱pu��^9�C�K��Swf��nZg��l��05��ڼ�G�f�8}��9���0уƃ�]t�?C�O8��8�I����J�-r`;@=��>�זJ�»�]�����0�B��gߝ�h�����)O7���ЎQ���#X�06�'�֘l���#_+&��k�Q�uKl
�:dOL&3U�2�+�B��u��V�
�i�ԗ(y�{F�:a��KEHL@�1���`\����*N_�1�M5b��,��݇"\��F�WD�����u�_����~� �z��ŀ8	��R�!��^E�'̇)�pK*�i*q]�0����;�O]��:��o)c������{6��l��;�?,�z�\a_������EJ���t�&cٮ����:�`Co���y����+o��=��ы��auUw���o{���~��ab�d�
YJ�s�*fs�!^��������>��p�ٞ����W
.�Q-{�G޿�˩��U�Ti��ќ���/�匌�F�B�	w�`����Ł��,�I�~��s��������.��G�U8��T[3Z���j��epZ3ZG��=~�r��:;GEn�n��͏:�|>I��_�6'���g��������	�>Fn.�%��Rb�&�4�ںO����;�?=�u��O�#ȝ�O�5j��,�Y��O�R�m����C@x�x�6i7��.�Y�d�'��"=�I�1*���l�?������D~�������}xVҢ���^���P�� �� <72�v�����W�M��_��`K���\x�}l��0����Z9�,�̸��ȑ�&��^΁������q���^�����$��{��� �ٰ쪚=Zdq��o::��h�Sў�X�>2��&߃D������q[&N���&�	����*l`�ن�r��~�����W2���p��,��=k����j�`��՝!�)�k�����U�H����)ع�!��`��� �b���_Ĉ���ь7�㒬6�����S���9�v�ճ�vQͿ���אH�(�0,�����.��jֱܬ̵ǳ�nj.�w*�B ^d�9Ƿ�6zFj�c.�z�p�u�k[�����3
����������S�F����b���'��p!�����v�P2cꫲ&?�@�[݄�UTs�8a����M�+��1�D>0Ɵ=���x\�%�q�ς�	o��={��Nr����J@0p�B	�X�bĔi׶�X���+<ϽЊl�tc�v������@ދ�_@F/[f##ע�-K�XʕȪd����;>��Fl_���/�O�ܴ��ս��r�j.sg�����\i�ƀ%FD�C\�^���z��D�Ƒ�<)�Q�p��S���qx�˵�j�����7���b�֯;��9��X�c����2;o����w!v���q�2��z:B�u�vc��!�,ݻޯ���_����b��JӒ�q��	��l{��fl�VAC����¾^�c� �zY���|�7��P���Է5)�	_LwAn8\�Iy��O�P��\^�)�$�OΖH x��fZ@�7f��S��Ǧ}k�4��
�)v����ނFl�����<ٛw�S�G��M"ιj��>�����y���3vl?�
�r�w�y�߇׼$v�uAnJ!A�jXejC�Cf'�pfD�|-��l�t��@U���b]�M�u��p�k=���Л�5-��k�����f��
ܢ���0�瘂0��(@��Ma���]��k˯<�[��Т��"�_����mw}�=�C@�	5���,�m���F�Gp>�����t+,oդQ��#k�Z�J(�\lu�嵻��xR��έ��`MЋ�8�@ׁ�k���j⋛Ô4��qR�wm���r9�i�U���לoM��K�Ś�5�9���A/��|Q.������F2&P�u��w 2�_]�:���?�c��VG�&��R��/NOErnW�����)�
�t��v־�2�׀T��0�Ψ�� C.r)���mBX� f�n���{�u[+��C��})��U �P�	����?¹PHs��_7�g��Q��w�o����#�
q�ґ6������gƾ`f�q�g�
�ScQr���;ˆA�#)��쬠TD[�w)�G��hЪ�<\W� �)��ZQ�,��nҖ�yR�Uq�f�CF����Θ3@u�J/0�^w�$��� %B����*\m�����/�{���ת���4q��)�,/d
~:�"T?����>8�x`X��=�8~��Z��J�Qq_ْ��{5/_�_痶��ڿT�A�UIHW��3F�u�s�8�";{uGs#у�{����קZ��צe��g��w:��)�s^�]Х��юݬ�������E�ˢ�^k,NT=v?<�g� �8���Nw"���>�TΞ�=��_8f��J������Y������÷4����!bP�3�O��;80) �l�Y�[��u��k�W��e^�p��|�C�T��|���@o*Ma��q���`秵�ͦ�}^���w��{��1�7^�E�=�x������|���=�@��C��^��i��P�0�vA��6�P�1C7o��&9�=�����Mfe[���ޢ���µ�o7��ȜEU�-�h��q�z7V����U�_U��r8(X��i6D��ɳkh�U�����C�*�]۞�	U�g.F�إ5v����c��4�V���n�%x򱽯�E�1Y����ӗ֭�H��J�r�����v�6j_ú����P�6�n�fq>��n}��v��6�C��fJ��i�c�Hy��g.�I^Ҕl�ny��(9���F�a]�P��Z��-|�k*�`���g���N�_GBp�IDm�Z�X2��E*���W�G�F���믎��"[r�˫��	d���^��ƭ�Q��mNͼ� ��E����w����ES�i�-3Xi����º�����K��):�0s���"�;�n�aZ����ݻ�Z�Mغ��Ǆ�Q��[�݆�-z����c`T)��7�P���}[qY������ע9���F�}�Q����88z��>�[�0�P�Z�y��k�wcW�K���q��3ry��P�Ya��/��!�f��\bN"�$��x������`G�o�1��?��R>��v�Δʩ��4�U,ӽ,�D�@a�Z6F^Cr���XfXtS�s#a����w».�~ڑš��L�K�	$��� g�6�{5��ҹc��Vˇ��9�oT�9�kR��0#�ކ���"�ef#�@{*�jvj��T3t1ȼ���/aJm�6Y_�b����S�bn�T�Z��f�L��&.�O�(1�����f� �l�KY�	xhL��� �Ur���YuS�4�x*U:MꌫRc�'V3;�~�ޣ�ǐ�U���a��-�F�#��ɂ�vh��EF��/�:��0�Q
�����o7�8�34�|�4�2=vf�=����Z���l��qfх�2��)e������ �@� G��3 �+��N`����f�了I�e9S���#-wkaٓm>��h�đk�Յ��Q�a9X���;#��w`,hm�y���9��� @H}���z� �Sa��ﷳ�=���\Y�݂r��ND�4+����iX�M�&��oTt[t�DM�V�b6�HZ0V��K1q<enԵS��|��3�hɲ��� ��ڍ�^����B�~ҡEw5!�3�˹;�����eN���'���t��7g$�]�"���9�H��E��w]vFp�#��lw2~u(o#�U�R��nZ-
��ga��Փ䫨�h��sZ�M=Od�)/Gg��qO��Ϛ����;������r�at�P�Oo��fmo�3�%��TT7��Yp��l���q���ʊ��6P��$uǯB0)�u42P�WP�'��t	�;݇=�{���D�<�]�����8/�֕1���\�^Y�J�C8V1Mg)*�-�ʑP�zX��!��3[������-���5)�m�t-t:�(�b�lc��)�u���\*�_k�j>�34�;3&�u�^��$;渮W���k��ǯ��o^�U��e2�u��Sۣ�ؗ'p̢"�j�њ3��SD��Wv{k7��5�6oD�\�Ib��i�Uqm��Ӛ^[ܭ̡�G{����e�q�`���,\k�]|11�3}FU�KT�P����g�Ųl�I]y:2��9�N�u	eg	r��L�����S/qˋ���c��]G\���n�os"��sq�)���x-��2^v.��#��\�l��;__4�fQ�/��`}}&�}Kv��zL��腮F��������}��ݦ�̦�l�����G��rl.��Nv��P�g&ҵj0̌t5��)��"�*�.��jRcy��+{�Jri�D���v1�mc��P�0*�t���= ���U��V�7�s����f��0�ii��9��H�H`�B�Tbu�Q����o�d��͕|�N�p���iwMn�C�٨m�܌���=�E���^��hRd�e"�t#��6��[�p��_p����6귓x;�*��v;��1��Ԡ����^�V����5���1��b?p"�����������0��W縑昄�E�7���%��f�
�Sb���~Ig��K� t @8L�<���/�09a��c|0*���9R8
����zb��2RG�Wĸ�}7�eblɎ��B4K���nlN�>Iud��Y����wL�K�Z���P�qͷ�v@�M�N�����L&9g	(���Eb��0�y�o���7���Y�᦮�cۙ��]z\��m�HNtԦ��|N@�'�G���D��X�3����]Gy.�kj���NV�p\����8�4����7�/:�ks-fӡ��ʓ;��	Җ�1FZ��敔j�.�7�t�T��8�k���&omx�{sJu++�4��텵��X���n󦠘�pņ-x���f���+�ju����=>ġ�iU{'�v����o5ba�y��6\Ktt2��}�qq��Y���s+E�[�5�e�<�l��5"��x2ԓ�s�l�ܧ�S�l"����uT�6b���ܬ}&��9��k��t�o�F���0w��ꄍ˭V�7[I��vWl�y*9���=�ay��V(��ʭ�|닖�2/a����y��j�j��G9���◹\���r�K��u>2����v�0�<���+q�x��Z��L�X��\8�^<6���{�ign3�I���)b��j��g��[m\z�
i�6���cx�LR�X�m6�co�g��1���[i�m�cg�16�m�xc�4±��b����xcliⱰX�!Q�$?��b&���PK [�E[i�Q�\ �i��BE��?(�	�i���g�e����$���יJ�x�#I�����s�nH�� �h���z|>�咭��R�e�!Ə��"�1Z(�9�uy_+�|���|��]-~9%�Kt�o7���z�)���R��;r�<6l��ӧX՞֮Ƃ�IPPZ+���kaN�<:t�ӌ�T�ZW2p��!F@�QW2b�-Z�Kg,e�l�Ç����|����nky݋�l�7^�ݑ�Ŵ��űL4t�t�ӑ�-z��Y-�m�������#x�����Qa�N�����Jxzzt�çYl[���D_��L���6��L�l�jv5�iM�M��O�H�K�2�)24�O�U�T���9�ƯZ[�
�^.��ux)*(�C��d��m��?_}��y�~~�zz$�D���1Rϳ���5!��V˾@��Y�Gl�ٰc����8�Q�狹J�ߩ�B��&թ;]�	T���l�֍+G�4�z]6���{��x�Z���~R�.fj�H��~W�/�Ϫ�h1�Q������b�@m�Ezs�y���
�෴HӚ�M[��:�1�pN�&"/����ܥ�;bl�v�~����}eV@�Ƕ�%��MUScpws��H���8B4�4v�[L�l5�ee�j���D�]�Ñ��ZZ�9��L�����>	�Yo��GH�3�{4C�M`�^Hs�{�R�j�DN��<�c����F�uS ����w��GӉ�UC9l?{f�'��h��є�Q{�1��e4�n�>�W����=�{$٫�G�X����b�m?_OEV]��m��f�`W)	��.4#�]B��6��L�ݮ�.�K@��ӫ���1긧�s�u���[��y�n~��z{�o ��68&� �����z�F�`�<���.���CɁ�Nu�+�Y��5q#�`��C u�m�7xy��=M�ש�-��N76�1��L��Ub�������~x��|�:�j:�N��*q����n�V�=
�b�7W]E��N!9o�ݛm_J͹�tA�$��cA�O{.UΙԦ$����+{��6�����QТ�؎U�k����b&�2ۘ�Vm�(l��6��T��@|<A C���}\~�ە�J��eb��R5=��l��,�ڲ�eviʥ��C1��s\!�{�L����S�;�/���L���t#�]n�	���9���&r7��}P# �/}S����sY�l^.*q-ޢ&������P>�l��Zb.6�@�8���f�/2#��;�ހ�����1�K��������6��8i�U�Ŕ;��]uw�Jz¬1���pH$�c�C;Qm�îz��GC�˖�Z�f��`��2�.�_���a�z��Tk��^���Q�i�u1�m�e�r؎�myx�cu4�y�Q�Ϣl�\u	���7��":x���va�帰���ё��闆CYA�Ľq�� Uh)b=�,��M�+���W�� �U��ϸ���-��7�d�^�7�b��<�N2�4�%�W��g��Ԩ�f[���K�yF<�ȓ��/1�C�U�'�e{j��6�ɝ�����Lz��u�����3�la�`�v��Njh�j7{0��T}�ՇI��^g���n����Yp<�� ;u���X��!��z�6���Kw ������b��j���X^*�����h���/їdc�=@Y|���$���[ղ�ff����7sT΃9FK��Q�U�mH
���U.������~1ʣ���!���Wݴ
��N�n��H`���)R��e%}Zl]�P��w�X^hj�9��LP#AM�l��n;�.����������y�-2_�6A��$�� ]�{���3���0P�k�/�"!oP��Rz�Z^e-:��s��q�+:�q�Rs�����@C�e�[�3�5VF[��1�`�s��ԟn�[l7�����p�p7 �.��;�W���`�kG�cj�3��FL�_~�mW~aȘ�u�����"�hI�	o8���D���[C55g%� Y�!WM�����ܯ)�Ն������ƪ��y5hX��z�����j�`�ۿ�[�GDfW2�mH�^��9�l�>۹u��֜*\ǧ�y�0�1�@�`��J�nM����JR����#V^5{�+�����wv(��N�h5��%�﫚�!n��!�B�^ x�k������o�<(ylTS��'+}�@>̃B���sp�Ũ��Xl�|�Rj0T7�d6)x�k�r�7ʲI��$�e���ǫv�'}6<EK��Hp��n�Q�c5ڍ��"ndUH�i�~p�ӧ��v�8 D��!H�>�ld�g��=.�ޜ1R���U�\d�]1��t�W�D�٩{�Dj��$�j�'),��V8�S(�z�T��N�&�������m��ޠ-�ʍ~�	�riLN,�}k2d%m��껶8z�Q��,�Y��*9@�Uŭ�roK��r�e3�n��"��\n���(�a���{�����A����qZ�h�Y9���^�%^�ʼ�ľ^U�����
ԢF�z�n�yxY�Lpٟ(Q]�u-��t��y=�V�=� �W��*�C�:F��u�#�)�t�]�Ɣ넎��t)��Z5��ŵo��j��6�4���L���h��ΩWŖZg!VWf^:�&
�ǮSq2�D ֪�A�0\�|%��?�;u$;��}#u�6�5�ͪתnT�j̝�}'9�q�g����J��x�¯���,���f4�F4�6�M6�+sZ�wY�����[��?FQ��������y�Tژ8`��L~Wi�S %^㶈�o�� 
lH��ٛӖY�Bd�Vi��be�`�;��zp꽼�`0�n��!�gw��Q�hNJ��]g���f���WK3kM��p|��<wқNe���xQ�L`��-A�{a�vk�m���z�;y�dڠ8�2���ތ[�܌22*�5�oH���fLb�5�9�`Yw��e��*�3�Պ�۱π����h���w�p��	��`�iba�7/�6���z#�=�Sb��m��a(,����@���0HF@]��3������W�u��)m�=�=g�8���,��-CM��8zݳ��s���V�N[4v�E�h�Å! �A!~?{�2�[5`;�UO�� �|�o�uOPŊ���<_41�Vr�r�-����w��Xu5>%h���׊�u����g<�m�K�Y,�N�&�8�^��V4+-�굼�Yg�+�j�Gg��ù�G[E���j�d�n�O��@H(�_��#�m�[�z{�:c�\9����ױs���i�5j�Z+�&�ca������\��'p���_�xy =� Xi}��{�����uC3���ݱ�����_x:�����/���<�ѹ�I�#+d��o�غD	�h�Vl��q"���p.��K��E65N�ѽ�mٜ�&B���c�����of��W1��C �a���Z��j���Fje�.q�w4g�d���˳�J�B�m��x0����ʝ\�;���ˢ��A�a<Ξ̞�J�^��@�1�x���7i�=�Gyd���ɚb�ܣD�P�B�BN����Օ=��ŢW�ij#$�ou�Ƌ'��18�!��h�^�4�v�c>x`5;���`95�S��8��ĺz&�<3|A��q�5������Z@mF`m���o5�&n�%��
��OZ��g�>Sd��*�$�3����þq�)����y�g���_pnT;�^?�H�`2�۠�L �m?��[�/O߿9Q��>EБ��!U�Ov�gs_�t���޺���Auәxi���Oj9���Z���rW_eT�H=�}l:���������bh�PM����k���{�^_C�m����� �5�J�잫~� q_Xz�/:lՑ�;�Lc[э�T'� {�@t�9��Cd��s���@^���ÖXb����Eĉ�;�JچM1�i2Э^�������fOj�|⩫K�.xT1�隑��^�w�K�0@u�ٺ�L=̅�*��^�����$���l.��4.6�[t�w��;q�oc�}����p�H|���*�4��Ԣ�{�8�ޞq��ws�\��gu��a;�Pϭ*ݔ�J7���Z�͔��ʾɼg�9���ѾPR���~/��XJ�烇�a���<��^:���� a�Y�����1��t`��w�1�n�zkV��w���5q��s�\��h� ġn'Vk�Ni ��h��Q��\���^��D�'=NZ��S�wWO��٦�ј�������o#9Y���qy���ە���Yݔ�'y^׉g����t��7��G��}�S��ˬ�pNL��u��m����f��F�K+�;+g)�e����j<R5u����aT>A����c��y̸���q�q�z��Y�{�����m���lX��{'�=.:ʖ��H���S���O�����ò����`����1;�ÒJ�S{yN#��[�Mq�4C-e��˒f���5v�G���!Gu��5./�3�{�+�<���+@�u�g [���N�H9u2AW�����G��vt�( �	�A�"$�,���g�0�}o[h����oP��)&FG:�y�&�,ٰ��(��@8g�iM�a�����`wi�@�-5+��([Z-��:X�S�Dd5�@~����`� ��q��[�詩ʢ�1P��[0ێ�Px�@{�* x�T/z.ٝ%n�ü49�Ν{C,�p�
o���=�� �{���<>�V^5:�/��p2����]L�8��@�Ƿ��%��i�M3�KHi�ةdً�����5����J�r�$i� �K8��g� 87��ޚ'l�-�dȳN��M��+h�ؔadI�n�*,��X�49d^n�� �a:����J���i�W�tҳpq��}y��j�U��d�'�|��1b��&�<�s8�'NMY�s��^Ȋ_V�S�
��w!�\�\!V
:V���N�.�G]�׶9LG����]��,����wJv(|�}��[���84d�;�Z��K���@�X#����[֦�˭k&~�����`+cWr1K���.#� d�	��
�`�ͷK��hM����G($��k��k4����7'�ii��F��®\��$V��	ds�X��ˀ�ɭ|5<oί){�+Oa��s_GR�[͎!d9Ҡ�����|���k��ïN;��Lc(�oQ��Ջ_-������']ފgO:Ş�2�i�3��3\�^��w������f�Y 0�f�XS��U��-ٜ��)��	�����̌u�/9Pr+��"q��"��R��ׂ��� 5<8c�ỵ�#�%G�N�;�N7P�W�^_�^T����^�n\�5������ e��(�Y��ty���G�ކ��͎ @�2wIh��0f<�s�*�Y��v� >5��e󂻘7�Ũ���s�^T#�������ܰ�g�&�v]"އ����`*@����M7��C�lSu�p�����FG�_mo����;�i��=�ӿ�
#���^���ՐղY�F-��䀄<H�0`{Op^"����z�W������V��x����IO�gWLQ��dM��˭ìB�θ�߀������i�����8��4��K���	�:[K>^�`��e�OO�[�ǋ��E--3Ne��cm�q���1xc�L�I�lCuՑ�Ǻ����1u�n��еP#�=3�U�曜?��L#��>ߦB�F�R�}O��~�T�}n��2����_����weOo��'�c$�3Y������d�{�������wm����}wo1ɹH=H�����U��\��z:�6�r�0�+g *��UqV�p5���BVu�mh��7��_��S3]w��hc�C�1��7����[�8��f�P��������(܃�d��Z[�b�qH���oBZ���z�\�}R����5�s��<�$KD�ְ�nm�A�[�M�=w}Ǹ�=�G�m���n[g0��x2�mC�nBy�}U�om�\dU�@��`����NYNX��݈����� uu����V�7����6�1�wPaE�Qs�;�ƞ����ZJW��
�>���q���Eu�V�z&��emr�^������;$��5.Y�>:���H���t��;k���c�8���WQ��TG�����ګ��S_����N�n�'8�kpۨκ����:,ޭ�h�[ʭN��D�j����gd���Օ����3,Jq�L�jư[���m�W����G�QGk�T	p*�E�OMr�;A�g	�؍�اt�j8._�'�.��=�ǞQ�V#Bȉm�۴S�攢��Z�(NkNgkV%Il��$,ڼ"�=km��o�[�q!�W(Ŏ��N��o�p��{~�= �u�s��u�J�����/�7-tL��%G)o����H��Y�N�	ɯԆ�ɾ�P<�������cdחҫ9n�W�9O�.:wڡ���4$ﶈ��v�}�t㶗K�)UG��[��}OL�x�Y��3�j�&uS�qr�1D�҆d������)���UNw��tZ����sY��
�i[����c���X|�8ҕ.n�2��Y�$i*2A�ޙW�u���S2�]9u
�e��d�݉���l���;�xsPk����haH`��.>3��t��X�0��M����W��ҳf��6��lҴ"��ر� �Au��E�4>0ukl``�� A6��c�42�2��G�W��_�zw���=+-nJ�S-k���!"L5�U����\%�[�t��ʞ7�)�G;�����noi�i�.Am�<b��ưT���:�v]��J�W5�ǳ$����Č����Md��m�ɮ���s�	z�g���2�UR�m�75�5o ��o3��o��z�ט��/�+껤�Z��Q/D��e�_c�q�<^�����w�V��l��I�ٹ�
v�wN�T���u�O{zJ�Dc�ˆNq��V�OV�wI�f�+���tu���J;���V��dW��9�o5��r�C�9�MuB>*ֵ�o_&�>���s:o����^4w2��/0�կT����\���Up�ȥ�w��5�+����]PkJ�Ȗv�)Y�jC'd�T%ܗ�݀��!N�.�������]Ѽ����[r*��ǲ�Jl�>�s�IC�4�;�7{�#��7 �Qͬ�5�7-��ݑ��A���^�7gl��yI�E�۹��hα;n��	lf0�ݐ��]����\��S�������۫ժ7Y�&�#��+��|�W`�VE��E�(�8]W<Y7Wp�]5�_��qB��#*�;���e��ȅNe�
a��������7�ع�M�b}K1P�t���68!@�P!����=�����u��>�-$m�-�YW|��J�?+,�%�<6zp����R�>i˻i�-�ȷI�9��E{���z�W���ӧç8��[O�L���-�����Ƽk�h��l�}>�O�#��Y�VW6"���5��1��M�j�rJl���}>�N?,v��$�c:��1�5�f�iV�3o�2��%�nX�0٣g�����r��~X|�JKd���I����݋KV�ֵ$���Ν:t�rR�I1�ص%�ӂ�kŷ�;^4Thƨ�S�gO�:rn�2X�w6�ޗ*z�k�~�toүkkJ�mE�������}>�8���-�t��X�l[��ƴmrz����qm͹��@��VfL�[-��}���{����{>|������+��ަ]e�S֋y�b�pɇ��ڬ]Up��,kI�f�3�{�� A z���2�w?�/�a���4W���2���uQ�`ᙔ��g7O5P�3ɝ�ॢgd��s\����@l�3f���$7��d@��P`��Ő�_#oDi9@JP��e�uF�/0_L��X^�0�9��:���d�Y7ۺ� ��@�sb�Z�l����np������;�[� ����Z*�e�@���y�")���Pl/ Gb�����_�1�j[��n�Dsf�9T�n�C{�pQR#ATԛ�v�y�*��i`1p:�K�wz�[݄����A��HͶS��Y��xzD\�w�T����#�H�Fn8kʤ�۳�́����dd鶀8�Ϩp�>y���	��`%w�:|%Ն�XY��3V��M��+SK�v	�z��Y�X�@��at�`�k�l��ǞT=Q��"�s�:�$^���:��,�������Hǡ��{��
f0PA��i���~�����{��+�.�kl�X�#][�\����Pp�����
����}x�٫�ٝm`�	CH*�x{��V�7�Y�}MJuv��V�7�iT^c�_�v��t�<�P��/
ە|ݧ��[�9��)s���@UtG굥`S­��?˦�<�ol�Z _XX*���*�M�N��ڱ̬��n���Q��я7���	-�˰	�E,U�W���O!�*w&�n��
7�۴�0Kw��fP��-��+^��t�S�J���O�o�*��a=R�MA��%��TN3]��װ�[����atm���7_a>��4�"@\F]
�e!7:��:�o3+�	�M�=}����^��tf��`+d�U�W����e��p�5�:���GM�g&�M�Y���Z'��=�4�4��A�]UJ���!�>�$8	�t���Cevq�oi���S\Wc5Vmᇩ~� ����p�y�k0�	Q���X��kZ��Q�Ck��E�iw�\�H6�|��v���|��U�P���tX>��$�Y��2_�������}�a�bC)\��x�m������m����u�p�H41�1
���"Ȱ]�_�(��c=E�"�z�\M�K={�D�ۜ���5�[����T1vD�����QC��X�Y�K�<k���v3h���|��{��t괬M4�u�S�4�R�3WX������b��٫����j�)i���������y��t����|�R��ǆx����!��0�]���:��������u�S[R��F�����!��Ά���j����9�5�|�G�Ĉ1\O���jm%��MY.�r��� �|s���?x �$9�=l4�]�:��$
R�+�g��L5ۗ�g�tt[��X�y�?p]�DLb���[؛�̖pc����LV��+K�Ϧ�ތ&�r��tH~of>�O����"�?���Z�מ]����:�I�2�l���*:�O�V�kxW >��v��htP����W?����v���E!�rR6ŴdxX���34�7S̶��r�!���Wzn6(��ޝ���wyX~Qj���heWL�W&���ʺ�iU��"!#Bz��0�Hj|���׸�Oޒ��~�Sܮ�n��_r�ס�n�/������r�MG5�k��ƈ&��^&Xb��8���;�����;��n9��{���Nʷ/g[��#A=�Uot�0��L�ಱ���Xw;�_�7F�l��K�%�����0�Yg������Ϙ2܋���
<��EU� �[)eO.��%�~�q���>��,|5�����m5ŀ�X���B�v�],����4M��7sB����;%� e�@X�6y�;�O�)��k�t�l�Z�M@����y e���v�#�@�n>�X͡�.,Vv��ږ����Jb������y��q�4A yr�o5t��v�pv�f�
4@�VE����W��ڀ�����g�01P23�I�v�M#�>d�3{�^�Q�f���m�0ےl7KQOѓ;R�p3���k�b�i��"�;���LT��R=��@d�ߪ��-�oCJn/Z���Uq,Eg;�o��)���UrX@�2ee�H���*�>�PP�5�Av3^���.�2�:H�
�l�M�5�g�^D��Č�$I����<9�����y|�w���f�t̡�%9Z+1��չAZ����gfk9�YY�2����v��d�kX3�7=�(�B.,���m<׏I���p�ʁ�0ڸn�p���z8L�˸ٚD^�!u�ǔ"�Պ�f�gܵg6O��@�������䥾��������?n�⺔�����oM�hG��7�s�x^T�@t#b�Ú bJ����[z���ʔ�x�C��+{�s)�W ��^r<�h�QZ�l��+`[�Mê��8&Y�x8�;L�CU�6�!���@w��=�=j+�އ�Ĵ�ʌl��A>5�·tA0�1����fn{�5�$��Np��0k#Pܥ�^��񜢠3�k.�n��^^��q�.���	��n|}��!��|-�5�..|iZ�Z�Ov���p.��b�z>�Ckx�7�9�P|W���X�j�o^ҝ�<�hQVf����$
�m����0���0=DݏL��l�l������:��%M��qd�÷�`�h\(��ީ�m����5=U).�o;OChk���RF����7^ M���,���ժ��b���Pǣڬ#���5!V���ݮ�+/VU<�j�c�{�o�%���SF����3��n�'z��|�|- ��8Z��A��/z�k���o+�Kwyo!�#ȸӪ��T[�6%reEE�����5�<��` f� o ��B���0������w�8�;�Ey����>��������~����)/��s���p���ڊ���:u[P�	�Oa�~R9�T��-�xQ��3�J���gh!��-$_���|����!5��G
96� ����j���<�V�cΞY��41�Xf�������*�uY��1����銲�R=7��|��j�-mÈ6Wm��e%;�b�Vx��!?g�Cu�j���O>�9��l�2t�]4����XIm��ó�`Ǉȝð�؀͸H�&��>{����"@Y!�L(��M��z�����ae1�F��@"�9ܗ	vQ�p��ձ��Bޠ:����~�Ɏ�T�@@����I<rX��.��	�n�e������7�i��e�X{�8�Ϊ*�kT�4N�\4�eikM �V�h5�E!�F���n�M*j�Y����q�ǝ�����P�\�>C��ٚra�A�o	�J7f@����}v0���d���O�O��ch�jxk����/��r�M���Lõ�Kj>�X�&�Q3�\Xb����
�z�N�i�ͱ�MY�˙.���8��@z��`  Kӎd{Nꮮ󿉱��p�{"	ٹY",�r�o 	�n�:_/��)�jG�wȲ/��;O�@p�9蜛�����#���U��oU�~�K�{2<���F�6.��ց`s�N�M��x>߅��F��A)!��]�:X����O���D�P�g)��58^����s�޴��of[�n���Wޡ�x��>a�j0R����~�%i��L� *���������M��i6���`&��N�m[�L UM�'��{�cU/r�"�(�"�2MMגɣ�:˺�w�:)��e}��Z��K:��.0+��9�K����!G�/�f�s�������ʢq�U����f��ÏxP`<�H�س��٢a�9�Usjo��H���㕠e����w89��������@L۠�g�]�Q;�6�A�18��&Y�d��(�.�5v��E�K+7�r�]�(wW��~���.�׮m�gv�Zǘ�~�lRa0� ,��szR���]�q_΋�]�ʛE�K�ʧ	��Ђ_=ַ%2�7��*�P5x����� �o2K�.a�_d��<en�,�����1!W@kxWT���f��s�nɄ�tJ�Al�M‍QN�'v��քM�~>�a�;1ŻU����̽7"8싎�QV�}�>�H�����J�R�`�ۜ"(�v��^7�'�kQ�$Dc ��Q�ŦE_)wnWly�6�����ٖ�t�J�h��`�v�`Qy�N���h��Wy�s�޹ߦ�����	w����k����P�������Q�TY݅������� ލ!���[Ι����Æw^����gZ�2 8�8�y���5YO|����[lv�0N_�=���,���O���y�p�̓]�Ei�j�Rl���9��Br�D^����j�X�7��F�������٦��w*�[T���0�����&��e6��2p87�7j͸6[�^j�1��]#�&��}�:V"r�1�lt�����cHHx�t���N<8�x!�h��L�.{�<�15.��U���\lpo`�v[%Rڼws\��2���N��e�i��~���� ; ��Y�ruD÷�T�|����X1���'蹝����/���E�I�������=3f03�?��W��@���E^B�Z�ڙ�^�޶�Sq�<�����>�	|�)��V�u��p8K�U���.����㜾��Z;'V�� c��z����eM_*~*��ORW���|��]�7耂�@����u�1���yX��R$z�Z�K:U\�s!�D���*|R{'��	��_�``���%��+�7Z%n3]��z��Nlul�%ϻ:({�K�>.h'�����8����!��;�Q6oNʚ~��L����r�b���6�w4��
�Q�L�~
�C�����u�I1�1b4�_p���������S<���j���Q}��e��	p.}��|n^=ۑ���A��ύ
Y�u��AP��~+�(ff�=L�H����R��G�Ѻ�7�褑��ܭJ����b�8�$����ߏ�x)M�׼�Չ0$v����s��!��g�n�qn�Q.k���1 �'�#��x�;�ι�?�x�� ����d�u,t}rnTW��^�c7��z�6Kʰ�ʑ�*7.�\����p�L��1Ό�� ����`wi��<X0%ó�3�3�Z�.�`��[�˔�4��z	\|�{Ӓ�u{l]�Mz���8�� �D����gYV�v�h L�U^VMS6\B9���94sf��R��[y��k֋��4g4�����a����AA���.��#�7�`�N�&�3�]p�E0:Ȩ��?g±��-��/��'�\2*�L��'nI���+���z��'�|���X=֖����L`ʂ�`���Pw��F�F#:�2v��|48�:�3��VUC^1�A�gU��Hϯ��8�$v}������L�B=�+�^=��s�uotU}�� 6��n�8bt:KH�=��%u=c*^ �����w��҆u�N�S�\�e�$qW�����9Zqc�--��;��S5W��uU�X9j��v-:���v
�����N6�q����SoS����k�䌕q�f�j���W����r
3���q�<� ��8��We��yؚ��u]Q�/��ovao�o�I�T�̼��'����9P}��7�C��qÇE�lL؛Є�E;ڱ�S{d�rr��|d��L\����/��^N|��-;��}#λw�M($ǅ0n�ӆ�k`m�к��ۛڭ��*��V�P�g��i����N����V'ȸ�a]ܮZ���m��S'{X����r���t�z3
ƬBr�>�Qx�d�:rܨ�W�f#���ͫ����k!ǩ,bhJ�-l�_w��-Uc�\&F9w1 �.����1Tm��MgF^�n���ʘc��i�/�E�lx�ȳ���[(�ǉ�O��$��k͵3�VY}%�ws�2gN�Hv3�A�n\���hcX�[�u$�'ek�j�+1��v���\+�c�+���K��vH�٪V�#���eS[si�;W�
�1x�������]���j�4��I:"躆����X^�gM�k�j�ct0zv���x
�Aa���+vypє�ӗ["/��%x��}copp+�e"F�α=�$��� RՅO+06���$:�A��V@~�ؽuA��w�� ��	-�Paނ��W`�:�_8~���Ɗ�.�B¸�U�}o������A5���mL��U�F��Z;�3&�"��p����J�r���J��K~�;Ov_Ye�y�n�n㡜/X�*s�R�Lvr3UXa���w\tP~uy��h����YJ��:m�Y9��Ɯ:(��_����Q.Եp�{�|l�z��Dm3���Ы)ƔӵR�Deu
�Y�i�Q�KjR54WM���Y����d���Փ/j\��T��'4��c;���06�=���j�$Yr�$�vȫ�[��U��J����������Dbt��N@kr�g%5���Z��Pj;�ǩ<���%E�C5\�Ǡ��u�]o�ܫ�����6��5u�۲,�xꅇ�z���a��jkS%���d)#)�r�ɂ��*o'g���
���\nd��O"C����L[Ujb�=�s���(�H�,��e�e�[+�NB�,��3�k����aO����y��tIN�]cN��Ct�(�᫖w�Q�kwl���� ��v��f�8޼R��nm�:�I2��ɩ�n��;��+a7}�eo���b���Da�e���
��m�5�&�n�Zص"��uZ�oQ���ۍ��S�l��N�iy�3ĺ �<Uz�M�|m����^�z���|z�zښh�4�c��6�u���ƚxƘ���j�6ҴҶiX�ҘS���01��[����i�\��cF��R,��w*��5$UAeպ��m������ob���l<�UDlTo�]6�O���_jM�<<:~��$r�n�5adb��+^"��x�N�MS�7e�Kd�N��=:t�jv��Z��i2�s����Il�j��XϹ[a��T���������/�I�m��*Kb[�1c��oJ�ŵ��(�9��jT�æΝ:t����c)�76��-�k�ۛ��ޛk�+��˔S���Ӈ���,NQ�}��kzj��V5���?He-���a����}>�G,�Fū��x�W,e���K�2��Z��On�XS�G�O�N��ũ�l�v�Ƭ�m','�漢S�����ӄ�q�K&Y-'l���5|�\ѹ�F�+^f����nU�nU�X�!��"߼A,���֒~.BIRH�u�!ו�as�&�Fe��Δv����kBX�gQp����Ŷ6�Ǌ��v3�{�̸�ޛ�"��`bP�4ҫLK�uqmf���c��1@��xr����v�!���G�����-7�#Z�>5�<,��1X}@!�J�}��3�� �>$3Sq��uʟ�䕓 ���>d5�d|��U���=}��!l���lL�N�"��� S-P����l ���c�<޺.�V-�ڌO5���UνgL�W"�T���t�*��2�M;��D eD���IoG%�7|<���	�`)j0�ep�in�ĳiH�c�f�@o8uɅa�Zme��x"�@�;�Zf�?f��c�x����:,ǜX��&wT�i[b��oa�ַ���,����	����PC���=-��}��d>��QA�:i[�Я�&��a�w{��98�g��y�� 6P�Gj����wr�.���=gM�O+f&�]H�alVG��bM6u���_v@�ǹM7j�pA-sS7/��tX��,i�t�_q/���f�&�e�l�O�a[����]`��9���@�ќ�l
����c*��d�E=��%��B;Rc�H��E����;A����=�Q{�2��:[�`�����9n]��U�5�O��&^�>�
»����q�&������}ܪŊ{M�I����z����� e@فW�%��n�Y31u��DEV�.�ջg�V���KFe��
ɀ� *���M�@�u�ثn�[1<[@-S�I95�7J �R͎ʩy���gh]�nl�Nǲv���Lg�($a�.͠2�4�Tg@��8�����c-<
l��D���%O�8���g�/6��Tyv���z�X�xv�f��i�Zz�� [�:$�Y��ޑ���P�����ī��Ln�;y�NC�l��@8�r`�vK�O�=#8����r��uw2֚#j��-��9 pp7pP�Ƈ*uS���v%�k\�wpܧg�R��'x� ���h�|^���/d���Ct�lLx�甶�>ɷIm�Q+��iArc����vg*��뫔�!J�<��u˴�k}��vj��	�������M��4����f�V,/�I��s2�<Uy޵��٤+�i�g�c<]��c+q�}��~� ^ �=����K}w�~���j
)�	�ҰM���Cx��O��r�ϯ�p�5��]p�����.���<����S�o;����_Y�.%]���^��R,0��������9��fV
̻մ�m������ӿ�xG��15�^���Y�E�ց���
�V���
����$��컩�`��.��]���99����ZF��'�B6pP��Z�U��5^��V�#���r�ymqnf�R�C;�\����pH�{@A<w6J����E���YW����f�k^�N���7�1�zߍ��Ur��M`�]궞:x�3
��I�%�����Q����V	�@$u��k��(�]�S���g��?<6Ҝ��`���Dp*EW��d�����6���9�>����w�[��x�[�OGs�xͱ
�"�k*�(>�H�2,�㱳*5�c�]���0u����v?�أ5I���r���`6��+R{��n�7u[!ްvL�{��엑V���qE)ޥ����t��Ź���>(����8� � s���Z
"��o��sv�ֻ{��_ <,�	�
��]�Q���a�t��&5o,����ܫ�@L	N�f��������R�:f�q��b�uX}��n���gדݛ]�x��,$��'$p����� :� XM��k|�7���;��HҤa����#m o8�N��ٰ�n=(wM�f�����S��T+�L����K{r�q�#��fU1��*�x�n�i5z�or��z`+2.lϖ;dԀ���Ϳ�y7*	h��U鎉�!�@�]>�o,����Ys��}��|c+=U����y�p��|�:Ï{������;C�v����-���X�ks��� $@�Ai�z@�i�ta�`NHeP�lf�fT�9Um]��@啱��$�p�����mɶz�sb�V$J}���7��먗hi�	�=L������ꯅ�hcV��ֳ̒z�vw\���5�4�%h_G�����F��7�.� ]��E����L�)r�x�)��5�xf�YM���$��3.Q]�F����e��y1��c�c֛m�Ͷ�M)��u��f��y�@_� %���v�9[jT�u��8��Cc(?qثtf@�Dt
�@%`)X��E)w�t��R˱���[��g�Ik�����AXf��7#	��%_�$㯮��ߵ��5��+�B �pV�9a.�t�zZj���37ٸ��&�;V�o�s�lr����x_߯ǆ������� |,{]��g��s�7���$��l��0��;�����m��d��q������5֦�4j�t�i�,�l�#pi�׺vRۺ٪�����3�ki�Q�A�y���^�*�-	��k�-���)��p�6����c��:�}`Ubu�O����Lx��5	9��j�}m���"Ə0�4�z�Z����fcQ����g+�7��'�EADT̠щ̞]�p���g�ؘ+�������ݼ��<]��g|X���܂��iog�Ρ�f�C�n9�Ì���Ţ��;kF3�g�We�ֆ\0>2noQ�V\�E�§FR5�y��=��t�s������+��`��kC��Պ���3%�f�Ty,��T=�{�@:�[_��-���������fc����s�\��ט���9��E�'��a�k�����#��xk �u�ƻ{:)���k�u�)���w����������3B ۚ����P�ٽ�"���«�Jk]q5�3U�'�A��`a�4�욞�Q����1F�F��fCԄϦ"������#�W5��W���~�-_�3b��l5T7(�2��Ek�˳'����vAC��&62�H�����<7g:�f�wT�4W����0:@���G��l&�mM�m=L���Rp,f��[ 8I#K��+�w�
���Wʢ�.ݫ�;+��#���bxH�9#"aniZ��0z:�OX�rC����*�6�k��^�wox���?���9c��b�չ!#qh	m�o��Y�2J�UU�k'ST�=6�g(m�iW�,��ѱ��-��V�]�啥i�����5]|*k��fYoa�+:äk�魳�"�r��Lދ����w��:����ݐ�4�q1�Ҁ�<��w�(QF@����Y8�;0v���J�>���ޔ�q�F�І���֝;Y�t�������Z����)��2]��h���g kGrs����~�WD�"Ȫ�;pKhv(Ȏ�7j�=:��V*�ӡT�Y�PG&�WN��� X����*JT�T�s��|	�9��f��8@�@wg��d2L
��0�1Y��w���炻�?7d�l3��RW�u<�Gp8����W�]��X�3q��B��R�a"��~����=������SY��@�n2���g�Bњ�nD�;�g+��W]�~:�,
r�<&��H�!��W;f��ַ�ﲀ�Q�=|���Ouf;js�����حoY�����~��@}"����0�KƄV�E�b���]=d��'�����Ë�q[�{��Z��m���1)�ŉdC)~�b�5ok�.�x��Vܳt���a�H���*��8"��)�`��93m�� B<#�c>���v��H[��7���=���x�<�Y�w�+�����5�18�Ç����Q����׽�\��<�{ߝ��R������^ 	�y��
��&�J��`sU�����E�4� ��M�w?T���?��c�#����(�k�+�x�.!#Ϥh�&5�J�O�� 0ü?�$3s�i7: ���gc��en��e���,�x0��F̶鞂6���ާ�rB�U�ؒÚ����#[m�1�����{dq��X� ��ڗ�����9��`$��)�9 ����<�/隷�o0�ٰ4�ܲrˀ^�C^�}�r���v�c's&3��*Q���H���I�hNp�θp;D�ҍB��p�*2ʚ%� �Z`�j��\�s��9��>���5�|بɶ��d��jt=1��@�}7)F��}�������?m�όy������&�,m���af-dy	N��[q�+��ad8��sv^��S��p7~�#�Ρm�ovհn�d7�Ne��L�����|ʨ3��X��l���D2"3���U�;�cT�:!��Q�+.���b�.�k9�d�=��u����;��:��+x-!��w��lsU�|Ⳋ�F�r�� ��D(P0C@!�A�e��i(�H� �x� UE={����{aC���㩌���gϾ�8u|�	Y"�.�>�V� ��m�v������pc�_N�>�γ�<��T�?��}
�&��
����;���ֺ�H�=�U�z�`wQ�ў�@��=�Ɛ,���3��u
f:������M��H�[�z�G��ۼօPX�p��RaW�
0Yv	�W0��'�1���U�#Iμ�r0v@j�eI�IQ[��x9ISf�x4o�����n-��@]!ݙ�7�����;y�Է�+�8���j��0�vt_l�#�nq��ʪ�5^EҀ��X�2���!B��Tu�``p33�k��!����:�j��.A=�^�׎���[���� *�ʘ~h����3�<�pO6L��h
�5�T>��x]+dif{�j5[~Ϝ�P������AA����}�ch#M����@��V��������|3�y}vm��7��ƨ@�4u,�םɝ��[[�n�U��+s�-�36��Y��c���K��j&�v3#��{�q��?�?� � [�9��Z����9]�bVol��N��BC�榏i;S� �S�����O�F%Bu�:g͉]��gy��P�es�j����7N@���n�>��/`g ��(��ۤ�ލ��'[��#��vX�oOw��
p���(p��>���������r�Gi�8:Y��#8���x��E���A�wM�ck�ש\s^�f�'�5b��]���� #]$9��vÁ�I����H�h�Ikc ��#@�(1f����>�9shZz���t�&�;��	�,��WS�`�!�c��Z芪�*����1f�W��`=�^Jߤ�Oxͽ�_c�}1��-��Py	D������O�Y!x�� �hڽY͎��@��{Y�ńy���j�e�<�C�n��u��-�4t�a��s�6쌕ƶ��m�MUn�lSՎL�|��gHbٸv�n'�Sg�:��j����ǒ^�F��T5����읂Z0���w���U�*��s�2d����	����� �sdUy��o�T���R�.�F�z&������Ě��Ko�W7��4��EYp6��(md�����A��X�0�t������]�,��G��$}{S��k�QV��	uKV�Z�啷Vr��FԮH�Wj'"K2����oK�\�*-k�����§'�Wp��&�5z�r�ݤM}�A�4z�u��[�]��Ҽ��t��#\��ɬ�1��}jܦ���.a��jY��s�PӇ�%�\�(�Y��>̀��ª���]z�\�;�IM஦훨o�)=��S����H�\�c�q_S��ݕis��mZָ�4��-�:/8�:�<���)�ĚWӧ2���S蛦:��;/k���DŹ6M1��-}|�W.��m��8Su//S2�֥eL�o"fŜeo3��r:�M1�Ԯ�i
��
����K{�ٗ�f�d��{��M�;2��Պ�fP��J��ab����w��V�&��$G�v���K��p(@C�?��𴯔ƾ7�\x���Λb�q^W��������7h�l!O� �
,!aN.2(t�d��8B �a~��f�g�ްpm�Iê�oE����{�	�G�2��UV��9I��W^'d��E��+q�s�j�q�-���w�qJ��.mU3��yՍ�ۖ�3�n.�Ȋ��0�+1���t:������r^%�ۮ��"w^mR�Td��34��*�R���������w,��W!�\t���t���}�wen�yh�AB��I�����]���Y0�w^"��7�'8���ے���{ӯF��8W�����^y��n^ᇮ�"���gTt�,���&��V���� ��=��}ٕ���F���P��^]!+)a�兇n�'�S���wm�u���ts�u�EYc���M묕���Wy��������;u)��&���ٟ���<.��*,�syw"=ĩ�:��݃�,���L����GT��%�a*��R����Gl�%^p�w̷ٙw�<����]� �fir�>f@�t��F;}N���p��87՗A��]։�1g�b�Wu������dє�d2�'v��Ne�u&�ΎA��[xcuv+�_^�a��f��͕[�qUh̯��n�8P`3��ϴZG�d˔�V���}��5E�J��匲)��������*���"e�[��v�+3!-Zn��M�:t�ç;gm�s����݉l���cw��r�^R�2���L��͜=>�>�I�k�ʅ�,�|�7R�>)2���VNܣ(j�W.��6|>�9�ĵ��[�s_��BW-�;��w;��(��l�e�4t�ӧ�Iůů��b�S*����W"x�@oMsX��ٷ��W꼯����}9>�ٖ֪L�c,����L�e��[��Q�̉M�>�������oqk�)򤛢j�-��Bѻ�S��m��<:|:t�r�>\��d^��m�%�9��ߵ�[��ܭ�I��MWnXfd-��3�l1���ְeKI�#)������w����\�ݤ��y:klc���Ҿ��R�1e���S������:�rM�3���M�F���o��
  �� [/䳭����Y��pű�U��ZƁw�ε۟f�y��zWK�%ut��[|:/��7�7�:7^D�95�� [O*{�vd�X�ӯA���5����֤�wZ#B��o�X�v��ݿ���~��2�mv�![�o���6
辇Ѫ@I��y�t#eoP��m�iV^^й��M��6n��P�3�[�e�,�����e�dB����� WoUJU^cF��t�y7�{nM��/˾wՓ����d �`�����\�B��kֽ1{�̾grywwofV���/C�7=��1ڧ����m�V[x�Yy������k�@'c�t��Ǟ�ͼĶ�[3l�5�3wKAq}�)(���o�r��k��$�F���{w{�Sd�9ۑš5%a�hI9|�&�C{w�}��nw����;:�S��/�r�����X�ޛ�\g?p�v4͋����]:�#CZ�tj�Jƅ:��X4[�UnJ���Zt�5wي}Q0Ů�����(���7��n���3+z�2�;"��/.�s�� ��� $xLX�6��/�}��d>�rx-���_�m`��M�7>IV��$UU^.t�<����l2�w6��j�E`���1w�Zܺ�S��۳�h�(x�8Dķ�c���w�\��4i��Yn�o��;�q�g%���'�GK�Z�4�<zc�,X�t6l")�7.õ��Ce�pQ��zM�@�`:=/�v	�ג
��s��i�z|=�sF�fˮ��
8:[7�������\����*�g�5��j�"m.6ro"�P�b6��.�h�Q�T�Pn`�h0L+��Y����7��F�g�S��-'_i��\:�Ԅ�y��`ef�#m�q=.v繦�{^w���D��P�ϵ<:������ZX��;?El�nZsI~8��$�u*�:����F��������'[��>΅s5+�O&��p3w�9�3�9��z�I�	Ps��%2�Kǣ�t@�e�ɫ�)Rs�wk�FY��ت4I��������Z�*���ok������q����6�gJ�3�t�Jowlՙ���4����v:;5�"�6-�����,80�c0�!�h���l�*S�?��4q������Æ�hW��}j#���S�;�,@��Bnlf`�=1,3v�1�Ѡ��-4p��K�5�
��"#�#	��r#[�ʀ8�}��z���F�N�aJɞy�M��퀴 AP(n�S V%�4ko;�1��vVe�p7]�0�l��m�������z�Vy��[�D�#�]�6��a�Av�ۖ3+�J�q�z��p�h6Xж-}��<�Z;�۰����p�l~Q�q�|��$G~ڍ���p�)*�p:'���M;_b���L��Y�T�^U��ɳ�gQz8�(	��	_��z�6�� �ݔ�/x��Ss���@#<hT> ��V��K����	����&�u�M4�K�����{��N�5�ɭ�x��U�UK&��<^��=��5�r����n�rVէ��~"������]�Yl�_�	=3�&��#���i��<�/gne��e�0"��)�$�m+'`�x{�=�������ja6ޣ]}��F������f֭g�v̾�:0k��M���>f��5O�J�����%�x�p;3R��V���m�Ob���یY=ddU$���a*����W���YC��;�:���\�Ch�އ�=�����5##����K8+7� ���kk�de�՗3T�j�L7\�`�n��}�zm�r��%d��<�gS;���{j��[r��A��5��
�b��J�S(�g�m�Bz��o7A��L�0;�c�q	(۬�J�5=�ty�Q�m��f�	����������P7�����C.Lƣ7*�g�S��x�3��=����dϏߗ�h
�� y:��*��	�P�_K�R�L2�o,���iHb[�K���E� dL1���	����|�u�|L�5����o1�����֧��nD���D�IjK�f���t�S1L_?�����>�ll�z�׭=DE��aB�{k�v�����êL*�`/�|~�b|�GI����`�2B_J��n�db_;*�b�d�*[��Ꮋo����!�Qf\�]l��8����'��]���.W란�Y��SoJ����a%[�]�g:�7�X����.@W�bj��!R�2��2��>�t��w'�r2��7f��~޲��^��  A_���t��|���
�*q���Q9��1!ݦG%u�䴪w���SSy�ctL�Ok6
��5	_�ׅ!���4�i�g�\�=�"�I�Y[%]�� ����&o���ٚ�7[2�C�؞E�l��^o2XU���"WP��ʫ�<��{2��_����V�Rd
�:'Ȭ���0�4���*8���ٸ�OF�vez1�\�ȇ�HCH\�z��f��Y��,���SIY����"��KL��r�@m��-�E�[��S�����O�R��}������w��L[�U�;��� �`1]��y��.�6���?]�×^��|跚V���V���!D#HTg��Ϣ?���-!ݵ�?9NSW�xB=���d�ڭާ�~�W�����Xs�WUN�lfە�v/<J���ڥ����>��ݾ��-���g`�lzy����<wk���m�#���4Cw�l��m�|/��s���}@��&�U�������ƺ{�q�j5�D'���7hu\s�|ㅍ�γ��e�pk���<w<��}�T��9B�0�s�<?Q�[�{D��↩w�
�Ժ�U����L���K)�ۋ��9�`ؚ� 5�y�@>)v��N�g�#Ef���qT�]����Ɠ����u�=.�|lX�ȿ7��n����Qb���m�x�������؇?s_µm?�M4��[��L�E�!���&*$馮�ܝR��c���'uMⵠb�~�����k��5efv+�<c���):x�]��Mq�U��M{�q�m��U�1�fxb��)0
@��ccGe��o�c��Xw�*�+���0�f�c+����T�ꔬ'�{��ف~�m%J�t>�����J,p��{��h�鈲h�deq��j��X��a�m�(���q+\�@������f�WeO�_*�7�|�c��?���U�q��r�;��j�.�W���N��ࠃ����6b�ҕ�h����D�!�Q���p�U{��+�pB� ���0I��μpU��g޸�e��I�����q�
vp��=��y��ʾի�}Y ����P��*[����N�����X�y"2wwh�`ޭ���Ϲ�*+rB&�L������@>���ǎ׌ɭ��=q(O]v��S�:�1ݔ�d�ِ^ܣ3LǪ�����m(��3+z=(�����Iڭ8�3�����OMl���j�z��K� ��+z~⧆�#mng�5���ϸ淸��\�� ���0X,�o�c'�zF3홢t���/oo7�;�z�ڈ�����w�n�w��"B�#3�e�CJ8�uuT��c�e��ɀ��z��<T1���F���4���%0;
�$E�nK��T�È䄗m�Z,��.y� 3��yrZu�U�'��S�Q��9���L�yz-��Oɐܬ�V��wZ$��ىKYոOM�:z��Y�w�̢r���{�@��w�]���T{�gT��Z��\�r��")p�ǦbcTX��^��7�Ԇ1X�-�̺�'3J�Z���1r�\{��XOD�9?V����q�f��/hӲ��2@W[�Q����N��"��L�z;0�c���x�����[\�'��Gl�e]�9�kSPȴO�j;LU��s�S�u��/8E���|��TV�Ƚ�xдpv�P�jC���+�
�X��5�f�FExtg!}9 ��B�N=�xʱ���-R9=h�m�����l����>��ο`)��U���]�3��Q���aC��k��x@`��ނV������˧�ij�C!#z�� ���%<�w�xqC4��u�ꢦv���@��|�B�����>Q*�m;�e���Ev��iꘇ�k\���"�cԢVnW%�u!��~y�٬\w���`�"�\8fQ;���<�BK�ޟN%w�{WL��؟���Bk:�_<��W�_p�r�Ч-p9YN�8��]<FqV+#�/��y�����k�j��6����w��+��Ʊ��T��q��r�l2����<��5D��g(s� ý˻��HƤIɵr�c��ʳs|-�e`����:=�Y��߷M��W��U'� $M�#|�@n[hv*÷��]�ò�!vu�"x��ivTN��љ�[��aN���洜����V�~��;�iϮf����W���G@��F�,2���*�U�pn�V7�3�'Yb�R{5rLކ`�t��cU�#�A�i�67Nv�ٽ/�>>��w�Ru�������xf����� ])����v�LȜ���y�&�Jĸj��+���S�53t����4�<�w{{ ��M� �d[۱S>z���#��k��Qe�?_��/{������EZY;^Փ Z�x�EU��$�9�Q"CN�̣�/��)�C ֣ה�*V�*�%m���u��P�}������GL3�oM�k㣶�]�|���� >������蜡�j��B��7r'BU��Q�VC��:�u웣��V�9�ك;]>�1R|�7��!B*�ݹ컀��Y{#��޾��32^I�P��0o;�_o%eAG��T�b\�h�z�;1}�y]�Q�9����۠^�;����܉�[�
|�z���N�WoU��mFq��բ�ݾ�ҕWs]w�����C�h|Ny��{ժ��8`0G�D�2�<myq��.���5���[�q�ca��Y����i�݅���ۆǈ��'t�r�U��ƀ���6
kؕl�s!�)�*t8�R�V�58��3��ѼX	������ζ��������>D�ܶ�wm�y0�ϻқz����s\	;|k���9�ѡPm3t��'���ŨÎ��I`wo)ݘ}�Y�*��,g��Yj�B����-�F��}��U�נu{F�Cq���}�� �]w��gU[c�o��o�q�˝՗�/��Mc�a���R���Po�?k/��_��|^�T0N�� �W=��W���02H�H�g�"!�ߟ�?� B�d�[��挚�27cǹ��{��I����B��!Ab��!AR$(*DB�Ȓף`n$���HE�7RIHH��BE�(,�DPY$"��!Cy�$B��!Ad�(*BHB����
 �򐆷�4PQ���PY(,B��PT ���dBAAd�hPB��dH(,BD()$"(,$���	��!H��$�$��Ē����PT
%���!
AR
A`)%���&�"`*$PXF��5$���PX
	(,�� ����D�J5�&S@������<�c'��?��HH�� H�!�X��F}?�������w��?w����������G�����?�;W����?џ�����S���=�������w������?���R$�$��������?ʒA"O���L�%Y$�#�?�I���V1;Rl�����?���H�H�����?�?w����#I����'���H���q>���I�����K'�2"	���	-�%T�I�ɭ�[kI�lU�V�j�[���m��e�5��ٖ�+b�&�6֋l[X�&�MT�������[&�MT��+fmlҬ[cke��UL��[k�e���3VJ��ص��f��k%�+fkf�l�l[X��km�*��Ŷ5�5�5�[f��Kl٪���VKl�l�kd��[)�ɭ�l�VkM�*ɪ��ƶKl��Zkfke-���Klkfkf��UKl�e5�-�e��l�lͶR�[f�i��l��)�*V�-�KlҶUMl�m�[4�̶ͥY�ٖ٦�Ml՚ٚ�-�5���-f�ٕ�5�Kl�-�+e5�[d��m�kfke5�6�-��[3[%�5�[)����YMlj�k3[6�lkd�ٕQm�[&�M���M��l�klkY5�j�lkd���Ŷf�Ml��F�S6�5�E���,�[H� �<J����A�E��KRjڱ��mm���6�Ml�[�[��n�{L����w��"	h-E�H�	���'�N�_�����ߴ[��G��ğQ���������H�H�dy�����T�xN�L�c����������<��$I$I5�G�S��t�7���I"I��H�H�D�����{?�o�J�A"O��?a����I"I�Y'��G�[����>'�q�O�Ln�7Fѹ"I"Ii����ޑ$�$�O�GR�|�~�4|�|��ԏ�S�?����$I$I=�C�?Б$�$�#q��2-������꺟ȋ����j?�����I����"����D�D�Ⱦ��,|�~?�4������=�n?��p�O���$�H��'��4�A"O����}��?����ʞ��7������)��@�Z�o�9,����������0�O%��UUT�
*�J�"�QP!B��T�RT�DQ
�Gw�dQTJ(���%�J�Q%D�*UAI�%2�퐲i@R *���J�@PN����%R��)BPQ{*� ���@ѭk�-�-H2	ml ��� RIJU�Ӫ1��,�h��ZŨl-� f�6e@fB�@B����(��e�`�	(%����́�4Y(�IA���B�X%�h֚U,YEf���l�%J�k �ءL�*)B��
��u�,������U�� �$�����J��P&�9ˬ*ؒ,�a��,�3d(�2�6�f�` m�2+�P]�iD��(���H8�JR���P�������V�j�l�-`U��JB�B�� 'X � �`h,P �(�-1��iAF�4*I�Ѷ�� ����� *�(P�f��� 6,�[j�[T2��4J���Z)�а��@�S�q�+F�4f�F��`���hdM�*h�-���ұ[ 琠   @D T� ����R�CL&�2 )�IJJSL� 2 2@9�&& &#4���d�#��@��J~����4ɣA��4H�4�&L�E<�2Q��<�ڐIꔈ"� z@  A��կ=��M�*F�O�֥���ҷkQU�?�4�֠�����d Q@U7"���̏����eb_&�������V���eS$�����j���o������m�V���՛^���2 A� Nm n�d��B�ӟ>t�����I�g��i�.�?������yw��5�����y��^=z���s�c&��(2ʈ��D�J�"��� ~O�a!.H���"2Cj&�b7E B-�`*O�(��?�Gfd
HKl3!I�B�!Hj2ˌ�d�D�(�����+�Q��m�a��1��d�$��(��DBf$)��ҝ���?�-����8�m�����r �a���Rڳ%k��� �7�6�װ}���6��&j�C�)Z"�!Qn�
�op�eÖWq��q�c��������߀h<Y�l�/Q G�]��iGa�� r�`'v�&��v%Ywv��fL �C�7K-ʌPГL�4�Ҷ��{[���N��P�P?�Z͈���Um��C5�Im��F-53&�Qe�N��ެ�p��qͳaH�E���sI#n�L�h���X�C�y��$dX�T/"�U�Ij5�k�q�3�P:�!`z��j]\����	�cw5��V��[wE���)�i	�g4�]���Ӵؗ%+u{)֧��rj�m���)m�z���n`ô���7�FS4�Xj���km(K%Cn�4�VԆ���L���Ά�d�e��¡[sbۼ5��̳L?�`雐�B�U٪�e]e�P�q
T�o,�8AqZ�14�f�)�x���װm�m�{Y�`İ�2�%���J���N!(KǍ���
�j��4���N1UfY<?��}�R�EDԺv���5�;w7�b:^�D�:��͈/�7V"FSʰ�4J��øʨ�eԂ�cYR� $�viS^V��Dv7F��X�G0U�ѻiB�E��2�k���rc.�z\�v\�G*�U��%���]�1���1Zڑ���c�4-�ֳ4NދV���I<�UB[*�wb��T�h7���,mP6}�3�bFP�9��a�`)Q�m���q�֩u�*K3	��KD�V�$�2�oP2P���^���jaDX5SKfL���;��ͻ����&T�����M&,}5���d
�p:��{[�*@�{��`k�E��\�	ف�܌���:��	1-Kn%��:�q����OBM]Sߵ<�z�"꥓i�R�
�$�2hƝ��r���ٛ)e'B�M�ZaN��T�be�T:%YZEF�P�f,��S�7*�bHA�z�m嗃uY;���T �d��hV��5>p���պ�M���aM����2�΍ܥE��Tl�q/����Z�{z0&'2]bmm�[��B�Bbvpѱ%�G��(�ZЪ�x�������cSFK�t�씶��ᙎ
�`�J�#+�	P��"��ӛSc����r��3�Rݔ��UQʪV��r]�3{	gj��yk0:W���\27��v(�ִ+:4��n���m��w2J$,q�E��X�KD�*�
�s(����lZ*�Ȓ9EJ�n�4�e�*�m�����Bm[F���&��(-{���nfe�x�
S���u�qQ�]��,�Q8
��4����b��\��j�b�Zo��ͽk,Z���݌͈V7u��B-����/2�F���Hnh��5���Ő��'�ӭ�i�B��Om�5[30�Q洩k�;��S!¤����鱐nȩ:c^�X�I�7d�{q��M$Y!7��������GE�Q�+h@��1ĕl�nܓ'D�S2�[b�2Zݸ.��jë�f�M�����:�h�Τh�v�7�������vE��n@����11k �e8��f�2��+V��Qҥ�Z�J>L�6_ԖA��#k��Ov����]2n�-KjM�0��ɂnl�M��%$ͬ{� 
�D,��c"������E���--�]��[9!����7�R&� �0�f�q�Է� Ӹހ�6��Y��y�ԭ������ �Vn����j3v��i��T��K5`�ݗ�0�k!lGИZ���ղ�����2�a����+�)+�g>�9�ӫ!�@L��l�lf`wJ
Q��Lu8�V�eX?�ͭ��6�Ykp�b�Q���h�h�pR�Aьސ�ӓ4�n}�Wn
��b�LЪ6�����+]��P��ѽʙ`n���pi�����X�`D�!f*GPڇ5���ks\��f��������Z�PfP���ddKx�Ky��ݳ�BCR��vjh�::i�ܙ�/&�[�#:�)㨦�$Y#R�h�!�Q��up��l%�dM�f��`�r�>�#��h�܆�m#��f	tP��HҚ��������Rb��>C�;�����ʍ�ŧsJ$������sR}&Ʋk[b��X5�m�����DLu�c�I��u%=�o]VԴE"�8�����!��B�mU�	[��5�$�[�5��a��ܗAF*�渆���iᔎ6�.�Pȵ=u���a�s*���9l�.�ei�����yb��2�hS�2h���ח����Gml�U�f(��.�t��x�kUƝ��ol�����N-p9�t�V�%�Wy�<Y�gw[��������U���!�Iv-ҼU�֔KS�d]��J�^ِ�⽃+2�;LUi̺ Sh]5Y��f�gi���tn���a��1�F�6b�Ҽ�j!�V�'7A91��	ǹ5��8�D(�.��6�𝣕r�_XN��Yr�RP�T�-�t�h�"-��D\7`�6o#�׍L��d�p����bU����,Op��aӅ+Q;�׶̳{&��a+�Y��dX�F�7rn,��aԱ�����Xm@m�wo�� ��8qY�e�͇�Kh��B��7W+��Y�$��Jx�x���*��1��`4+L�w%f����lV7�m��(r�*T�r"��hJ�g+u�fv~���r��N�YR�عv�"ưk;wB�Ƣz1k����h��ϓ7>4dӴ���n��d+���j�	���.�����E� ]l�V�j#u���#4c3w�*[N�6"ŗ��t��ۥ�ݽ�tt�a���-_�u���x&��U��dYZZ�����m��MC��R[��B�hmm\�������(�p�&�����8լ�H�69�<�o0#�VYN�	�5h��ɆI�2Pz�m"�KN�p��TI�JD��P��E�l�,=i�5�q�.�F�o#D��<��1R��q���0gNT�̈�ۦ�,j���V:2��E�阷B�U���1�R�c�MB4q�{r�m���ճ&:�c��d0J��2�#�t�xi�u�2�ij�jXɪԔHg�.�	�xpnd�8�r7F$�7�C	�(a{ct��.@�QQ��kڬͥ��5�E�Vo#���6MM�"���wF�l�۰�_ Y�Vm2Y������re�Z�b��ih���q�R�܎������h����r���Q��,UQ����eK�e!�擶��{M�gM#�2H�Zq��cX㬳�����r���<�zޜ�b���Vk�d��J������
��R��:!%Zm�bA÷��I��v^7ٴ����{�ÁI�T5�P3WJ���s��ʖ۫r� �˷��6�B�.�䔲���q��Y(�E<�p��9Z�� Z;/m�sr� Z�ŋbhS'-/xv嗊ѣ P��@��8���JF�\��n�]�E��B��s'Ve�GASSN���c�i�i-+nXƳa��2�(]'����kuk�,3�85rna��z��,�Kl�4k2`C�;@D�K����i�T�B科�DD�cBA�$Y�/-���w��T��z�����x�w��Fa@��-�˂&�!���02b��2�4�&8�l2���j�d�"���M�W�1 I6�i�B
#?&��� H�,�#'��! �,��_&�LIe|҉$Td"�,2�,�Y0DM�fO�ͅ a�	n6��~$�È�??ȑC�� `��LrEb�˻+$���1��!��10v��}�:�.2P¡�c��+qm�X� �J���K6�s��m�
�7ʝ�:���nSo��h�vv:�Jw�ܣ)��Z��b�U�wB�=�cUnA��8e�t�:�'��r�n�d�[N��g6Z͔�3>�r����8dd�}�T���b��W*ˤF�]�,1kW(�붏:�,�yص���#�+q'�r�;�̧J��Y��fb�\����ލ�đg����^7��06�te�%O�r�f��]�����.鸱��W�N���p���
�g.
�34�ܗM�s+8��3��]ivǪ�\��mZ�. ���x�hw~��������]ֽc.��I�4�Y�u۶�뷕$��
�KU�r���Q�ھ�]n��.3|h���������|�|�шl�� ��}����@Y�#hLμ-����"<7q����ݴ5v6�Wt��"+e�G�P_��u�n��oۨ���ahtK��PٷSyfؙ�m��hޱyP� (�=�}QG��<�aA��ws�ۑG.�J\��R�F�2�2��%�2Cv[׀�I�@�,H+�L;�u���/�k'K"�;E;��(򮝾�+���$�r��vO�0Y�@�s;�8���对�]uDؔGh)�d�c�˫#��a_���s.Ӭ7%�}Ԩul/OM��Z˸
V��zo�[s%��&�n�EEC|l���[��v�y�\9΁�7�s	G�Bl	��s{3i�[�b�A0&�?�gLʑŌ��ܼ��#���G�!"��(�L�²]�z3��^�]�rpfKNZ+u����l]���Yt��U;;1�G]����ҹ���j�<����N�5F��R�^�Y��&v��b��5��h�0�p���� ��0��q[�N��bo�I�����
�m�o��%����;�#��Ո��RX��Ńd��]��d�l��Zu	��� �7���I^v��ި+_}�oS1��H'(���I;.h�x\��ͳ�mw�-�j��N�8����J���aݹ���mN�|��� O]l���Ν�b�྾:t���ʘZ�4�B��kY������+)`yD��������.�F@E��)�Y��ݾh(���T���q{X ���3�ǉ��5M�J�Pؗ��uK`t6u�S����{��a\��_����(�cE�;��⹋�k������/������V���]*#�9��Xf��S*� �����6�RQ� �ܕT�O�L
�wR�F5g�+��D�ǻ��s{�8�щӧÓ������b��WWv#0��P�U�|��{�b�M��*ݪ����V�W�M����{ӭ�)����v�����h��w�=N3�-�i`aɯ��S�+Up���0[�G���Pq.&3[*xm�n0�ҬJ�tu�(��ܡ�k@s�OOyH\`x��s��J�S�)^}�V9�{=��l��i	���;�;z�a����C�J���:ob|M>Agy(q���y!���u:�n�o.�#2fR�|��KM�X)���(a�����t���������t0��r�Er�.�]+���Y��rnT����lh��x���Iӳ��1��q�ȕҪ6b�:^y\Mn�T:���K��A�\HӮ�)Q�nZ�T>�J��D��̝���e�V�TQ��y�\�x�Ó;,E�I�X]ê#�`�!�z"b6�ս�Ϫu[�OrZk�*�.0�k]̚�#��s)ˊ\6_@�P���{e�o���L0���At��L��R��km��
o�Uds��ě �#��̉P�XvȋrLeZ*�%_!A�k^�866��\1�j=����T����'��} �/"!� Saj0�����Ѽ�IX�:�}u:`��q��+�f+GS<��J:c�ձ���(+Ɖ��X)p��6�R�f�.UX��2������e�".�ZQ���#|WiN�Ջ}��6c�[!��N�C�E��:�N�]J�yN<V^.d:}�b�>��y��Ρ���u��!5)rN�]��r�0��֣c;^�f�����D��$�c�6K�B5,Ō��1k�n*s��Ynl�	�jYqg�![V��C��m0֝W�����k6ۿXr�ޭ�[��a�th�֜�X�����p���\��R�Pn��]j�7U���J�va9��V"U���Sj��l]u|�e�l9ox[<+��}X�n�q������
��LX�Gø�ę���u���<ĳ#�e�t0A�T}��;٨V8y+H��n�t0����[��\:�]�uw�Ǯᒦ�E�H=f�v����L��n��L�]ֱ{�ui��9Z.���r�Y�3�EQ.��KƆ˩�+�T6�wWU�8`������x�u�2�B�kpӹt���h�]��M���
V�wͶ���۵����lz�̖s�D���0X7��ػ���8�6e��R ��nr}�>a^e4�N=}�<:�ӷ" ��\_@�2�MH�|t�uA>P���u��΢�z��)f���
��D|u���ѷa�7��	`�{5��$z�U��Pn���9�]hg!�Q�5Wf�zi(�0۱ݗ����3M=�s�R���Z�Ri+�؞�cީIp���}�k6���Fe\Vy�q߮�A+K��<v9��S��\�n��O�1婵����o6��B�FH��m�Y��g�/_�X���Ko�m�f��;�wd��ƻo�I�վ�	��5	�={� �b���X�U^���^;���Ց�{A�]��0RH���kRYd9�C�=8h�����2�x���e�",1�9�n��̜۴_K���hl
�.�����+Y�G�fG;��Y����ҽ�:&����UqmU������**��{�jU:*�.�
'�&by������z����F`�}l��[��ܬ*��+�tz���SWJ.���Ig-����kA3�L�1�^'x�xh�'LB>}�\�k�m�%j�r�i%������F�W[�
��ضsz�ƅ�|����s�`���=��o�\=�9Y:����0(`\&���6��h���V�������ŝ��	��)��*bs���gEϞ�N�h�9�F�2+�f9m�x�;�c�#r�o��C]����o������߻�%�R���F��8t.��_c����^�܋0kVR�t��:�od�	d�o�;;�8F]�uJc�����k;%ry�P��MU�N��	c�<cE1�ד7s�٦m$��$�I$�I$�I$�I$�	�&�p҃�A=�&��v&rɔm�R����_նQ��{����$�"��Cv��Çn�X�^�Ѯ�]�����hN3;������Y:{���U$�;2��m�Ź�\]�y�!L���P���gC�`D�K��f}y�r2��A�)i���O�� + L��[��/�fg��� yq4��{O2�C_�q���ϖ-�Pl�0��҄�³vZF��E8��3N)gm��y,����P��/^d����� ��� �C�0l���P����b�$6�-a�z񓐤I7��X��ajkZ%ǵ�:[���oH6���4#�-7)JP�u�)2}�'ƴ�A�릈<M���45P�r!�]�TFDF9�8�[�9�;�}���-��@]��¡mf�Y�=�b,Õ[h[��.��.�5���%�ۡ#\�(�Ֆ����͔��XC{qD)0.�C��R;�O� ����Mq俐ڹY�ڤ.�8�i�r�N�G*�a�(u�l���b���yշIs��"Q!v7.���u;oFR�yʗS�feΚ�Q���ެ�Z&v��9��4�f6Ǝ\t:Ժ�a��]p�UrUP��11��d�ws�j�Zύ��e��n��7)HF�HA�OZ͌L�3,hYdj��K�+7��lc�Q��<.���{A.�:�R�G��M#o#�-��9X�e��u����}Ҍ�V��U���k.���c��2��;��#��	0q���v��≷!�p���P����|��j�FӦIW��T�vVk`�W/J����/e)��F�^٘˨��c:r�Mn�h����D�׌`V��M�teE�`ks(��*i��}��]9�&�U22�����I�g�o��nW0MY6��e?�����?n�S��}�U�|gnGλ�E�o�ē�b�U�/e��6�ɶ�7Fwd�xo;���θ��3y�; ^�Ox2�N�O���μ����l�A:�FuA�꼋����T�:��jBh�&�E��@ʕ��R�����3���][����z�RtH��Qb�'!I*�EM}&�� B�w[T+d���a6n��Xh�Op�۹�{z�V"��gj���T����aф:���q�}���j5� a���̵h-v��踬i�<m�]�'��n��;������Zϴ�JK�j�9�G�\޽Z�_��>���n��Yi�&;�W;�F�r���:䨛q#�yRq����m�^泟w7x�jE�X+>O������w`�hçNEjN,r��'L�-�pq��܃&����0��v!+���n��GYg�a6�w^��q��msy^%�wK��s��ܹ�\�t�ث�UL.)�*僳��e��;�c���"C��r�����{w3��Σ�����1��Rk�R3���ڋ��k�I���uVP����*�]`��/���m��Y�]d9|�܉�z6ȩR�L���mXc#�B��K��շӄ�4���oZĎb��BcYl�e�.�*�[3�P�a&���tǖ��
�;2�bعMa��pB�7\`^����0�nQ�'f�\Lj��,��r�"��7�fB�#n}.�A����S�`ѐ^4q��%V ���fҲN7�ÊrZo��d/����X���c����ō����=/����%y�uԳ�ur,�FN���ZR)���ɥ�D�H��)��)V�G�n8S���(ɭ�:��u�%JpS���᜜��ٵ`�n�z�X+VQ���*YraFfY!�:��v��Ъ0A}�.��t2.�S�TL{��`��M�]ԗ���Po6�lUVw�+����>�>P[w�8�dƳ	�d����¬oѠO�f'�]�c�w�����+�~*�)��3Π���ӳ�+�!�;6'�=���ɖ�P�����.v&)Թ!G�f������V��\����R���xڝ�Q2}�gvI�� ��?J�j��q;����Ze�;�U_Wq2��<�mn�}d��\�K� i��d�Mh�i��<�2_Xѽ$+�� ����e��q��nZ���Lx���P�,��q�7fmk�¡��#gJ�z{�?\����,Q��t�(���D$���Y�ـZ̓釟��1�'� ֹ��ʼ+-:̣ �I�Ɔ�y���'�ۋ{xm �J)ѭ��������:gwjw�{rW�#o��tu�b�Q��=6�
��V��/��o�|���g;w�\����Wf�]�,J��x-��ߩ1�'�����p! �Z����[XA��7h!®�M7; �
���O�հ)��-�T����gk_��p���[���5yS�j�b�����Ԭ�)�:���`����3���_K�5MjJ��k4,6�
ܭtnړ� ��Q��|i�ϲuu�}U����;�ܓ𤋮���N��b�)��O�J���,��Ԫ�ڙ %�`�HkS�*�>�Tbn*�����g��(�cZ ooym�m˜��VJQ��vӹ���mz	�#>�<r�T���)u�\9
���f0Q�/�b(��O*���7��5�:.��Q��?V�_v�Y>��q/�_Z\�j�_;���ʥ�T��K����[|X��*�۝`3�K�{I�Qz�=m�F��-����k����wg�:�f�����l=t��x�\��/�HM' �o����{nQ�Gw[��|���x�G���;�N�螺M����x�.���cW����q(����<&��e�<����J�����f����������\5��,k5����� ��X�	*�k�7V���XQ�%U��hŷ�b\)�˦�Z]�(j�����_Bfv�՘"Lح�Nn3׏-@�N�n��	�zx��-}-WJ�[%�w:��/�SM���>ϐ�:�n�M����jX��_r�@0�]��n(��x��(�>e:�M�!X��'u�[��-tk��xb��]C8h�,ca��%��}b�O�&�`ձ)��/N��J��A4��@��;f�_����i$�mm����C��L��wv�93�w|�l�Xw��Ս�U �h�����s2�w���(k5��P��r+O%V��FK+��UL�'+ש�.
Z#Ŭ�fmI���.�WvU�gfm�i�gM�N�&�Q�]�F�c�̬��+]����΅Z��t%l�Z��ۮsR�qQcm��C��S+�.?Z�1U���c����MS�H�LN�Y���ʎ���naͻ��wP��Fmeo$����d��٤3S�'i�&W-�r��H�\��j�s��AޮJ�����
ҕ4X
��)c��u��p�>ϕ�Q`Ixkh�`,]ޥm��tViW3��j!��<��)�����7Iҡl�а��:�}���^ƛ�LX.�
i�Z����s̵|�9��zz.�����\�+7�J��R�F�r��r��u,cdul�݌Z*��'�����J橮c5+c6��r�$jCX�3j+�6��Ψx�ƽ�sl�_Ms�sWK����"A�"����+��}l�� :��]=9�#,�(�N��8.9!K''�y
��Ò�W4���-̱Wvۼ���a���59��)��KH�3P���w������̼� �8��3fч�aܙC5(�!k7u������9-"M�=��,�F��WI"��	!+��nB���6ܸ�H~�eF� ��ss���#n���k�7K��)FV�9*v���rp}[LS�.�}E���u�9s3H�p�t�YTd;xx����}�/)k:��V���F.��L5	�G�u���v8`���q�T��x�͇s�a{�B�a�T�YJwMf���S��w���#n��;�T�ȉ������Ψ.l)1��t�����ms��{��GU������v��K�;ΗH�f�Z���l���ͪ�CS�/n�}f���V+[�gq�#c8)w�&u:WW�^��z�+ꯪ߯[j���P��k�]���ڿ�~
��P@RL�a�'�B1��� /�$4c�?� 싻��(�b18�!i�D�SI"e}�����F�v+Lj�W�#0IS�p܊�7�Z6v��u�/���^;��ߜٰ�A�Z%��(���t�N�� Q�V*�V"�w0L�bv���o�<�5�OiJ��M�w����KTJVU�ϳ_2�H�:�dܠ�vu�s������p�6^��v��PtS\t��48��n����A;���S�D����l�gS�F�EO�]c^f�Sh�V*��̭H ��.� 	TZ�� �pJ2J��q�^΅�k�B�J̼�O"t�-�
��E�OVc7Ʀ�j��l���|�@N�}�~����׿}�ͯ��Ƶ�V��V�5|��m|5�m�o��-z[�;^��lk���:��.MJM�$�I&^���D��2��FђM%/}]�/<�*4��ѵ�Ɇ�Jko��·J��H��o:�X�I�e$W�n��U2ƍ�@��Й�CZJ�׿:�(�űh�m�Kd�ޖ�b�*��5��66KF�%���Jg��z������ؽ5�"�,ɦ��FX�TmE3HbL��;������x��[�W�#� ��Hx����%��ݘɒ���V�
6n<��(Z�j����{���I��p��*�^����,>-�a*����.�P�´lf�e�����������eHǵ�6�}�<穔��+p��s/�7kWu�ฟ1{�;���{���}�/s�ȭI�S�����}F�|��Y��9�U*��>��������ϔ�^���L��1�n��P��VP�w���`��W�ۿN9+EN.�~[H�5�ͻsa���;�[�����E�=0��`	U9�Y�9mG�״�ߘ��"��>u�NJ�4\��ۣ�%�@�5�ط^��%J�Ѣv�S�(+=��Y]xd�A1�T�j��L�d��"��ꌣ�ے�bz���|�ԃ̢i�r2�������.I/u%�'�t��]Ud޿�Ѯ��+'��g�>�V�u$�}_z����n�++Eޞ�t��_N��ٰ�	"��S{ǣ��g{��Ky���3j :��8�kel6��,���X�ڣ�i7.����Vb�R,�y�͵O������rWV�N��a[��V��?T�>�ך��ɝ���d�t�<��I��5�p���N��ww1�����xk>S�G;O	��RN�ł���^�`^*���69رd�[�"��l�+ۇ:;��sVo���3����,&��`-�����$���P �u����k�i
�������-JF���j�x�;�s>�1��u�:�h-se�u��<���6M1W��s���df;l�Yj�f��7���(��݋�[]�Js���7�g�P�L��c-����o����<��c��L�������3�{��?x���b�*o[�u���w$D�F{~t�?d\͞>8����:y��1Ə+�6�Hς��\k��0c���U;���L+QFn%�y\�;m�����<���c���h�'���Aw��R����d��J��|�w��6���wW���8vX�l�����}&�T�B��wf����&���)t_�����A�2�fn��m���Oi��]��۸�Wja��W�t�|����f�*£�.�w�����6���)Tr�Ϭ���mvۥ�w��mjP��� :~:���Ma��*c5j߽�%/>aIiU���]���,�9�[��xx�x�}8WI��6�r��Y)�΢ye׊�r���xǇ����Y���?�S��xh��A�|M�|دn���Wf�O��Ь^6�w��-�a6�"��0�AJr�U	΃�BC-Qu�������-QH�7�1�Fj���x���/��Q��5�{�Q_
�sJ��>��/�>����>[�<��C>�
�{�rp�?d�����yW�k�g*^��a��\���G��}�z�-޿t�׾�1�U�s��bz�|H��L�nΘM�զ���S[�c�s��k)���[�yPF/M����S8W��) )�(滂�l��̺P#'tNc��"�z��uo1&\g�t�|�Vg{mXX[qJ�I�$ƻ
3Y�j梫}Y{���7%��Y�N�Z�77Qml���m�����S"Ю����=�j��ǔ�f[�;���k��Չ(��]���?^{m��y���Ю{��Q5s���u:��
v�m�6��*�w*�U�0���~��V%z��(��~�:����f��Pl���oݛ�(W�����^M��b���Z_{�I�v�yo�ͽ<6/�kߖ��m
i[�]�<5��,�\m�n/�R��s�
I��m�;.Ǹ�(h3��4��y�}�c]�s�o�uy�*4Ϳ��>���g��6�%�}]hY�wC�����y�<��'Rm��.��q��Ofu��-�f�_�́d9e{�v1����7s�w�E*e���ϴ�:n�w9��J���ᵀ�^z+L����,��|9�����O������Q�:�y��e���c7Υmuv��u��L	g���K�z�(4���])�](A��qҜ�e���n���G�]Б����2���҅t9[��px*�)���,���Ƿ;�W{2�!)	�����������S�L���+�L/n6����U�kxEM������)Q����g6%e� ջ�ߋ^��L�qu��^Yޞp%��o˾�w;��<�즚��ˬ�p.Jbr�9�kM{~{�^�z�z����F�������F.�}N#��xfPh#��[*�짛A�;EY�/�vۦ⽨E�i�� Q��K�ٽ�䚺��{X�ݨ@���8ة�02K�a��l�V�I��;y/y��zeW*9Ia�����|Fe�^e�g�@i��^���b�|�G�Ӄۯ��؝��
�0=Z�l���:(]!��/Y�>���;����<jw���ف�i)��d��K��z��X���3�߅9GN��WW�hV�M#څE�%��B�wA�2ٹΕy�����p�ϰ�eү��L��R}+pM�kǙ��N�U���{���'�(�^���kX�>��>����>�<�}���)�&˝�k(u�r�Z\�H�zxmA���w�W��,N��h=q�|�����%-��������f����Pꚧ�����b�D�j."����u�Z��G���;��͵!����q�X�.��T�����U�>�m����;u��Ju�Rc=�8n��~��<����.���~�f����ul�����<�3r��~{٬�^��a�3��Q�s+g�Ŝ���nL����k��������p캻�LS=�������wg>;�aE���+����}��N�'�F���Ʋ�9���ll�֚T�n4P�Ѹ+b�ۥ>h���o.�1Rڣ����,҅W��@��/:M2�W��z�����i�+��*��i�UK�<ƻ����-��U�ech�fû�0�s���{S�96=	3�C[��M���OT��tt�\��/[{;�~��5oS*_���e_I]+�f��חd(^�A�.�ϧo�y���紳Խ�4����6
�!�Cʹ�J�0j��D!y[���S���B���{�O->�x����U���;�V4O[[�n*2i�^L�V����c�.�L�d�ڊ{�>�7U�@�J�v\c�-�W����=j��4�kٶ��+��|�z�ư[�]�m���A��f����i��!"x-�����9�o�o�o<Pٺ3� ��_ �v�Ob�X�(X�\�X˭�i3��5���Y�ޒv�e�V���5ZB3ƶ����;�Yck�,�2�W`�G�aϰT譐{+f���6+�g�	�0`�C{V�*�O�8���������g,�;���5S����QK����Yˮ�zfܱt8�u�ht��HC0w&��dVM��:q�����Y(�9���%@���Ae�{�����p�1R�1���L��t��Xq����twC�[a]��Ս�t����醪�t�Q��m\	i���s�1�<Y&@X0�h�JVX�]��	v����ƴР�qou0ȫַD����E����Es����f�E0kǕW(�7�PB)OmIC��G����޷[s���y�u�����-��^�*Н5x^;�Pu1���e���Z,d�#��9�ĭ
�m��lю�ܶ.�i(ob�DL�'ΉLT�N�U9x�AaH���3rV+Y� :�k4�ȺG{�W��2�%�����̻��Ņ$��bʚ���kr�Z�g�C��`��Dκ<�e,�P� U�����"����T�g3{np1�]%�v���C/��a��R��C�]��s,Hn�����p���6y����YI��β3��Wte�x�2���ѽdYl��/ N�wb��WfuݫJ�M��C����{S���ͩ4�w�Tb]ձ鹳WͻM.rknBi�[��(d,�K�J�)Ց�,�{y&�"+�QS���f���M�?����~����fK��51痟t`�y�e4l	�$�zKwp�+���ͷ�ܨ����ܽ=<���,VM{nm��ܷ5̛����Z��%����.��]/J�E�71O}W����W��׎li�/:�m���o�sQ�]��Wy��xۥ����|{�5U�M��1���hzi��g��?����9�Ȱj/'�+j11�r����]]-N�}̪�e���{�r��������-w��s<c]�=�����m[O>��+.w�c�m�͝�3��|���Ϊ˸f^R�eHV2���x���@M''_�Wj�>���@K����X5�uϽ��3T�G��58z޹�la��=���|j�shn�g.��O���<�Ȍʝ�ʋ��w��p�6)�6��9-4��赗U�kD���O��%˓���%�>���ޗ�u�2��0oJ|z��A�%�1;������sQ��6:KN�mJ�^�j�l�J�+�����:�f��(�D��CNV��w�e��v:����+�����i�|����Ȱ�M�6��>�ᬷ^i</�{/����1�y����F�o6����`��Q�v�+��p��t��`�y.�V4e�fD�Y��K-J-h�?T���Z�u�ZڪI�9�W햏�)ʓ[|�~��a���5;q�w�ό�[��T��k�rm��hei��L�������w�rA_�;���W���s{(�Y��w�{_U�MQM�]q}��oc��/���EK�z�4��q���s��yן�?�C��x8�E�`֧x6�iJ�O곁��6T�:CO[�U���gO�����"Q`C��~�����������{,A�Oy����((^s�����bg궝Q����� ֓�N^{
�{ti��Oq�~���|�R��Rw`k��'���ͮhεLϯ:!�<h�����s�]F��*�v{[i��{0�<nMD�Xrs7^b����с�����K-�Z�]�i��3��}WP�4���ݘ}���y��W2��H�ݻ�s��vp��wy�KZ��Y��͢���vfvlӧ�M�Y�s�I��C�n�k����̇��y�i���g_�mL��I�s�"���{�;���gh��o%��'Q�P���+�mf���W�smu+�$��ooY������:pϫ�}�{�6�m&��5����-����� �rs75��y��F��]0�a�n�oDS��ٸ�/U��-���_<=��P60k�Ŧ��]Y���9�w0,�ӳ��{��:�d����sxD{K�	�C^9l��wL-��|�%��	ν�a�14�V��5�.�m�疾���\���*j?�qfRʄ��xx�҆t;[�kOZ落~[��؟I�Y_��R[�O=[��a�1�/k%*�S����43��cʤ	�p�>��b��k�F�c�ƒt;k�����S����V^/ �S���G�����oQS������<2�^K�y�k�̷xe*�|�L�� V�\������_����E���OgT��unD^�V�jt3�T^Ƕ��o`Pе�~������Gz��'��g�%�~:����/h��K�[WU�1~&���{�5Z�����Ţ�{�=�f��?x-[~����w��"�2���m���8������fw'���7�3�Ų>����h�7x!�q��9X��AX<�� ��ִB$Urh8�"ޭ㛡�;%�44�͕yijɄ�}%�����q���������f�y����-/��[ ��ݿk�b�QH9$A�[�3O&T���`6�߬�N_9N��pGձ���x��0ؖ�xxy��*��G��|�Ʒ��x��O_R���:�g\��di������:O11]�S�&`td��R���N_�`	��y�DZ�ɽX7��<���M�U�`��M�����V]�j�(;E�[Z��#!H�+C�Y��p>hn��������?ZoW���z�����?w{��n��P�"�[�㍍�~���?D��߬�ݧ?N�������8߯�����n��g�ʉ��4�qV��qy�����c�t�Pܮ���W�y�30�".
���t�SU�t��<����eU�rQa��WR@e���0Ű���O��E�?W=״"ݿ'�s���B���1D���iL������ �I#�M���ļ[R��v3��r�7�U��d�]e���)4�S$�ϕ�&��� �Ct�k��ʮa]�f)��+��Lne4^<��.﹵|�iQ�9�P����XUܯ����!6��L�sy�m�vW4UGgG;�t��:�r��E�4\B��q�v�Z��F]�8Z�8��n�j΃;�v�6�P��+9۱����W�WN[�K$m���|����f<h��F���M�SO[�p�/a�:c�1��޲�2�R�f��w{_�T̲�Z���R����:d��p�G�+z~����7�=t['홲F@K�G�mi(�*���������y�Y��_�Q��H�x�{J52�q�~�џ��?��ԡ�V��k��g��k���Vg�q�ӛn�:aoX�W8�.2:�KD)hQ��y�}�����n���K������"%5#kow�M����S��R��{���[þ\��[�f�ǆ�V�HWN+����{���LKtu�vJ�+ʹ�R�����>^#�دo�)W��Ͻ��p�\�3m��F�]����_J��"k7%�oh}�:�5s]�l�]���2��3�u������rް��f�#��P�U�n1T��M�����Ygđ2�V�2�k}�uQv�mGl����<m7��S,�58�ǬX�?����f/1<Ltwxӽ�}�1�[f�s;�mp;jgm����p��&~�~��#�}�,#����vT6��m�u4��Q�̡73Ud��N�?lk���?�k�D5�XW[��!�����?���>�)��u��v�kگ���E�ۑ�MwH���ٽ ����Xz�q��~�
�kI���s���s�f�����{����+��hYz��<8�(�}=��tw<��h��{����%W���{����}��!�|�3jW�~I�f�'��ʻ�<�U����%�HbNͯ�yu�2�_�51���-8t׳Bh�T��M�ʹP���x{����n��߃�N:97x��f��Ih3����a���e��}U�r�'7ՕNnz����Ѳ�����<�8���-B1��}��VSghP���<����C	����e�VQ��u[���ꢧ���/�5/ĴZ����;�s{Q)a~������=�C�qjSf{�#j[. ���_���DB��X-�^CL�wK�Ou��Bކ}��饏"m��+��p�؁����]І5;�յ\�mkۡ�N�%��ǈ�����X^�?x���Ԇ#e���
jD�	���	�Ġ���(`�
�����D�k��!��H��2��63:͔�.����� f,e��|d�|�!��j�y]���{&�D:$L��5�"�t�[;O������}�p!�����P{|+�1�#��rr�|s��8�ġ�������k��8�i}
鯅Z�P�,�b�0(߲�\u��	!���Ů8�ܘ�z�II��å��λZ\����*�[55��M�<�f#W7����a���R�I��j��Q{��C�]�dB���/m����
s��b"X��V��S��a:��9�C��������]��W� p����B�d2+[IWZM��X��n��y�"��.��UoC��94��Y��D�@�*ޭ���<��-���}IZZ���R	�a�Q5��G��뺸��פh"ĐF!���-@Q�b-�������=�~W�l2Z7Գ�I�62Ԗ��R�\#��R�;�V{Q*{B��E�vw�6��G��:��N��5@�C^��J�G$S,X�q˥H>���L�(L� e�].x%L{����P1I�6��h�dC"��.jA��:Tv4��UDY	�ҭ� �m;]4�+Ç,f�h�O��TT��6Ś�r����ܛ_w�) w��N���8!l�s�tR��N�"�*�r����VZ�����1�,c�eF��8���C5�7�ki��t�"��vO�m	f�Uŋ/��Wi1f]���mvj�<$}{,$VTcǍ�ǀ!����uI��F5�'A���{�f�4���1�uZ�Yzjڌ�5Z������W��-�ۘ�wv�Wu~�m�����H����v��^-�%�!�kpM;����qF�[���:��7���m�ם�=x��K�)���:� ��J9��P�����E�1'��'�������	^����-Ƚ/
x�nXɒL���ۜ�.���u����F?���?��5�nV-�̈*�O?���	a��K5Cc�C%�Х�ĕ�����=�a'*�[��̙��"�z������!�ڦ36��S�l��.��<7f0�7���_����	M����Z�6�E���f�L���	�>�OߦoG1*B�5ê�Ǽ}���~v�"a��ʁ�z4����������\	���3��{�6���(��nyG3�}k�J��_��?���3?-�jY�G�t�|�섪k��W:9����r�V5��X��ƴ9�bi���2��X+���S�M�q�����̒��~�#��.~����*�%�c{x�"}�ղNgf��P-���L�\���Ɲ�(ɱq���I��l0Z���K=O�(�m%�O���  �_n�=�ɻ���%E��'�GKz�)�k�f�i�d����ճ���+�t�Ws/��P�UZ�՛��T���^�����b�Գ׬PV��gC�UCu�T4gE�d��Q�h~�=��혳g�R��&~��&� �l�~팑�x�u�`6�����΍�BOD�f[*ꋌ��*f1�vwZ������Ejˎ�BLl\`�n�U��x��=6�_��Σ���g��FJ��9�p�*�^T{*����OL����	/M�.���ם{0۸�9�hJgk	m�3y[�#�]lG�nVV6^.֐�Tm)M�'"ߝR�8G����L�W��R3��ڝ[=V���3Eߩ�f��9��l�|�OyK'�ٶ�F�vL|�uwd�ŵn�O�8|Ю��~؝�G���f�z�)I��Ñ�b�|չ�oh_j�g{��.[�TLk��3w�'4;��t�OϞ���
�۲�P�=J���d7,�hV�@Pb�Y1je���N�#Y��vU�T���@@��p��	
��4���k��~�}ˮ�^D���W�����Ԇ�k��K���]�������a{���ݼ�����;�vi��5���Mw>�whM��q����],�Iu�Ҋ�V��x��9n���/��֣��Ƃ��t���UU_<��3i�O��ǽ�y9?f3�q��nR�iYɤǒǧ��(�(�����S��H�u�(EK�]M�Γi[�9ʿb�=�{�6���ߎӝ�?u�t�"�-
���3N~����by]=7gچ�3q�iR{��v�Δ����ᆚ�Ωlut�Ԏ;\I��5N�qS�Uh.5����V���#��jUG�ezy�yC�f�e��3z&a�����P3�n�D��e�)i-���2ΨΉj w�����v��~�[�8��G
'�y���3L����4��7(��7R�nW��f�吢-�Bn�*Di0j\�d���9HM��#�{����K���*I�uY
6}����"36�՜�ݍ�׹4�l�L��nQrv7*)J�f��ǫ�Z���@�K���.+��S*	���M��QqI�>�X�nܺ�3	mQ�dX�p6��&{9��
�6��ԵY�e�bcm��D��fbU��T%�<�E���b;��gߺ�2��K3��}�<���.��騽�P(UԊ��u���Ž򷽶�Uج3`/�݊h����a��{��!�A_&�gΌ�g�nw���̋�K�`J�3#y�0�0܃�C�l�(Û�Q|S��;\����p�p��l�wѹ\���A�Ӥ����onN�]0�ջәEUfCA��X������g������3�&;���n����p����ov۶#O:�w�bcO91��X���x�}ܺ�=\�;m�-��|M�����錪Uג��������971�Mږ���.Ϸ�%?z5�n1�w���c�`~}����d�)nR�7c�6�6XWr���6�ҿӻ;��mM���Ҕ��j]|�2��~Re�Dϳӽ�`����aJ��=�ǽYO��][�6b�V׉{_��"�4~�{�m����ة�����:1�y�n�� �/8�QT�#��m�X_���o#�K�6��e���T<[�Aٚ��u�Rvb_1�5������ۦ��W��֭�7����I�����X<|.^�9`�s��]M���M���
 Jk��܊{�Ʒ8
�A5�|yK'9y���R�OTSd�]K(	��Z�<A�ښ�ه����P:e�1��a��W|����B��5)o�{�@=���l�����ͷ]�"Lv�yy��Į�	�\Qܖǜ��p"�[3\��a��<�U$�x<����^n%Eڨ&c-����'�����}p�m$1tf�;[
��{/YKD/W�X	fQ�zœ/$�쵕ͽ�'&��X�P�B]���.HzҾ���9��nl76���:q������L�P����a��0���=g>ݝfF�#�~/#3k!�ذR©���h{y g�����������y(��)�{Q4�8�,h�<�<~�ڬWR5���Ş�X�~3ַr�9.��d�)��I�u��(��7J�m�Oe]�5�'�q�i��M:��J�_Q\�5`�OɆ�Y�{y\+;�ѹ]��F�m������Ȑ!6�3$��٫L.wkUw�R�7��1Y�ؼU[��'��A�ȭ��3����;�H��������L��2�\�Y�x��߮��g�;h��q�+�1d2�ФH���Au��h�v�T���s��-�\a\,:���I��-�)>{��U�b��7���n���7,��M5��3VVv7<����d�/%���sGC��ai��)������0�ۤ#���ah����Y��O�����d�M��v����m6�vvE�h�,/��1��q��k?e�t���|]�LIV.c���D+���3�u���m��`B5!^|1wz�S���Ll�{��=�6��M�ι�8%Y�Ȯ�՘�b�k������}��up�U�b�5��]C�S��ָ�B+�E;����2Ţ/b5vb:��/�L�ԢM�C�����c���B���D�ѝ�%��E��^��wc�k�.Kf� C��q��u�0��M�>�}0��7J#�n͇w�̯K�S�7eu&���M��ѢW/�s��$�����=�Z�Ck��g���O�<�����ҕ�a�Xk��
]���z��w5�-�z���2 �D>;%x�����q�/�V?I+˹Q��4��f��+�m}4`�\(���.wk��Do�����S�M��~=n7
�	�:ǚ�����Owd�Zw��Y#��G�?����U 3�����z�K�m{�fi��7�W��8���kD�4r�7�(�9T������TE��"��e��Y%1����b�Q3gv]�Zmws�-F]�b'�!w�6Խgi�nI�h�������+���K�L8�JY9,��_E�VV��ޖ3r��h�C!� a��t3�L��' �Z�4��8��v��P���>
�/l^�I{��5�B��/��E.�Y}��XV;��0���N�/.b�һ˓����ݒ�(�5��wV�LN�4�S��g�����B4W^5V1H���8�C�x[w�eu�܀��K����o+A�J����".�ú:�G09K��,
�o�)ɖV��0��&��K=�� ���a�OY4�fj�5�4�L�!Ɯ��	�w98��� �
��罶� ����v(��;���J�LOe�߈V��V��F���aId[�"��x�ݹ���!V:��s<u!R&DZ��x��8��f���%��d������r��o_Ԯ�UF죑Jd�w�"�T�e������P`5����ۑ
�"c'p���<Uu���A��9�^t��G�Ȯ�|�u?F��Yp^*��}n�I�I@CØ��U`O*��m�
�ń,��&�F�N��۳e�8��n���Wk�G@k�"����.Q�uI��vɖ���>Έݽw����s��������{�{�Ć{�w�܎\ ��ﮘ�H���r��Dm�c(J{\�����Db�����X���4�$�	2�I4��ѥ�u�\دS�{Q��^w&0$�3!(̌I2!��Ώ;��Z jf�p�	&o�O�-ƞRo���te����Ǹ)oۚa��s�e}OV���S?������d�hq��o\X0_V_s�go�/6s�ظ�ɷ��e�F0���V��I</�W싾a9^�9��iM,p)-���ms�Ջ̇�Z��R��5?f#UCtk��(���o=��Ʌn�#n�/so˶����4P��v��-*M����䢣����Z����>��mc��U#4��jh�W� b[:�
���-t��,x��гʃ���4]�f1m0u�[�!�ћ�*1�g)�#�z] Cz{1��?�n=�F�*�V����Z�����R���T;)��ގ�%l���T=y��Ƿ؅J@ӌ����]v��2s~��M��y`��0��gU{�����Dy7{b+lOc���f����>�@S�U��-�M���G56<�����q+xj��_�@�6��Ed�̛��;z"s<(c �>��ɰeM�Vr~�������r�����_��#��T�M����$�+�d����L�%����w"��(k&[S�}"g�B��&��/�P�~��]i��q��.��}�aއ�y�R\�2G>��/en��B���~KՖo7X?g��~=K,��N	q.ͽ���]E���O�:���N�K{�c�aY��g�d_K�9�l���4U�t�Wo!W'\{]Q��y˅�iJ=�՝��Wc1��O�s���_z"���'�(��>��w�]WK�!"b!�)�����+Sc��מ{7|Zy�u��5��mKLUv�\`����O�;ѓ�w�#�&��u[���F����
�)�����UՓ1��������&�D<�z��뽎^��!�/5@k�z�c;���5�Z�̀����t�H���|�Qb�fg)�|�T�������GV�;eV���g�|������� ��j̘�����(�ǭ@�I�!�w -e6�f��� �|�[�#_��T&X�b��<퉣*g���(hcO���wn�b�u�W����~5���_�d#��uOM��2�~����J'߻;��f_-�L�����ҵ�˽T�ڭ�G/9O��_"�������dK��<�st%ldHՕ��.����]�+Ɋ�L�OQ����,Q��h{��Uؐ�x,ɧ]]����W�/Z7���|������\��C���V����g-��g� �?��@n9�pN��If�K"��_�B�L��v/m<��ݯ߰�!�:������7F��V�����/.���2���Ǫ�K����W��8mkaت�I+����W�R�}gI�"��LVkm⪜�f��sC���z�i�����f�  ��J]��0&m=T�"qe���.v�8�ƤSH̳��T��[�����O��W�_��� �`���sE� ~�g~^[�vжL��~�w��cHRN��HȨ{p��(�w��3��(4ť]�7V��lq��7v���,a�l�vR����ؿy'���/�S�K-�69q�h������"b�P�pj�9 �[�[?*�V�H'q��O��Wњ�c"8���\�;�Go�>0����f��8��'c|���z��-�I���?~/L���G:��}/:���G�ﵚV1+)KX"�.t��6YYv�q�;���/��k�xQ�#*�����7��X���\{l0�T���OyQ�+��o='��Za��_���ֲ�T��o�T<tr;�=��*=��F65��K���6<��\�q��UG��g�k���c��t��*Sǝ�Fmc፨��ov`AeA���8xUb��=�ç�~�t�M��3K�\�����;(˨������nڏO5L6\i;���C��\���L�f{3���&���O��!y.��Y���U�r�MVݨqd��>�M�����cZo2zf*����"��h>�2��\`ٳUC%���K[��y�.�7���j`:���_)��is��
�_I�Kz<B��p��H��۬x�"��o=��yY����-â�v4|�|���r�_׊j48�懑��$��;�mK٦(hy�����1�JO;���}�l^��W߄�s6~F��-���f7����)Ňs�Q[��t?�"��>�A坕X�B}μ�}��G.g�v�s��Z�s-�b��num4V�T�#����,����n�<�c}�_��O]`y�{I�����Y��N�eA�v�h�imzUt�qC��Mlz�4�����И������q��
V����ں��gw<n�%��DuYUu��Rs��66v���� F^I�u��O�w!���^4�b�m*�W����3%AZ)a}n;Tz��7��'/�܆3��k����[1Z�	�{Y%���V�#|�P&t�ca���2��b,0�Mv5��zzg�%*���X� ���ЖΌ����g7	
���	#h�?.�a+���6DS�ד����y=s盵.M�џf�W��?[T[	��k뛯VK���qYo�Wc�C��kW��fߙ�W�c)U�Ϊ�P�2vD˦�OZ�&��f�10C�a��8�j�)�g�����`Sb�w3���qm�J��G��d���\yi�h������:�k��z�*����7���KT���Q�0kS��]��l�ы�,�ycmo�/}�
���iQY��ei���N7��j�[ѣj�7�.R�O�Qo�櫢b=]�c�c��*Z�ڐ�9n�EF�m���'��l�;lT&-�9�¨�ýw�ӁӴ��9qw��'�dNn�q��E�Mw������]�)ň��=Y��"��L%د�G�4a+g�V��HS
���5'��J�!�F*�#�n6e��dI��C��IE�cL�Z"YC̩�]�����d�e7
�͹���^���B��N��密J�K�gT�4WK���{�8�M�ZJ��gf�U��-���i�$l}7[��.4�4���)RU{�![��R30�D��?7<3��fu�qW�!t�{?<^��.xwɪP�G-P��T��;*v'�|��[)�u}���w��t��؁��D����B�=�vc�ѕ���*������!���][�[���|�r��p��7F�������{���zw}��eI=�y����	�μ�m]\�vn�:7(��*����^���n�XDq�>��8ɮ bw������:l��b�B0Pm�	�	���,%�Q�HuVG�����k�|i�U2���Sw9]�#*T(�<p�������@�Qm��9Vn��r[I��B�j�i��(�5��c)H���t�)u�7+f��#���Qӣ·m�WKa�#��+�h�S���ޟdVbP�Y��Ns\��\ƻ$f��/lUB:eJ=,ٽʰ����(-7��q�m�Vb��W^������j����u���q3�:���h[�������W���cF�����:%:h��{������A�J��^K��NnmX̻�#�@�y�\�tR��U'�g*���T����Q�����P�?1�zp�TVX�H�ƬU�Av���nmDw�r��b��p}�NIQ�=�A��3W�g^i�ہ^�a�9u�-���W�a�n�
��̢x����~`��6[D�)$##?O�a�I,��8���{���r��5�#����:��2�=���GEJ���ۆ�9%����mb��=����m���V�p��쩺�"����]mQ��e�*�2E�[�s�.��І�Sym�䩻\�.;��-Q����/l���S�v8i��ԥ�	�X�]Y8l09� �w�����t��#�#�V��B ���u4��2�ʝW�l��8y��бs�c-����ږ1S�K7�����%7��ͷ�/�N�/XDc�]K;J���V=��ʉ�Es�ӻ%>���2$�y���Mh�A��_�T7���V�X��N+r�ڈ��g�5�:���V��.��t�&���S�<-����t{n_�h���5�;�Gf�}�{��M]7�hwuI�z������ ���F�#v��7>>���]�ϯ�z����0C4�)�;�)>~����(g���\�ey�L��K$0Q$MΞwTL2Lu�a�2�]�H�hIKx܄�F�Nsw�����]D��$�(۝��E��d`�vlb(M|�����}x�ޝ�;��|���~���2�͏���s�`M��9�� ��nHek3�؆�bvgr��~>运�׋T�gg�#�s���\�Tj;F���
��-~��훾��
d�9�W���*��OnEiY�ϻpY,:۷�B�f����)��Ѽ~��w�٭W�eȞ��YfE�����
f�U�R��VG\�!;a]!�1�ל��&��d)�×X��M�7=zAᵎ�&��ʄ�OU!R�/ [�秈�����vj�y'�8��n;���D6�=�\���*��j����|�/t�e��Y���F��NQ��֮����\�ۛ���1���R�t�c��-�D�
�Y|�	�m�Y����c��vv�ʝ���`��j�4�5��?���~3��o�+VS(��rٌ��\{��@�n�\u�ӿR�;������[i�",���ȴQ�i���뮣류f#�^�e�G;p3Qh[8�|=N s�������xםD�T.>+z�t:ۗ|w*���B��\�C������{���;��2����x'u��u��t���=�����x�۩d�+ƫ7ՀuxT"��/��:\g�?�^��ۛ��_>㛌̄�^N؛H�/pi븛v��U'���ęsmX��x�������I�T�L(�E�ꛝLq�#��]��9Å�>G�%��y��X#4�n{�d���p�WQܻ�
��3�z���ԧ6�L�/��P+9v�x��~���m���k�Df��ٮ����c-��q7�j���p�-��f�e��:�۽OQ�};t��U���w,7��y����<DzC�ći��e�j�<�µ��yp<�W�?����(���)�q}0��������܀@o�p�EV!l�ζ-������t�ڮ^��nqj<0�S�W����f������P��_���b�ѿv3�^�ߢ���O:����B3�G]�Xi{�R������X�~u��=J���t8��}�l�"��b�;n:�*[ܮ��K�*	�]i�ȡ�31�w0���mn�|n��E�d�Wm��wq��]�9�{���p׼�S��u9P�����MQOz�h��\��|��V�ݤ�I]��9 �%Kd�'����bhɜ�ʗ�Ч�5�R��=�a�L��y^���4����a�n~�گ��wmU�]_:��nr�fl�ř\Q�r
k�N�����@��xy<_�m~���|�Y��R,1crF/�T�E]�Q0��Q��F��_�b,�^���z��{�O������{!��`H�eM� �;j���*~��
w�r�B��Ն��3&��6��'ޯ{�	#�����f,���@��\Öcd�]D��b�&"q��b>I�9,��Q���c�?uŜWu)�Et�xkU�����ڪ��(7Ê4� ��y�$�')��6E�US�1:׮�+�����mi��u<S�lv�0��{;^�w��?��-���$Zfb��E�ȪԶo^�5˴v����6%�֫��Y�S�;��Q��n�[�����z�v�e��S�!�4a�6^es�o.���UZc�Ra�]5�qH	�e��؆V�Q=����u?jڨg�۾��pU�ҷ�
�SO���0�6�ři[/�f�q1ll̼�S{hwX
U����/)V齻3���-�9@�MN�������2�Tk�yʍ%癟���Yɟ��P�����ca-s�rz�T��W]��0���k'9���h�W'�ǖ��h�q�z�+*��j�|��~ �l��g�y���i����o���]�^�d�x}�w��r��܎��f��v��ת�0����<KgC���O���Ι~R:�����i9�:]�F�����B�j�o���.���|���������]�S��6���AÊ�J�ꝉZ�R���[z�ג�[u�X�󉁰R��`���ľ*��<M0R�Z��7nl��}jV�m�r,_i3me=�'m�5�s�t�J$���ć�I<�����}����������?bZ�(����L���`�u�E�2��5�o'{gl��mY�@��_#�n��Q�-��ԫ�;{wY�{�Y�%oJ�����1�Y��3*1���CI��B�z��+{B���1���o���J��ĻW~F�;���ѱ{�=e!;U��m�)Lh�����m9��W���yw�[W�aW����8��mP��z��]^�U�Ľ̼�x׿^�~���m����C]����X��:��sr��og>ւ|�M(�#��k˥F��˔�f������xr����ݗ���y�p�Ǽ�>��)w����	��?N��a�^���ف�1���^}i�k�Ϯ
N��u�F2��r�H�3��ؾ|6���'ƽ������u��1�/���vr��Ͷ��n��@N�Y��}VYφg^K�Y�3ϴ��U�==����NNelϛZ�Lo�Yi�."&�Gjp�n��:ީ�/z�w+Um��ˌ�����aan�mUVa�덒�7���W����gh8�o��LRh�x>#�Gq��(F�2���Q�c��utК1��8�sF���ݠ�r':�����p��(�����aF���WrG�*gN�a�7��9��Ag>aG�� Q��ՙU�}����*�\T�alXr#wrk|��O�kɨȍ�˷�Ĳ׽�/�z]��6y��-o �~�/q�}�h�Q~nR��T��]��%t��}��7+Ս�glhi1���([R���j\�jR��Ci�ٺ��ι�5
�Z�������l���Y�﷫񗶖ǜm�ב�w��lnI��w/��n�b�t�ۙn[�𿢉U��Ѳ�(]
��Xb3`�5&�tܗ��V��ww;Z���B����/��Պt�]�^�<1;�q���E6a�{r��9I�yV���*w����-�pCJ:��"��R��B�}.î�2N������]�VOMb�S��A�� 3l�J'�����xl᧜�F���zw�Uw%��W�iȟXv~�p>��}�W]�>���\>V̔"5g�L��U>��:�e^Ş�տY3!Ma�ʾ�9�5��J�޷��@dņ���y)t�)T[jkM�-�(]=�����d��	��P�-;��yo�����+ќ]M�*�6��g�UL�o���o��]��\�\-�}&�^��wP+���e��=3|&nW�4�߀��~1U
��4{ 
P<h���t��%��5��5o5�zG&f�U���\���(�nQ�N�;e��!�hx�a}�����Aw�-�z�ҙ�����B֑r"��n�zt��3�!��t��NJ��Cr�Y�%�W����4���oz�@U.K�����ە&JC:@�5�B�ѭ*.N��ŨEp���]�,��Ԣz��,��{��<P�͸��.ۣ�׃F������������hǓ��7;X��(Y�m��r��,����ս��f�0�>lo�]���m�7{:N9n�����D;\5x�Ȏwa�r5���ƞ\!�RgT�7]b��g��y,���vgN�'h��i�F����:�&$`�/��f�o:�Y���8�p.L�%ҩEI�k;�R����
��ݫ�9r$p�fsT�W8�P`T�Z����ˬXF�3��b,��ܵD��d��4Ês��oc�/ fJ٤����û4b��p��j�i
4�ܖ51�NL �a]h\�m� c#*\�(^1N�GLtϏX��eE�h�͊�Q�W9i�x����H袍0�q��F�=,u�`Yr�-��������{�ǰml�Y�Q�p|�P_U!-��f]h�lL�� ̎\[$�Zy����7>�t�@�J[Q���(�Ã�U��1�&d��I:�k]����✈I�CԬ�}�Ǳ��?�Z��A��|�|����ra��c�cCb4U�y�!��P�&�dђɣA�D�ch�6����6���E�hǍt��Q�4UV!6���Rh����$����>�/d���KDh"�;�5�V
��v3EQ����|mU��_�����LQg�Y��e���K�[��[�{�u^��^;|'+��<�����>E���'�}^�E�3�Xɜ���ҕ�̎wx2��$���>�+$2Yd�-5z|ɟ�^��+���2�[πf����;~�;��0�Yo��J��d���>�)'n�K��
8��u�Mt^}����#}�3�9����m>��s�2_�z�t�������}i5�ٹVʙ���������q*��2|�&G���Zi�f%껢ssrK�Q�Dc/D�}ܕnc��Du֝'V,-�E����h�4���)�1Q��X8��`=�帧�����H��P�+WaCuE�Nw�:eY���r+{w�L�If��/:t���=:]l�K���
�'P��[�~�܄N��.���x�:b���"�k���;-��%j�Lln�ķV��^��P���L�q�7!�V���(��$�x�uq܌o��<��ތ꾺}�+3��WY��0�޽������-���.�=�;9x�4�؉���n��ʩp=l<@O���IZ���j�f��l�V-����償�ŵj����'�Tp��Ź})}���{��!�幙�뫰p�U�#�ۊL���*�'|��w��J@����:�[�gI \��+���y���M��軻��9,��W��l��EKL$��R$j�Nϛ��Ӭ�[�V�~}̔:PWu��cn���[}���E
����˺�����S\�{�_�	���͙����z�wz�T>gzy�nQ}�W���\���"f������ʆ��'W�8`�ӝ��|\�,�E�y�zF��y�۱��&��3x�k�����I��^���Q��S�,�]�~��f�������z�����$��x/���L�P/��M'�uj{W�^��ʫ�&ë{Z�3"��X�-AP�[��*�ǼK����a��a�<��f���H$���^bh�0��a�֕mk �z����.������Rb��p!�C8^u�%�ev����2�S�Y��l[���@�k4$��<Q%�T����>��_b���zn?+8�o!�����2g�s�U�,~���AJ�#wnתTڜX��ܾ��/z���QUY~!�8�I����Z{��N��C^��c���~�T�Jwڹy�j�n8DS�=jCj6�,'	�m=T�����Ѭa$�F��[�~�*X�e�ʑ��.�!-Ea��׊��A�rpd�b�^L�|cnM�W�K��Wgmk34�:fӧ��ؘ��j��q޽h�-S�j&4LN�8�Ct�gҟ5?��25ڢ"�&-/��$�:�O���S�����b-M�V��լ�mn{�W��c��Y3�ve]�wZ��1.:����z�YT��8<��ە�xp�v0�����F7Y{��Xo%�өJ����lN�P#�=Wv�ΝJDM���{����>���ڮ������R�d�>��Dg!�ߵ�^��'�q��dg�Nե�0�{����@y��hE��P�j"�<:-6�{!���\��V�+�s�)�'c�)V>x���.�V�܉kb�r��r��Gi<Pr֪~��@��X?���n=�����~,%^�S�����:q(_�y��U�/uQI6�����1�*�s�������Bl������k�+3!�F�?W3�RO���n�P2��I�x�OѼަ��~������VAZ��J/p����o#�Ɖ4Z߇�-��ĥېo{�+c�e<�)����h�Z�;vx������Oԝ�����>���M�����hL�G���=�(��faў��[���)jގ��Bm#���)���@:z:5;D�e4��6Z$;_�"8�l�^�_���4Ӝ���#��VdhkD�E1����D�[��H�r��7��B0rp"�e�z*�;�'Ôf�c�������=[�+x~�31V��=s*��~�Sp9�xR�h�8�^$��N���0ѷs�%��ߧ�8l(�]N󕚇�o�C��^�{ν�i��m���y�����J��p�ۅmC�˙|�{�x���}�]l��o�j��$���Ѱ����Wp��7M#[��t�M�=(�a��ǡ���T��L�]�o��e#�7��2��u
*j:ٷ{����B�S���w��׵}��;���Ȏ��F s�=�H��1��kd��=�j����p�����uc+��s���k=���/Kw�Y����6 �Է%�2uv[=�R5L�VO邴�{�����*s�)s|-3�q/��q|�9J��1�#>m��n�m�y0j`Z�T����P�x�6W]'���ݸ��l3����#SQs:�<lt�ma;h鮌�\V�1m��-e�;�mg�m�Ḇ��h�`��=S\�7f����qQ2WB3�N,D�1��u����2x�0P)������!bw"��a�B�Vdnش�Z�2�����?A�䆭p��5��a&�'�{6�w�6��C�*8`Hv�`���f:t�["�T�Ffv��n���N#��������iq��u���,�ٛ�rǅ�nP�[_��	_!���A{�̥��ݏ{J��~I�I�v�u$�>���*�4k�m޹����v�%o���T�o� ٵX��u���`�N,�s��p�.0�'��D�?\v��w��|��;��5;�;�)�+�Ga&�mu#Þj��	6\�hl*��T�s�!�_�����VU�3qb N��#�����tI�-�Z�h���(�A����k�{��������y��DL�����(��0Ƒ$��m����]��R��*/�42��(�ߠ����~��1]/���a��M��|�Յ�a� ��q����7�aS�G(�d�HU��C�98E�,'\�+WѹY`j(�;&���i"�29�6�8W��>#�Q�y��
ޯ׳��փ�0x�P���0���L3q�p��^���t��ɳ$#�6%ή�5��_�i��moق�SS�ws%X��f�@�4
x��*�Y�2��խ�4OF�ژG�Vf����&DC]I�9*ȂՐ�fJ�}��:�{b��zX�[���do�!�a0iY45���w�L�Y0Ӧ����-��桜�7F����N���W���XѴÇs��dg��Y0�Z�ɓ&��Q=��7MTk�v
x2x�cAq��`���|��Û.0�/�5皋�]ow#'��2N��k��z�m��ܣӌ�	�v~�Ɏ�}Wʸ#Duf@�M�	�q��뾳ǣ'M�R/��/��{</�?!)0F�,�B,:w�?aݞ/�Q����L��>�c�����j/� �7��]��.d�;V��f�n��=Xی0��DNo]i��$�gS8����x����w���c�>��MsX�*]8Ey[�v�$0ܑ���]���A�2Ta
ABI�2#B5�]��y����y�w��_J�}o��|[ח��ؔ����өY%�m���Ou7�Z�`���]JD$� ���s���.v��V��*�5�>�Ľ},V�1�=�$�x֥+�t���M�z�gA�5�{B��D��%KM�S�����٘�Cd6M���D �d7����/����yҷ$WƷ(wu݉&gcŝ!��9d�s��z���=;@���u\��z�tl�znf
]������?̚s���>^��o;v%����4�p-�z ����Aj�{�KY�F��h��H��ZÜ��s���Ovq����Z�;h�f-��p�آ��N�Uv�5�%���Kjm�E�(���gT��7�M��cs#t2����N-#���Nz�7TJ9*cFe�;.�g%���KJ�W0�^:<���D�Bd� 9q6J���L���9�&@�֡���4��Cs����(u�ڻF��p�	��ۼ��a�:�@�Y�7��y|�uIpGj���,�QmR��g�L\wA����E��ʭo�tUp�t�N�g����:�8m�$9u����:=��L��2Q��6���+`z��PW��`F�ޅ�i�_ܭ�Z\�mG���mӝy/�'�ݗ��XrKm��9pӺ��9j	G�ڰ�VU*f	Q�+u��և��ܽ
_FM���
N�Q�
��[ڼ�_o��ty��m����3 ;�{X2�q��"䒮*d��&�7��Q��*�2e��O]�9�!�d��9�<�wnfĴ�cR*�W}�Qy}�(��nmgB�5�]h��Wۀq\��gTdJ�Թ̣}(^)JdJ%����̃�QFA���������>����OKj**+	DQjKQ��*�Z�Ebŏ�c���-\��5&5U��[���0Z,XѮm��y�WH�6�O]m�kƊ��5G6�
��-�Ѩ�5�[��
,m��ъƯ_�����.!�8�,f�n�����P��Ӌ��������z�S��g8���\\d)�ca�l/]s��h�D0M���>4� @�n6oy���};��Z�'�-��n�}��G���rŭ�����I���?��oa�k�&���C	�9dss�(��q�<Y��9m9�0��K��G��'��tɂNk~q�υ�Kb��`�+�<4�v�umged)Ɯ6I��[K�O�Ӈ���?~?0���N��g����V�!��<{Ju�X��S怞7WZ�������rۀ��C��zE8�a�مc&g�Es{�~�OY=�('N6���}@@"=��-D���Z�	�7�k��C���s2�G1�F<�g��0�a�-��4�Hd�5�sկs���[�����՛.���^��n!��j]���}�B|"N�M��.T�WS[��ٯn톳�>�G,��c�c�R�Z�E��s
�T��6�6mّz������c�3������=p.�h�C����O�'���ғ�¸t��,VGb���5NHR��y�#� ��ǩfze�|�c;͒�s�i��[�:�L��m��/}}~DYx�C�w4�A�?* �|D��l��@�K)��Q�{n*����}tj���`��ay.2*q��������V�9�b�P~Z��e�}L]קߌ8�?��s���2]9��^�vv8���a��H��h�n��0��.3sv/#,��UU��5�5�Viԡ��1ࡵ��>2x��8�j��N�4-UF�E{9�[\�6�V6�6r�9i.yv-���"L�x�;~!��Ψ���"P�|A�;�,ི"8Kt���k�d[���{o�H�Oý���{��j����I�ٝ�>ޚ�ڵ5����`����rؑ4�8�N1����vg2��N�>U�������%&E�3r1��ax�h����wa����c�6G�u���KA;a�#[&�Ӵ�uՉ����X��s���&Å��E�n�r1�dI�.n$0,�5����� �^%c���E�n��f8I{l=Q�>T�ym��żD�u�S�d�o�q{l�X]�!�A��v#��u�v�iy���6Z[\O�ދ��_N`�;�مJ��֭��r�~L[ZB����yS_��Ç��o&�D��1�n��ь&u��"����L�$	�z"��F�o1Oygj+U$_qŗ���4�F�����1��� �Q�g�|t!�Dz[�H?FsF�M-p�[{��T�̞a{�rœ�#��[��(j"*f�v#έ��z�c�:�є��g�yDԭ���Q�ɇ�Z
xa�1!q#��f4���O?t����<�����ޔ�Q����L���Ž�ե�6enx��L�1(���Z���Ib#��0Ev:8d|�-�۩[/�"�ip ܷ�h,6��9�l$�˶D�O���w�U�渷���0S ?��pr��3a����uD�.f��(�q�kY~N8�l���3��Z�
��&�j���x#��8C�tԔiiaT�k#4լ$����<d�_�������z���h� ������	��iM}�z22\�D& �ar6�L�o�s�;<�"unoOn�L!�9�#I�a��0��籴�:�N��7n�J!u��n���Oc�%j���Нlǯr��c���:�v��C��D�gh�N8;yK���|�d��br�X��;��wm��c�b������m��r4����/\0���Թ׺W�U�,��gi
������9�PF0јH�N��z�Ku4k/r��&�P+�L0�h$�<����f���f��n4Gl�ȃ�ˮ{֐!�=ti��*bniĥ	쩥[�7�Hsf�_�޿�1@�H�x���BB���t^���_tLlvf@�©�ɲ8����_��цע/�������.�Fk�ǰ�0�E���L5Ƽ���v��oil��7��r�!.,�;�m��a��t��¹��k\l�Ɍy�Q]I�l����z���dXkp鯿/��1�����>��аE����ȣ�_�JS�h�J8j���?� U�0�G�E�R�e�TL�v�'�]�-�w2�S/�����������iȭ^��tw�1.��sH��z�0�T���"���b�$'���MLi���|���?~�8���,�.a�#V�c&g�5�~o$��nU*��#a�O?��b���)���"���bn��&���v����q[ΰ�9hg���1����Ng�V�{1���q�1T�������Æ�g �#��b;��A�:��.݈�Ǔ�{�"-�\�i�
����;�%�+r���7�ḭl��x�1��a������;���[�UW�N�4��O.x�S�?9Mi���&{��E�csq�a� �Xkixk=v�E�x���+rl{&~3�A.�_���
���`�Qĸ��0�~�c0o�^z��r�q������7aJh;��>d�e�K�V��6��s�g>�]bR��/ے�tv��53����`��)����)���|�F>z�x��i���w(�Jǣ���[QNnK��a�ES�\h�����r1��"��g �q���0fѨ�"����R�y�ߘV27�8Qχ`	u�Ӯ��n���x�h1 ���p�M�ȣ�^�!76��)t��Ҏ���T����>(Eg�*���K��?q[�ޯۧ<&�����	��4#
��k��tƖ<��􌐰�~Q�ߍU�;�wz�KQ���`g/��r�l�Ҟ\#6�O�t�u�&�ЋQ��h��
�rp�K���W����k��n����Q��� ������o���_��-z՞(�$�v�p.�H����,0u�:f�C���3�RxsV��ȣ��� �ۂ��EJ�(	�N��UhuM�=�Ɣ��on�'g|䠒�.��erӉ��S�B�}|�;�ai�j9O3���<��2�s̹¸�\tҷ�#��,������MEK
5\�lٻ\���ȳ15QD��\�Y/�߹���B��1��(a���"��7�mΧ9U!&�J"��(�i8zy�$qx|S���?ީ�sE�>�&*����FkL+����F�[���3vuEr��K����$d���IG&h��4V��>�xhڮl�Zc5�"�Y�u�c�6l�����O�v�i�-��y^�j<h�EC8]�X'�l��kͯ�.O^][�:	�K��#L�q�9��<ܞL���L�C��r��񢡉�X"��a<ّ̚����v��3�_d&O��y�Y�?
�E�Nm�<�K[QR���KZ�(P7Z�je�U�\�u|��z�!Sj��������n��[��Ѵm��֏2���ļZ��/��m�L��m:�N��;`YĴS7]���}ڻ�{���İ6�86���sE���&X9h?+5�[�c��Uu�p�8۶(��i��(o\�_q�m�ޤ�I�I�0�W��c1�a��@���8��."�F9�{��-z�c{�:.wki��񗳇+�\��-�E��&P\�bڋ�A�a"�Sۈp[�p�n�oj�}�K�i��2��36�F��y�b{\T{���^�C+���Y"g��Dg�d׌3����T�3̈́+�y�؍ƈ�5V�^d�X9�>�Y������-4(=�1k�*9TG]�ױ�����g&�sMœ
�`(��FQq,�!�H�S>�s�s^���nT�>/xH�tI�����l�CP�Q�Ukr[J��B}8Дw�Aƨ��|9QB�rz|��d����&o��pI��`��4���H%�KI#�H;�3Q�A��|�a+\���<sZ6_N#-��.�e����~�����6MđI��ЇP
�P׬Z���a2䊧vlǮ�]l"Zzx8T�k�K�����Ӥ�4iC��kX.k����C����N@��Pa^��8�u���pL3�V���޽��m�q|o)��4���ǵ|�}�y
����U�9�5��#�m؛��6Qhj%�x!�8�ᡗo��^�<��	�O'1�Ma0��0��m��4ד���l�\���||Q�Ƶ�{�g��ӷZ��e����<�Ek�na�X���<hj��W�/7��٫I�;�'w������:��<�]��NK�:Y���%8mQ��&U1o0������ҙȹ�rLJV\_Dsx�uv$S�;��6�;a�52.�v\�j*a��#�����MѰ��8��A�Hv�b[�s�%�QM8�}j�;y�z9�S��c��&�nf>y�+��ʷi�(eD���T'n��j荻Y
ܔ��yػ��F���5v�#�^Rݗ�"	���Ω}]&3��l�)�Uw]��82x��8e�wj�%p�xx���v��7�_i��ҹ՗}`�Ķt�0aj���co������z��.�na[��Y��>u�6E"���W��>z7��D��4�ح�{/�6���=9�t��*�
��4�A�ʾv�ECs2�w#�.	�!�Y��X
�{)��A%�3(24Q�J�?�Jʀ�F��qՃ��0�TU8�X��6��2Z1�Q�S�B^,;VP��u��%����y��b�@PmT_e��|C����&"���<eC D�/�:�$��g�1�Ke�SEF���O�`α��d����u�Ӷ�IR2{���Xf��'�;S��k�"�15���il3�,ԬI�Q� 2���3d�����v�ȩ�	bC�A�lX�%=�9�"o7���(�EM������T�*��ȍ<z�X��D��P�]f �H(�ДeP#F�^1a�?	��f^���S�Ǡ��;N�g�p�$D��uُ�}������o�\�|��hƮ[r��ڹ�-x�r��j�r������X��ս�Kx�x��cZ��m��5�����MW��{m�J(�\��x�����շ-��������<��� O��u3�>�MD���cv�nr�v���e�Lu]�S麏sZ]���Ы���b�	�w����^�� �nI���Z%dK�������m6n���^�`�j�s;�ʽ/�I�̀�@���F!��Sð�a�bvj�Ww%�<#F8�㒁�
ְ|�`���8��*��{%Qx�(��B2�\ᓰ�Q\�����dE&�l4Dt[�U:�w��1ʧg��iN1���j;	Ɨ�D�|)���}l��Ec�V�b⹈�Mɨk�tIZ½���:`���1*�;�d�/J6��-�G���\[�tFk61("֫l��n�V�;͹9�m0�-��d�gm�I�v�0�3����o�F?	��&U7;a�n��P�������K���iQBn�*�C�ׇ���Q	��<�D4Fsg�O�W�i/�)���|"�RU�E��v2�5��u�6�sY;sR0�r��1�p���p�0���<j��[�銀�ȹ�k6���d�TU_�sd3}},]5�L�eh�s$^�����+���kA�{C��q2"��7[��5�8SC��B5mj7��c88F�L�fW�i\�O�kM'�%����|�������13,fj!6s5�T�q'��jY�OO[��<�+g����\=[O0��I"|���jk�Mݦ�]���[q�$\0�����U�q �sqyOdV-e��sE*��ul���x޶���v���m�@�q��� n��*���=L/�{\_5h|����f���]�p�j����L�_�x�z1��o&,�+<gԷ������ӧۣ�?��F���~}����"�]>Gg	G2ګ��Qh��6��XnH����r��F��
	u�w6��j�K�')3��	1�=�A6�[٢@t�`weX�gONy7��_�K	8X���7�\�O55���>؇=4�T�=Eu�����ͥ�����t�2{�YWO�L�����qA�q?�u�3Y��L�4��9���Xd��d��v[���G5kiZ�[\�>0���>G?���:ܿe�HNZ9��w3�w9#9����S"����;i�cܗ���Ň����D���M����守'9�-����ٻJԜ�ӄ_4%����n��>�[ �-����-�l_;�vb�t���B
�Lsg����F150�J-�sO���_;������'�m�찉o8֢�ؘA���\�ܥ��,M�e��;ѯ%���r1ė	=4jɵ��q�X_u�~߂��O)�mE?|p ��!/6��J�u�h_d���s��R���ԭ�U�@5V�˦6���ht��!��]J�`#��,�Jo���8`���k��uܴ��~�����y��G#��f�ч��2CIalON:6t��\�FԺ3̈́uT˴t�Rv�sN�q(��C��6yM�:���"�ƃ����_��29{�ߌ-�%1Mņ��œ#v%��h�棨�;��s�V�Fr���`)�1Y���f|
#-Y�~tt�����x]��s��`�C�S[����p���odq|<,]>�Hێ����"[��yd]���2$�0ڇ�5�[�j<f�nCŋ7��:��4��{p�$���I�D�)�{ޅ�;VMs�����;20᠈6nl8aZ��"�+#�6e�k��d�p|R�a���n����Xz�*�&{��gۍ����a�C�B|�����O��fye�b�z���^"��8/��Qǝ�`��!>�NQҾ��Ė�i��dw�|�#���v@j;LS��aq���Rx�v�����Z{6��-��o9ќ�a[��	���e0���5;��Nt��pci~�GO���E�)|GI��&a�����`븥׺�vH!��};����e�'ɘK5��22d����㖨Wʮ�o0����&�m;��[#���Of(��׭��]t�՗7����d('&�y�+��0Pխ��]����г_H��0��ǒ\0ggL�=,��[nkM��9t��;mgb�`qX�l!�.d�m�YX�<�u�{a>n�� ��64�6�Dcz�X�Ð��vɍu*��l���..@�b�_��<�u�(��z�"�W���"�o�LP�ΑV��`¹!8����T�����\���E<\��o{q����#�մ�q0�;ʺf�e]���O|�壙�^�ZI+�jO���w�	O����{[�@g-mD:m0�����8��jf�Lz ��|)�&� z�e�-�;pA���ɳƘ\���p;���Q�LH�E��i���H���
߯-�,su����}��'������m=\��z.9��D�`!��&��A�b�Y�Di���i�uc�b��/�>�� d�u��yj���G��>�����p�y��B}���6.,\.vx���
��&%���4�h��Cux������8�VY~�������,�0�f� 郅g8Ã1��NLC^A�gCv�(����"S����(��_$�ǥ1f���a2����w�ן�Eg������/A\MfVÕ%�wG\	�$�SukG=cq�����٨U|��L.������E;ۨ/-T'(^ɤ�t��Ǣ0����Fe�	���Xi����&�cu��DeJ�w"]�oc�(�5�tى0���y���(�q��aӏ(`� ���O
(m��w>]�,�`r���R�e��k��Δ{�C��,Ѣ�KJi"`����z�8i�>�l"a�sfL�Y�j&�i#�v�$jjSW\�^M�=�<3�����6�P�"f��X=���&Ⱦ�gY���j��./���`���.h�47*��Flh����a�98G���bc�C�6̌"���v���;��d�2T�X�Ew;�$�����N
O���٩x7Mr�PS4�Zj;,3��H�5�}J�D�!���^{}.֏W%�dL_c�����WT-�-��ӻZ5�G�^Iţ�xq}�m�as��r�+MX���)�h�1N���]�q��m=,��ky8^8L�� �0��G§�*VUv�~ݜ"��I������~AD���0�����d�ȼ�&���I|,���I�a���A�gfL��l����w
�N�"��1���va�:~�f!�]��EmqZ8�F:�,u�����V�{�M���q�ۊ��	����2cؚ�k�6�h[74���oX���~�ⱋ�*�&jydj#_��!ȣ|���6�LpF$����y��:܄g(DW5L�冢�9/:aJ�/�rb�̹�V7����p�Y�\ہލ�L��8Q�2� 睪�m�̖���"�kv�Op#�D�>�i8�����9h��+�Voe`��uf�Jbp7�)�g �I:�j�����8����@n߉R�Xy����]x.�������Kj�v)���.���`����m5�m$�p�a�[H�9fr��y����4� bg<��"�<��% ��Ӊ��r`��[�4{���=���k�|Ś9��4�3Pqe�\c=mmM�8s��7��9��Gx{NS��r���'�u�k��:o3p�v�ӂߌj/�
����n9�N��nY�k,�V�c���	_��L�a��}LQ��T���ȹ�#�LM�p��7��I�m��䢏X�
/�����CcQ3�[��66+?X!�=�M�11MAf�;� ��swr���8c���쎆k`�I�n���$��a�m����[;bo��T�h�����ȇ�������x����T����,+�xݠJоݶ.��
�#��A�dB͍Q_��o�k���`ul9W��[���ov}�ohIRJ�w_|o4��Cb�yd�]�N�� �`VZ��^ۿ���r�� =?�����`Q�Jsj��Ű!�.h��a`#(m%�aoEM���;_:a��=�cw�@��dE�q�;��1v�3|���_?@FJ�Q	2f��Q��s�^�h���~�m �l6d�׍�_	9�P�?g^VQ���_�/k�<ʏO�1.A�7�7�<QvP�AN?���י�8�̾����� QG�kf
,8'ŗ��t��"F�~��sEŋ��Ax������ q�k�K�*��6��F4�ٍ�Q���%c���l^�v[ˋq�j<BƂ%��쾾݂;��?G�[cur��+����l���0��f8�mA��ͦ"��Q��DL�������`e�������cv�:��J���9N�MP�M�dS��u��{�iu��$[b�1��/.�\mOF"�6�}�)�(lN����Ra�{�%�d;��;YY���[�ʐw2.`�^��*��Gzn������Sz�
��8V#�`�ۮ�o��X��w�!�qm��)�\E��Գ;(<J���4l+������;j݇��]:I�m$�նP�tK�*�747w@I�7c&���nqØǃ� �W��ˎ�G�{h�]��f,&���*]������69;���N����ޥ�;+.�:��Uż�I�V���Cl��y���&�r�ۥ�F�`�	B[�(.8�ۮX�)Z�!vq���="�H�i�V_
}�;Yc7!͝9�v��t�`Pؽє̩+�k�`��E��p�%�A�?"�&�N��zO@��3�1ʌM/�ݠ�,@U6i���3�s��}T�C�,y��h���t���'�q^�y�\%#����t����(m�@����������]>ɺ�i�#N]lu�$��R�DA�3��݊�(��g6�K��ڔM,t7!ɤ�aF��:[R�ƙJn�eƓ8��	|��r���u1e�'r�rFiĝE�q&��g�������m�x��uk$��)s-��G�#s��ne�6E�B���&���ɴ�s�$�#��+��[v�Ә�\��C1J��PN�%T�Yl�C,���|���}{������k|/V�6����_�j��oJ�������5�5�oKomk�o���v��`֍�^�^�����okj�5���5�\�xū����z^��5{Z�����b����׍h�*�m^*�ץU��? !}�;��P������{����;��N����>�up��e1L��d�Y�����Do�kƸn8l�:Erq`�I�RA������6�u�r���x�0�n,r�e�J"-q������c��A�5���pГ��½��9"]�&&���
V�<f��v{]3|q'E�'�C�Ǣ�g��g��F�bi�d���������O[#�L���
XE��h�3z�@��\���z+9nMdK0���<d[9����hl7��l�ϯd�T�
:Z7��ZZǱ�8d\��Q,�5���a������+��dwT(ce4Q�sY�O�<VS�ha��F�5d�il�݌fHO���)���Q�.����L0�����L"������f#d�e^�4�y����n���x��c��@��=w}Q�ҳ�.���?�C���jD��[�)���[��R���_qcw7v�C���s�퓎FTv����wB
���2�wGF��M�(��0�0�d`��#�w�y��4��u�ĥ��L$��ӂ���9(�y��/A\r�Ѽ"v��:,u�㟚y�e;�$H�}:$��ݍ,�.����nd+4[[��j,6{"�n3<[͉��k.�ũk��my1�hʗt�P"?����&��	k�֔YΚ��*n~�.�
��,�7^Z������p,>6DSOJ������ke*��z�t������Q'�Kv'��h��꼻�D�s�}-�n8�k�{7-���s�#�~�	��:���w�	�p#�~6a2��[�ƱR��SU��}�������.L0�a�=���x�0כ�1l��7Z�CzA
6��-�T��fK���L���X8<���B�ID�[
%������+�+"b!H�^��spŖ�c,��Ԣ�������ҏs�x�FSI��I��Q$*̕����8�>ހե�H��hb�A�ܾ�a�/��5y��f�:�1�;��ⵚ����z矌��%�ᔸ��x��M��ᾞ��-��J��SY�ƩtQ�b��ɢ������W��]�<�kQ��gB&s�DM4F��X�&��IZ�0��l"���c�Dc�M�L��k�B2x�t���6>�g$��D�q:ȹ�J�})�n(Ȟ��'���#R�TVL+Z�~��-F'/��9�̃��8'u��܆.l����0��6�g7v:j`�CY�[
>���w5-��Sy�8QCt��,*�&|���/��6�-mf��	�m!n8�c���4<�}v
���1��(���i����x.ُ��mE�%��oS�ӕ{�IS8wǩ�]�3��/���!x��fQ���j�{X����7�/9��k�Ӡ��� l�y7���&���o!n�l���΄'�M0o�8�4�X�p��mV�p�1A��%s����4k�ݍ-!���ۭ$f[��D�߻;�ڝ��4��-��t��>�6���a�a��n�����\�c�m�<gZF��4�`>ci��|�O\�Սh{�`��<��Lv>���&7\-a�E��i��=�h&�Na1$ζE����q��>si�m:̋��%9����HA'�oa�׍DI���$�N&��Wg{_;.�	���OsY�g8h���XC��a����K���~�z�NՐ��f�f�����IF�)7��{�}]H�n����$-�2y,z������zVC/����frSN�]��[Y�Y������q�[�V�sG��YK��� n���}��w����0���c��q��G=e����[YVG�	6;dm���#pS�΀`� �O°�
Z%�9�O��,�ǎ&����㇏s&`�6�^��2�ǎ��|,��W2�G�X�\�6Xjx(-���)iuۗZM�����֮�� ��:���H/g˽��ԩsV�\���(��Lc��ő�Q�T����K��/j_��~�+�
�����(}�̚hqIY2,=�U����ڨ�d���n��";�E�(��Dsa�����rx]�s����ַ��C��pd�|j9�j0\f�É���qZ����S%�Z�Le�z�p���t��"���{3�9��;��g��ൽ��L��k��Gw/�$ң�n�#�wH�#��m�U����g>0e����.��HQb؇�42���3�����/����3����O[!]n��5����:u5�Er�����-]�Km����-��M7'G�Ȏ3I��$�b��v�
�����J�B׉�r�l<G���Y�4eI��b2��Z�'��z�A��v�3"�|�	�q��8�u���0���Wͭ�5w}�ǌK<���ٚ��� g[JZ��'&�ܩ�SSl��Ε��x��2����_OɆ3��=�H�^<��ef��k�s�W��\|Q�R�=l:�'쀠c?�k������*�?��r����4æ�`�.A<j��S�Uz�k��ñ��0<�8��Lkm!�(�0�M7fk�<��y:�8č��m𕮥�X�:Y���:;���Sn��^fŝ^�~��fN��B�q��`�����k��>s��RTA�ZU�z]y�F_Gݐ��[pI��㹤�c�u�����[��a�D9	��[^R�h�6q����U�3��]�k_�vvоP�r��y���a���|�S�'�jڈ�����N)��]N��Wv��m���k(�`�����ds-fι��W_]���	��nNc�N�0yl=L���D5N
̼J��f&�_G�q�w�{���v`�Եb	d��
F�'�DN	�~8�$��n_ω@S�gEG=� �*��a��/Q�}���c��߳���N-��.��v29���AE�[�lkWm���Sd2ZӴ��qO��J$���e�e��!���+U�V�"��=M�����8n��siF\��@Ӱ��;�UK�W��]ʈ{�V�NQ����)k���vgf���v�j�2��)]��[����y��C�6�a�a���Xq���s�A��q<����{/
���ج4!����Z�C�3�i�9ݕ\lp}cN\?����:�Ά:09��0SO��L�73�>�un1����&������sCuѢ1k���-�Z��Oe۠ڜA��I�me�^N�z��3��p��N4�wN#gBbe�T�=-��-sa�� ��1�U�+��AS3�(�[��d�Z��L1�yl* �0�Ǡץ]��f=�����������#H±��@�E��7ltf�Fه�������\��`���(JB�3���l-��5��t���}�8��a��ns��By`8C4>�R����C�;�ߍ�T��H3+A�٩W-�s_bO0vWs�Z�y�c����LqeAG��6�(b���3il/oy���{�-�]G�锲��I�o=_;��H�m҈<�.bc֚L��F%�ɍ́�c�|e1tٝ�Zh(��w��38�q�:G5��%�0$�ƍ�b��cY�x�#�����l#9�8#j�U�j4#�&F��a�����%���=]�?{}�@��y�R�?���]m9�Q��	�(a>:\��gԜ��3,M��NgK������s%�B5�o���7v�9�����nY���(��t�f��֟3

��F�!���V��7�����u�a�avȱI����͜�O����n�Ǭ���a�_r֡a�-DN3�����Q��46��<���QL3�b���k*v`���(ʀ~�<�(r=�F����+}�So�K\��%�gW�1���Vk��E���v^���d�r4fV�q��n�����[u��i8�S�vs��8E�4��Eֽ�P��
L�[>��Ӻ�W��?tQL���m"%��:����}�y���g
p�޼���άz!�8���\��co����U�Q��D��@4ö���(�N���{���̔L��Qϫ�V��Z�������~��	���GkS-���1�GM�L(�㺞���}6zH˪��3�L.|�帿{^�5��凱
Ax��Q�g�V1�ۨ��J#�U��n�T�s�,���/��8�A"S�Ѳ�F,�E���=p�6��"j�;p�q��!L�ˆ�j����l�<�C������?s'`(v�%�ތP0d��C�z|��*��B���}�����������vԱQg;�|�_A-V��]�ƀ� e隑S��O��V���^�_X��m^\w�B��M��c3!	�5(e-�hVZA�`І�M�t66�(��/�д���U��݇P�eq��u5n1p췹�9���c�5�����U���drM�o�n>=����]��z�<\�p�˴U���Ұ�����n��}1�gb�+{�:F��N�µos��C�9�Ny��s�D.�S|����Ͷ����ecb=�ǀ���魴�=�Re�k;��P�zg�Cٚ��Q�h��졶f]�9��
�������,W+?B
�q���<疝 4���n#�Yׯ:5d%��t��5�������jV�������h�o1�9T+չ꼞���U��+�����b㕨yK3���'\����MaQ�U��W�SCGJ{��ܣB+����7p����̵+�jm���Q�F�d��4NΊ�95g[����`�}]�.��:�x��YUw�HT��"�V�w���v�іNӻ�R�Y�Y���ܜĖz�6�P0���ods6q�����S5l9v����q������q5��j�/��l*1P�OR��(u&e�@>{���9�u�V���a�E���/��Z�e�p�[I��B���	KoU��6>��Ά��:�o^�װ,c����wS#�������7u��k��.N�f�J���ݎl�"�L�/�.��E��#6ޓ*��
��x�ӻsr(>�eo.�;�e�;���{���J��^��mz�n��v��n��U�W�<�ck�k�u��W�x��;r�ۛ��ڹ[z�v��W6���[[�c^�oJ�U�U{m%W�U{Z��zU�W�����\�b�^-j��kU�9���6��U;��7|^�zڔ3�5	������������=2��n"i�fG�k�;�i!sA�兦�`޵���������靈8��m������Fe���M�i,`����FV�¾#(M!��Sk�y�. ��Z}�3���e�=7Hi�L>+谙ۇ��]VRB������/rt��]'kh9G���\t�>[�Uޓ6�V��ٳ9��c�X�FƼ��ɑin�h�ɞ�h�10n�;il�Z��]푳bPz'�2�U�]��&4T�8��:^1���4}�9ir(^���^v�ug;����x���5�y�<\�����M�N�P�����È_�O�?t��f��s�kXA��,`��tSa�\5��K�7Q%7y�S��+N�1>dC[qj�	昝d��:j$n���!��gN��dB�lƼ�)�l�Nz��?�R/gRTc1�'K��H{�k1a��i*��U��dd�	�̵�}�4�`�q�a����ta����[K� �S:?O������Z��z�k�J�Os̄HNvR�����:���w�5k�9�Y��~�i�C:�R�{r�����}Y��ݞ�Qp��ـ�Q{���9��;v����%z+��=�Vtl��o���5xݮ��))�>T�3�<�g��juখi���j�B�wy��{�ʕ�l��78�9U�C�Q�����2�����/�XB�&Rl�<��6�u=	�G�e�/�"n�\���Z}�:{�{�ίe ��mo_��3��yy[�y}W��˻9�˥�9g_ I�L�l+{��! ��}�Î�7C��������a�\���n���|�k��
�:�U�'ۈK����l��=�x�)�����{��A<D���I\�v�E�\b�r�T$۶�\5�&Ū�mnc�9�Go?b�<>�s�B�w��W���2��}�ʎ䘍3{�r��/?f�@���|�{�c|�))]@��>_���gu�QHg�.������7�g��}�R�z�rT����/r֧x��1���9�r+G�Q�(.�Z�P��������AU�r,�fʔe�<��WD�����5үNa:�F溸����etͼ��T��ދ(G�&�^洢��<7n�_z���ڞ����X��&�t:�>Kı��Z�N������'��E���+OqG75^����+x�<;�f�"W�b{����C��ϼ���>��x5:��Sg?Eg+Қ�Rf�{y9y�O�⚋W�ޤ��"�2���O���E�*�Ir�g��mG����a�K��X`/M�E]ѩ�շ炳A�%�T��L�*[�fծIYJ
~:�RG:�;��"S~�Fm��8�k�H<�7��9^T����C�'d�r�r�6�u0={S�/�"Atu����a3{��AI�7\/�Bi�o��lvn����w�lNٛ�׆%&�Mno� #���a��Ξs�l����D�-d������;���Ś)�Y�q���uY}�Q�xa�_�n*�GvT�.vJ�rVV�zX%�JҞwy�[8l$0�e/�ٻ8������F�}�7w�s�+J�#'����^����i�^�6�����Ϟ=���q��s��\9KL��*I8��u�.R��Fy>Z��dWfOb���OT�u��47ٓ�c<q�}����bF�(�p:c}���[h���O�0>g��xc� [�N�}��𦯽~��S��'q�h��%4�^�|�ݛ����:<3�vy�9��9��N{3nC�XQ�\dJ�.��=I��<��(�2��Z�'��V:��6��=��g�:���&.}��a{~)y{=at!��<6wl����ϲ�����^/)^��d=8��}�Gs��m��]�o��o��+,Oa�f1�h���}^K_�3�)-²à=�|Ŧ��|��� ������ݭQ�졊�>c}ZW�f�u6��{3���I{�-�7�ѥ�iW��
�pmn�F�ew��E�����.�֑4CJ
��r����;H#'1R���3o��B� ��r�<}f�r�e��5�PR7b��`�v��>�uwa���V\��{6�ẅ́�f�{7�Z��)3����x�4y�ʮ�;mW�7�+� \_
��8փ��时Y$��myl�F*)L��2�fw=Ш�Lnu����x�[��~N��b�޲��q
-;�c-�^�ukK~�	����w=�j�R�R8n~�<3�q��>^���>�W=�#7K���wb��螾ٞ:�~�~�o����^��f
����Ew7p����?p�~�F���mw���2��:����ܘ�Z���{bN���`�26�Y�n:���3���6�'*�VqCu�Ԇ6���|�p�2냇��X�;��Z�8���g���{3��W����I��W�<G<��	��s7!ؼ�34�Ue�'�U�,`�w����^�(W�T%vOv�'K�p�{E�wM��９�=�_B�h_c�r��{�_�T���0^yWG��{r�c事�d��O-�r���+��o��f(�ᨳ]�C�+��3ިǇ��Q����V�Y0�}����'���E��)���Z�����~�]����ܨ��&�����
��έ�>aVy���K�r_,�,�U�\�T��֓�hR���W�����R[�u��M��3g2�p�yДwv+=۝&�������Q��Vo�i��/�v�g��<�VS�xS��:��iP�v(70:�G����g�<zGZ�J��5�Jy�|����%���ݱB�}=��{x�حjZ��z��yP��חh��d>�(<M��~�E�ܧ<�3ي�C�ǅg����9{�}o�(��r�hr%���i���	�]�UN����3u\E�'^�pwլ�%j^�}�Ǘ�\)eJm��jzvZ��������~t
���7iд��������r�T1�M���F�Vd�w2��w����hj�%<)��o���{�+����V�e�������ǿ7��h�S9c�C �2�}�Z6e� ja��X-�N6����
��I�1���em.���12j��)�����!m����C_>)��\�Ǐz{�<���60����I����y��t�J�{�d��q7&l��>��T<����OQlo��9=���ۮ�3���[el�~�]�<�O�Ni]깑�z+��v�ϡ�,�}��Y弻�#��q?>G�>��f������'�u�HE���z���}�z��������o�]�V��bE�=s��V�]wx�ګm��~��P|;�I�� �!I�1|Bs	T�+�����D�&��y��yн�W�ʫ����Io��t�^��r�J��J�=7O��ڭ�Lmj�Z����mj�W���Z5���m���+m�����WZ�����uuL�HIc �	��[j���?G����[�������V���_���^���5�/�BA$B� HC!$ 	���D!�B����C�Bd&H̃ @�	�HB%2�L��hP�4� A���0�$�	B!	fL!��R�$��D)��@3&F$	�"`�"@@!�	dH��#���������>����J��W���;�>/��7��������|}��_;|��v���~�~���&`&D�D��L��!He"��4c6E,i,�Me!��F�,�f�,�H�2�Y)IE4�&d0"#)L��4�&2M)�d��JQ�J�JfI�A	�JS2�R��fc$����)�DLf%44Ĕ��K4�#@�$}|�~��?U��[o�gO��4eN�)��8(
�� ��"��H�������ػdC�S��K�UD��=4p����T89E��x
�
����ؘo8��5o�xP+�&@�y�"�H�[@�@p_Bu�"K��R�;#]{���c	|j(t�s�AfL�����X��Um�w��_~w��y?���^�-��T�m?{��^Rֶ���j��e[j���-_����N�j�7���Ȁ�ٸM��V!��y�*�+�,���[[7����hqD@t�ߴ�Z�=��P�K`G��f�6�HM&B�͢�q)❇�I>'��w�����)��2@�D�c ���<��ܗ�!Ǭr�L�FG��g)��$���NR���[w1�*9�P �^>�zQ�-���<��Y�U W!�@�E�|7����j7�ّܲ^�R���B&�P}��}ЇH� vL
`���4�0/*�5���l���-������i�����/�V��6�̘�[�x�&�p|[�^�����ߋ7ǜ�v�.|���~6V�[�o����Y�%����6��������~@pE�s�t;�"lSp� �Q�9)��[�$w0>��Ff�?@�;�r�bNN��I$~��&FgR��x�1�N��A�MbO۰�%>０� ��κ��1#�e&J=;��^������uF��Z�m�mU��UZ5�����Q[Tb�TmX��ڶƱm�5�E[�h��Ŷ���mlk[�[�Qmm���j�ڢ�lTZض��m���i+I[kڣcY6��ѵlU��ح[մkU���FQ������`��>�A�7�==��K����Bv�h[[�"A4���0�bN:��� W�N�m�0m���dG���_4�0�Q�@b4����9XEV�6�[d"�!D�(M�.�K�;n	d��,St�2.�il���D�{F���]p,(
�@��3�	�ky��"���Fn�@@W��֐�
:['B�Z�`����n�d׮s�a5�'RA��D鎔Lsn���)�����