BZh91AY&SY�8�՚ߔ`p���#ߠ����   b9^�  ���#Rj���JVf���؍���R6���٪���ll�RI�P٢JIR��UhkkKm�3�I�*RB��5T�M,��l%34��ڬ��A�U��R���Z��P�Hֶm�ik������L�+(��5eQm��Z�f��Z�� ��.�{�6�ĤUi���*l�Ƃ%m�2�ء���*��[ZKd6iUl�m�6ek,d�j�I���P٬�
����VYD�m-if¼�y偪V�lx  [��:�h,�Պ(嫰ӻ���u�ښ���;5ѓE_v���lUzq5��[���RW!�J�V�[	;�T�"l�T�ZYme�6��  ��}�h$�r8�M-�ꗽU�yKYT�=�;�=S*l8z�=h�ͻc{��l�T�[��-+K��x�.���v�{��7��B�wp��9��՞���5%SS5�����m�w�  ;�=*}{�Y�g�T�/x{��ޚ��St�笍۩u�{Y���m�U=���|��J$����%v�5����}�4�K֛�޽_f�	Q���H�j���M���֙j�6ĥQDkk� f=�/X=ٟGϾ�H���Wu��� �޺4˻���J�-�t�|�y꒫m��r�)饱���j{ލ
��-�놕T����gz����*ǫu-0^��w^��l¶����c%�l�
�� }��_j�@�^�B����۩Kw;��6���R�=��U��M���^9Tu��^����ԛoy��Խo��5D�n�U
�{o�l��kI�aim| ��7�钪W=��+׻J��z�K����J�ˬ������m�n7m�{p=J۹L��9��T��q�q�)i���:�4�UK�Q�:�kRS��kR����ej��Wfm�| w��}�+g�Ty�w%@��移�E%K�ㅺ�`hm����UP��7zoS�IJr��T�B�qwSZ7��]�^� �x{�@
�z�k&�&��l��[i| x=@����Moj���u���8���XQU�`ƴ
�z�:<���ח�u���=q���tw�n^޻�u�-�Ɩ��E�IK���  �>@���`
���=�
�{�=U�]�epz�@���+׶���ǃ��n�z�vn�z���z�{��thz{�EYL��l6[kl�_  ;]௠��N((9n�u@�6�
�&�=z!�3����{c���w�]x�z秇�$�g!^�c�        ��R��4�aL `���{!�RR�#L&�2b0`E?&!)TT`      ��BJ���� 	�    S�UTM2      	JRBzM�0��d6�LĞ��'�����f�,~0��"��d]d����%�دf��twg�#lC��n����  ��=�\�W�|<���T�DQQ_/�����XwC@�����~O��������� _  ����UU]q����T����2�����?x@"�A"#����	� ��%D0B�{��A�A*�B�� �*�A �@�"=��A	�$z	Q"=�/A �@��"=(/A #�J ��%Dz	�AG�(+�@"�
="�A t*����U�%A�@ �%Dz	��J���A	���!Q�T�%�� :	^�� =�/���@��=��@���A*/p���:	S��:	W��<)�@�(t/G��zS��:	��z��A(��t��B�t��~��'���z({oM�y�T�wr!��f�Q E��.��n��W�ޭ��M����LT�3���v�U�P���^Ѭ+�$랮%J�S.�^�hk�9)FӔ��ڀ�j���	<�t����{x�Z2��
����y0n�[�q:7���y1 mVm���/��vU�{��9�2�,Ô��aG��m��iZ���#�Y���nn(]�uwR�)��Y����e��� :��MbCvj�z�Q�X�lKŖ2b�m���yL�V���A`�3nkt�Or���1�$�r�M�F2kl��"�2ir"D/5�!V��lEa�+6�n����ض�n�x�D�b�'S�	��.�T�Ѱ1O!�T�#�������Df<W���VqQ��2�
f�^:���޴Yf�(v�S+	T�*�@V�Y�%XJ|U��)�-��mj�d�}O9ӡ��lIu>��đZ�E��wT�#t�O���P��j�72��*![�yy���u��i�w��\���ׁYF"�*(���Dl���D9��L��p��8�@n��{�7�(�.L�A�r���@���L#�n�eFִ
8��ј�-����:��F���R:�����O+�$%j��N�x�!Q�#��]�Z(ޛ�.��V��.�^#�I�`U�^m�ѓ5����V�9�F흐�l��֓C>�b�H�9���q�Y�:L�ha��[X/3�I�Z���a�3B[0e�U�5�	�1�j�C�V�uPD�Ii��b�k0aq�ɚ�|���m�ɸ酴3#cq�j���H�܊��A�JXI����A֍MB�p�T�d��/a]f��q���t�ip�����i�u�	]�qV����Kp�q������ <�Y�(�+�V��6�
�!��WNZ���� �aC��M�n��N^�ӂ+'�U̘�n���V�ю��N�O������l�C讜����ޚ׈�5����)F��/��v�)I�H�
Ӹ��i3[��T�_*:)�61�{J�J�s.�<5 �5�����Pҷ*�L�`�b��J�r�̚�J�-hf��b��76���{�-`�uqӲ�be�ȶ���Z�WMJr���'CPWB�t���sdzR�����Z�2�;-H�7J�x[�
��ݒ¸Tb�ȁ�ن�kp
Iim�1���G����P��T7MX̥�6e�(��a��vA��y��M��liӉ^ҹ(O�`�����L����kk��9�k�N�4���j��_&Z|m�؁uu� �Y�eus��o-9��B�U��ZZ.��L�#{���ь��VF
�[�ǎ'y�3��L��r�)`�E�L�{YH���hR&b�N�:�/rHě���,7X�(X���jf��<
��+8��vt� w$wFE�f�ean*�]�,�p_��h4�Q"E��Q��Ym�����`�,� �2����h Lq������Y>gN�0�":̭�~˭J�*�Ez��)�e�)���$���S3w��wE�C�I���ۖ9��.�2b�	f0dT�����pn7㭅F¢sk�9x�w�������b�1Mi�5ZDr�̌բ��i��.����w#�V�7z�ZV��@��h��iԵ��;��oFv��/�ց$ܧ�O�{��wuuhfmZU�q�,��m�z�h;�TWd[R`�6�6���n=eRiL��=���*�&���Y%b��n��v�-d$����,%S�4�*�F�n��*�e��Gvԙ��,UémD�I�����w1 );.d�n��-�.C������V$۴�����Ko5��[yKm92�r�/MG�)X�ԥ�C���f��6*<�#`�Y�g��A�ۓ+j�����cY	Tq��hLH�7���p-�9�+�KC�Φn$��6���ޠ�����0[c�Z�� �I�m���)��Y��ճt�h�b���B�*U���gHs�Ӯqz7q�I��h�eRA5���q�Nn�U�W�p5Ϩ%m<���Y�z3���X���r�qusB��2�;���z��k�o���g6�ڴ�Yyb�U���{E_es-�^��L��Ô
�l�֭��5�Xke֡�T4�8��jm�S��t��]�U�nQ����k훻�n���o@�w�n<�
� �Оӷ����	�Ԭ3��()Fj��ݒ�nLS���̻cP��3��,],E<̤MК�7FSZ��T��[��-5�I�*��f7X�A2��%ѻ�C��e���c��ifkt3s-��f9F�"���	@��Zޫqb�jۂ(b��r�T/j��MuM���p�@!Q��Z�Yk(|ʬB�a�GJ[x>�k+I�N��`a�t��2f��`�+J*�̡3�yI �&�m=�H��] �'�ve�$��o�ִ��N�四y�h�����D��	�>�nR����
4����v�F�CS�|�VZV�6�y�g1���#��Ra1�"�[;c
zV�x^�]�`ud�!VHse=ԧ��Y�D�!�]c��wr�Cr����ꁊb��S��akdHμA���3�X�G~$�"ܽP�)D��Emm˫"�E�r�0-m��[�SKC1��8��Q�3,mm�Gv�n���E���b��i(V]����uTc!��֦җ�q�*�7��X�b�`��Ve�f� �A[u�bw�p��Ȇ�ҩ���]Bv�b��4.D�#0��R���Yuw@�3�����)��2Nc0e�ĵ��~O ����f��un���g[��o�v�lnt�w���e��ә���v(1{�Sf� f��\U����i�IAj�^���
fX�'��lm�sf6�"�J�1iC�ɡj:s4wi��`į9&~�[tV����t-K.��T3R�oFf��p"���I���*�9wXX�������8(�-�%�Ԗ�30���	CqGQT�b0�(|�m=��Q��J��W��=iY`�ub����R�lY'n�D���Fd�T�i,li���l�(�7��v]�v&۹�,�V�[,���s1�Z^O xKSv�7����51{�;\��$�C%��+e@�ɼ��J%�XkY�]�ɝ�O�)˾!aY��yS�)�M�d8H�J��+M��x�Պ��m��X��:)m^P�Գ�Ћ���owWλ
<ðUo4{�c�u�^`80HѮ��-�[w�ʣ]�P+T�� U-3)k�ac�(�t`82���>�(=�Z¦訞��4�F�j���(�4�z�M!�6�;��[����e4C4Z�����ܖo+�\�����!CWEWq!ڢR��C��Y����G{�b��0&��A)=�����&l|���Ä=*�ڎ:��=hn�jRGskon�%o3 ��}�M�Q�L�a��;�)��f Q[z��[�5�l�`s~N�ն�b5���;��Llٴ��e��D�iY�@j[L��)�U+J`�Ska�^�������Vv=��u��n5�t�t�.D��OD����h�����Kjвa��OMm6s^ǅX��#C)-I��[2�JU�f^�C��P00��W+5�ˠ�x����W�5@S3W�5ATF������^��Z��̨35�ZZ]��CjԔ� 4Aw����V�*~-�;z7T��5��;�I �W���x)ws�ӽ�Pd���唋S�&��`۬��5�h:t�N YG6R֚ �_����1��3DU2��0<�6��zYx�_����pXhnf��n��c��AnXbke�jԵI�Y�1� �HY��j�n���N
�J!Ǌ~�Mig��a��f��v���K	K4۬���P8�i�tT�tÄ�/-�w#in쫭I|h�a&�c��h��6�đ��i{�Kt��Mb\9x^���D�/2f��̀��b���N]$��M�
���	�4��bVv$ո��*uR��'�/\*��Hp�gReւ)��n@�ǹu�$�Q��Ҳ�ٹup��V6��t��`�t1B�Z�iZ0	�k0m<i�b�/Ō�y�G^ً�Q[h*@u���t6�R�S�n��t��/e�*a�V�op�qTX��[%����$GI�J�`�B�1KqҥXiT+:(�+4�/,ջiBkf0�mt6�<�i�T���;ZYD ]���J�*��kUF�[�f�.�����f sM�pc̦ƶ֩x�� �-��h0VF��G0c��M�8�ח@�Ӻް�9iB�wYv�9��A�Hf�ՂEI��8�;4����/wE)������������ot|��85�j*�~�j���Q�)�&��.,�V7�Fqm��Ce(���m�Q���0t���Vf�*p�*YDw5YR�9���,b{,��5Hm �MMJ4)-�ʘb�\�eР13YN#/7啉��.�G��Y����]��LV�|$��H�m沓��̆�i�ͺl��^[�񽫂�V���ʕ�ϭ�nA6�W�q��I�������N;yt��iCBP�ˑa��Z����Gv%l��)�GhZ��&+E�+0 18�2�K�Ux�4�ۣ4�_���S+J��m��M�:.�f�P�Y��n�2VI"���ыp+�-��B�A�)�f@N�ݫl9����V|�5z.���7Z�,��q��35����/h�t�+uG��������XޘСP&��yYj�*�Kd#���$"B�2���^<!�GS
���ۊ��i:�!;�n�ޚ:CĤu��;��X͙�U8�j6�rn�W�k�M��L��t��	d�,�Ɯ��wl�V�Zz^m�����B���$���=����:"�H�4Ĺ�Ѱz�N���h�+�pKk�YLu@���u���Ѷ����ܳuufR�j�W�t-~ځ
�n�x�Ɓp^���z�$A�n+�B8�X{{{�WM=ek�6]w�LO,� ���ehe5F�Li�ZN�X4^Dk@��1��Q�������C�9��6�J�e�fS"c�Ʒ�`�6��l��u��b�ѭ�F��Xӎ6��ƭ(\���K**j���$�x�Tz���Vo�����:�C�J��dM�ᢎSz���6�[Y�at�@�G i�İ֩t��q͚����Efmإ(%��j��B[��Ô��4��WU4�-&�a%��h^.�e͸����C���q=J�4�8�j�"�yx0�4^^�X�QŮb��iYNIr�=-��G`E�!�i��d�/�qArpr�[xv����'Z��[m,�����ݴ�H֘6	cY��V��8��Un��{{t�d�;v��sH���M�O�Lә/M����1�FKǍ*&�M�쩻-U��ֹ�Ĥ�<"y�
�L�]��\N�Hۤvó���*�������kݣ#�+�M���f�f3Ra`fw
݌bX�YD]�(��LƳzk(�tŇ�@���
��j�Ձ^5FTx�m�'(hn�V�JS[�A^13
�ݚ��o#xm�o��
X��Rb�Q�κi����GS�qR�#����d)���.)I�*j��@4�8��/w!A��
ϊ�YGA�U��z��*�e*��D��fc�3�y.i�sR0٬�kDz����k)bnk�yeh82ڔ���B� ��[�3eMh�#	�$ٺV�{RԺ{��Z
,�q=܄���N0�GYsKV��k;i���U�nQ �Q+U���`���$�����3�OV���h
�cH;�aouU��eX��C��]�D�
�qm˖�L��	�*��M�v6���q�[A[��t��0h�:�rOu�c� SG{kyj�K��d;O��%��d'Yu�-z�Z�bw�� ���d��6�v7��-o>���zM�l=���	��V��(;	[��^�U���w�عi��HX��αNŚ6��lx�s0e�!��]:ǈ~L�Ԝ��w��x�����0X6gJ DF�7�5��ڒ'za�t���"�9�Sc�5�i���n�Ki�n�f�YvCz��b+0�lw+M�b�`��If+��m���-�V�9n�vi5v�mČv����QAQ�7h� ۥ`2�;�/t1EV�wa�_k���T8�9�V�s����f�N#��1<F�p2��,�X�YU �Tֆ�
�f���>/"������=�A�U-�\���y�U��4�)I�w�Z�E���h̅�p�]�o
��E7wJ�u74]J�C�A�:�u����1Wz�OK�oFl-��u���3�Q�F�7F�Vc��3T�V����r��KE(ݵJmZ�`hbP5�b�V�j:�/m�@��*�r*Ƣq�w��Jre�$��wX��p�E@Rۭ	� �	¦��7$ئ�ո3<��J
�V]�vcTm ��!R��`��K�%��wX� ���V�z���Q�Ia��QT��o�u�� ����)�R����"�ۘ��1��.�1i�f<�K��Ƶ�x�)��TXMc��/0kv��U���;���Xa%kf���vK�r���q��ҡ Ѧ��r�� J����5�$�p��x!)T	m��a��l�O)&��7%�t�x���,��nn���x�Q�)�6MQml�x�Ĥ��7�����sVcOr��B�ZJ�W0�Fa2$� ��;C )�8"�u�\�s���k��+3-t=�� ���䠚���	�E`.}�[|�Ya�h�_�1g�Ҿ���a?� ��"�����`7�.���a�b�j2�S����V�7��7ta��}_ᓄ$�T�@�Ư&��4���������~���ߦSSE(�vx������N�捠�P�(��hSN,�UK����������~��xo�����_��4�J]�f�|�����]Rw�;�z+r&Z;�&�nz���(M0����j8���O�sʺ�],��}�Ïk;U
*�M��G�cH���=�}՜ǐ:[�M9��ә/h���Ӿy��GI'SoNgF㜙y��Lwef�1�;o�v��R�9|!x��Y��*X�5tL��m��u����9���B�k��~��ƻ8���p������C8>=�����e��vf�G���>��h�O�+d����4V��*�*v���Y�+r�u����)9.Y^dݝ�`��U�-TǡV�p����n�HӲ[]J���F�яQ&Uu�@��������"򺕼�-}��%��5s->J��U��v
C8:�/���UNE%�V+@撴0����Mް�*2�V�&�f�혫Q�A�f� R'q���k\4��_D�.��*���VI@K����R��d����x�?�������v� ����.�lx��}�v�Ħt��0dQb�V�鶃������������X�vj՝� 5�R������|���\�!Q�Q˙ߖby/���DC�D:'����w�8��Ǣ�0!:��/xm(F�F]��5ˢ,���u�5vp�Kc�E�TZ�zj���f���E39���I4��j���w��J�^}��
(�b������ђ��͈V�5�6�����Wv宵l􈥣vč�����;D��j����Nt5���y�Y�4T��K}��9�1��p�!���Λi��MvT������b�YQ�N�=����W�ڽ�\
��.�i�K`Qh�{�r�仗mWp�1��'N�o�`�n��ruN����X�k)򥺱C}�,9}0�z�[�r�f>����7�Sge�Mil�ش�a(�b��q�:i��(��
���B�]k����^R�Xy�(kw����*AXm� �{|�ۥyІ�׶b���R��&��E�V���dJy.}r�#!����g̧��}���R�a�)�ծpm]��)���|���+��41�j� A�@�*fi�c�ǂ�����q��H��+\�j-��~̻J![][V���3�=G� �h��f��}�{Qb�F0<�Bx�;�2�W�VX�KT0�%��5i��,�d�����[�G��ʵk��5Խ�s�	����`-L^��ڹ����7�Woet`Rܝ9eJ��THp;�ozodA\U������C��i�ݚ�]*��l��].�ޛ0h��K8�W[k#��[<7�e>���rn�nP�at4��u\;��z�35�2��̑Z:X�B��s��Tzfa�V4�T�Gp,̡t\b|7���YB�]���4�T�yG/\,D�������`mq^�JH�a�z.t�]Es�P��v�&�ywH 9 ���e��̳�q��n�	�ֵ"(��E\u�><�xl����sƒဃŦwV��ٽ��gPC��;k8D�3��	�m�X����qLuά��!}}���Yζ����R�K�5�w!�;y���t��Լ�8r��`S"E�k�L�Σ�~ٝ���J���2�{���r�SK��ِ](������|���h���uhPC-�d#9�����d�`'A[5>A��1*7Z�=t�VK�pif������17v�
ڰ��1�x� ���t�f�+n����<��>ت�${h�kz�f:��	Z:�v�͹R�[�7�t�����M�DfwaY!�)NWʅ���S�:oC����u�VzY>�b�7��WT�Ou�Υ3S���&h���x��4�=Գ�I�sK- �ŢX�չ���bbr��h��m��p=ZN:�[hmE  ��"&��Em_J�s]����5{`^e�j`r}5�a�et�6���6��ճk�H	YS��QE|�l:Ӷ)���$w۹��{�;X�hC^q���k��di%���`�ǹʜ�nq2��nܭ�#�[��k�C/mӈ�t7��Ϯ���"]K�Ǥ�E�1ᥘ����M^�5����t�_4�S���_�F!��M]��i�p�,O@�#&���z �ܨc��S�s�qzgC�Z��K�:�>�T�%��12pUck ����{3�$���Ǿ���C"��t%�m���L�D�'�4{+V%�B�wfξ����ٵtv+�I2 m4�7����.u�d�G6�� G�
�β��xCe�`.�9�ms�6��J���}��_K
�H�c�%i���D��~�5'�m��=���ܫ79�0��YǗ�h
+K���$'D��|�%��[�hp4���MAd�q+�*vݰ�}�ʂ*K���
�<$�^�mԚ��6C-�*e�}寻���7.�v;��ϋ{d�M\��$G�%���YBѶF�����ӫV�V�D�\a�W�t�Ǌ�N��JP��K ���)�� �PއN���kL��=ͩԂ�-�E]�	��q��:�9EV��"���(��TGi�b��X&���]_+9�QW����n�황l��ȴAX^���xM���p[e%*�@@�ե�K�kf)�.���~Kos��!��qXʲ�J}���;�,��PBc�����P��3�:Y1t]��.�6��iT�m�^R:��j�6�27, ���;��Z�l=��ٱ�i6GE�A�k��k�A۵�	��y��L�������wj4/�%�c�/�D�l(
��1��`�+'W�o���J�t6nͩRMvk�a�=���NM>iT�m�f\ՠ:����ki^�f(v��Qˑ��&��WQM
L۩X�d�)��s��n� x�O�?u<�p�g�Y�y1�ZkR�jX��vVL�B�;΂K���T#da���2�Tf��N��z\h��5���(Js��ه�7)��@��N��p.��`��l�'^�S)���'`��l��˶�='�O}���\ʬ��"<�@1t$����"�@����>�D���֦I��oL�b�*��q M�L�1��ҕK�3P�hPC�]����|Q�轄bK���ˎ���i���f��CXͬX��wX,���n�k��m�M[uYha��ZYb���sg6��{�@W;4��Vn��j']ա�8���}��ԳZ4���R��R�J;Y���9l����Ūc��sSx��-�{{I�:��J�Y��ɚ�ۑf&ݜ�Oiϑ���á]9��N���ņ�_l:ڥ6ntCk���Z) ��v��.�	�DȄtv�ga�w^��-�8�]���
6�k�X�)��2�v�2۱�t�������������jn���5��T�a]I��+�p�7�y9-���]�\W��Օ��ۂI���<���]���.1x-Ь=ONSAj��l�9�!G�єh275�Љ�8�N������I&3&��L��6�k�.���l+��&���@���@[RQ�M�ЎaB}���.j����"TI��8���3E*쌈�ގ:��7zn�ev�����J-��AҔ�^v[��yڢxOCt.���Yۦ�M]R�wq|2�J��P��S������x7�d챭�-��=����m,���c�+�3�\���h���9��Ϻ!NX^��ۣ�誊��Y}h��V캊��W0�i�}R���F�.\wz�T.�D�;7��5Rψ/3:�h�oj�'Eue%ۼ+)����(�XL�3^#��ĥ�FiyF{�(��w�;���Z���]4�+��Vp&[�c�ya��
�ʂQowYCi.K��
���Z ��sA��w�3���m���B�H�)�]�g�Wv�Z0D`���6��\�\�Y;�yz)R|n����T"`��i5 ��;�{d'�'v7��^朊@�km
5���#ƤKGWǗ�r�w��Ė�ekT�����ݳ$ɗHɈ!F�����g3Z�����r�m��J����f�˦��;m�ע��$��)�u�ЅZgB�I�p��EM!V~x�ص[��V���' ��R}��:��[��qS����v3n]:��'�t&��A�8�:�iV#�/�����
Κ<k��Kk�Iܺ���/�l�JXޝ�� 1m 8j���73��,�`{-��Qc:�sj��)��T��V"�j�«dǹ��S�g�`��k���(�����	����`�g�=�����)b�X��)Waf���^nN�>fZoK�b���9+Fq���ug!cU�������.e
����=�0�����;�44���1մ0�'�Ѧ[�Q�J��ٌW�w"��Q�W��1�jA�鉗�oݮ��맒l�|M���:���M�Ԑx��vF��Փ;�iC�G@i`�:R�<�:��z0��ѩ��ق-eo=�N�,�P��t̄��]*��v�`��4�u��?mуNk���$.$�o����8���}!&�LËh��%�7O%ݠ^r��L�lܾ�y7�����:/��Dw!�P�-h������W\��iX� ��ff"�W��j����4lS�.�;D����נh$�*5t0�b��r�V^���3,H��Vv�r���@��I;�F0\��mC�j��=�p�T7R"=�Ɲ�Fuf��m�YnB��!Z�am��ZOG��
+���;OkDv�坽SV:
GM�\��8�u�aT�-E>����Qe�ς��5p-g����%��W��K�����e�bb�S�M����_D���NU����i=��G3�Q������U�(�;��+��%�hj��o��!�:gL�y"���G,�D�ڦ�N�t9al�X�,�K�nK�&��Р�D���rr/��t�2��	�5<����f���P"�t�4+�L�Vr"A�qoJ�����{�@�����
1It�%�,��=iX���=)�7+�K;�4��S[�C��2�-s�c
;;,�Pi[���ٜ9I�Vmmm�ŀμ��p��_6ˊ�t��Ѽk��׀u��	Ҧ��W����Rk8��p�vņ󭋈A܉�����������S��PΤ�զeƉ���.�3�^�|��X"a=���[�:�K�AYݾ�%�[�h.y��� +!]�zb���;��i�u� zn��6�I�l7WR��{B�T+*9G��.ƶ�Ǆ�n��=���Zﳆ�E>���O�Am��h�0>Ѷ��d�WO2.�t܏[(qBma�Q���X�M�Zmd�ܤ�S3�d�s�lR�����O�Q6ȥ���]�1<�v�*�h�Ĉ���ժ�w.����]�T��iUd��!3ky������8]�Z�e��Zh�R8�����C���z�-��>�`�˘օuZ�.hMm҈��8@P��	�/F�����`V����܎��).}YB!x4hX��.�4<z�6��%V�����@杇�JH���u;eL��&3��O qN��,�J�]X�q�u#��7F���}-���3�}�i q'<|,t�1��Ɛ�ݸ���˛M��Na���=[�(�P�f\Z������)�����Ve��\�����C�m������xJ	�.K�#�ste%��ɐh/���%�[m�H.��].*.��G����
�aVdA���+w�[(�khY�iS��X��M���ʒb�slې,؊�k����X2ʕ�p���黻Ug��m���Ĺ7��46��v�]� �є�K�����k�n��ՙ{�;3����8���ʕƶ�D[o�g@�&\��ܱ�]����j q���w��H���[�֝�]���������v�cXʆc7�&i�i�Z3�+l��{[|�m^�ꕍ�C*[�Tb�nV�v6{'d�w�r�2�K�qjԏa��b��M��,��e	-i��4��QjQ�r��QWN���\Z�KvG�Ut9\nhx��L�]�l��A
�q(�9L�I��̩��2�{I �p���`�r����;]��V*`�鍌����f'9��#�t^��zV��ך_��{kiFBs7��+������3��**$� �;��b��U���>��y�2T{&���M
��\�v����P��(�}�E�˽��
��ۛI�E@��71���
}:��79�H��oT�ܥe:�6�p�Q�EomJ�=	v�GS��wW}�sʗ�է�JgrUmv'�am��9G�y���*8�v:�tr#{t�b�9.򘃇vG0ɰ�zz۽$C��]v���'�)EZJk۸�U��ҧ[���;n�ȩ#������p�=�c�K��D�Ve��U�S�s�І���t:)�xâ�5� �Ɓ��A��LV��ctb���v�n�|��\�;n��Z׺�Ŧ��Z��Cfԩ�v��E�h	3��⋣�}�Sɘsgp�����7��t�:ͫډ�X*��k<(��2G�����О���έ��F�g]#�q}/����2�Z׷.��8R6��&��!	�� Z�Iʭl��s���n���Z���ť]�)�Lij%uq������rlS�I,�(ǯuNVs��&�/�l\�H��w���/RZ����s�2�(����PV��6a�.\2�S�^�*48u�����
�K���[�lQ�+��(��GO��-���Z���,8�(��ږ�ܻ�����۸/���o��6I�&�e�STE.�dI;�VsF�)�,���7Z��>��K��8�T�] �A��5$Z���� �$RJ�|�v�"��������ޑ8�2��I$�I$�I$�I%�B�u:���EL��%,��C��>� ���SÇ��
����<��.���;8v;1;�<�z��US*h� P ���>�^�mҧ����V@���}_}_UW����P ��}o��ǕO�?
�/���=���h���7�U����[�y�����`�s9w8��8i�v�z�Z�}fT(�Er�evj�fT�C�T�J����!i��'��#A��iЙ�q�I����ZT�,�dcU�h]�[5/7��p���rٗW�ɥ�U�����HKP��E���Ț�d�vadK�gf��y'ӓ���:ct�Van(R�i�
Хk"SN�mv�+��Û�4��}��͛{��%3�Z x�~z&��7@#{��1Zx桊97���46�)�}B�n_-n ���7&'�reu��F#to02�t�3:d�Z���TBṵ��d��-��X�d�7^x����'*$�\B�4����g�pdv�5��B�Jĝ����}tcU��\�B���>���S�*��v�r�������un��gÓ�Z*t5�@{��m;e
%se�=;r�㗛ʻ���ba��J�$��N��ڴ�s w��`��E唫j�����l�``��(l�����IKSL
q�ϒ���nv�Ҿ97�i��FZof�%,��4a��.�5ԣ�ʖ�G]Z�a���\�<v�`8�v�c_R��jGBA�V�Z�Юyل�1���e���&I�V� :D8s���:%������{MqS>�f凉J�)xR���j�L�aW�L��KY����:���� mv]3+�)8K��}�'��pKF�9��2P���m���hݐ���a�(�)Q�
��>8��z�k	��v�Ȣ]Õd����^㒔TxM�r������j��Х`Ȉ��rT���MO��H�or�Sc7�۽��ɘ1�� r.�X"1��0bν%q�Ӱ���Z�
���˶@�诅�	�!�R��f�)ܜ�(ػ��[���bY��`�t�ME%����]d�w�"��2���Y�rgQ]��س�R��u�����R�t�.�.t��3��c���ޤm����/A��Mn���}$�V�	��q*9֛�-ã ��[Y{�S_�_R���+:b��KT\ͻ�%˽�[q�t]�v��S��h�[�@a\���d}]��H��Z�O��e+f�e⣅4��Qvv_w0�������gr*�~6��Bĺ�O�8��yts�ɘb�SWj�_C�Rd�L�9Y[tzٵP�wl諫��n��\[�Ӻ�5��M����ξ+�����Z���5tᲖ�a�t�*�v�[�s+K�Y)^˸˹��e�Ѻ��������(I7v�GP�������w(i=y��75y$�*��C�r���{�v�!q�s䜕C�,T[j�s_�cp�g.$�(�0Ui]cH7�h��vXs-r��n�������w�"�uR�kW(u9{ĦP�`Ii�u���T��0w@ﲃ����5��#�d���[�GW�+&���0k�+�2k��TR�٫�Os{n�0�vbׂ�d��W'���|��4�Go3~�y�m]Z��j��T1u]f�R����G�C0ߎ�A��3����Ą�}�@o��Mp	[���.ܮژ�i�`�p���zv��Z��v4��m�'M耍x�u�+ٸ��y���%ˮ��(��>�����8Q�-��_Q�&i׸Ga"RI���o���h-z�[���Q�f���T�ٖ�c�w�&�v��o���6Ȝy���[�1���F��K�΍��5��k*S���!EkN�k)�w���+b竩��m��\v�9>|;cjR�a�?��s���� Y[��0f�@�!Oh@,+;�biJ�Nu9��;�A��d�f��F暭=�@�&�R�(q�Y����#AP&a
� ��q�++,΁��6G�9�j��\稞!��2�P/�O���k�W\�9�)<�K�01�0r�8v�����t1�\
���w\5]�'��"�]�_q�$\� �D'}��w�e(3�9Y�pȧV�.%��*����^ڗ��9X��@�G+.�C�� �0"���թ����7�+C�$���	�b*֪�B.L�;J^ح����E�:i��M�-A�+A�^�S*�/4_BX���n��%xol&�Î>��H�'ٶmEa%9<9����P�Ȏ鶨��fn�Еtv��
�M���2󉧻,VT��°;��4���� ���T�z�uF\�E�w���V�ԹCm�-R�b�i����U����0p�`Z�q�����{M���<���o1�&RD34(���1����.|�[C6Q�h"����w�����s0�h,����EQ��K01.[w6V�qRM�Xӡ�u���[�-S��\�46��\F���K�ұAD\�u+�qd�#(m�G#���;��C��i�7��JK�i���EH�gE�ۗgR܍�A���mE�n����J���	R��c>5�@ 3��2]�c�;B�F*a^��zs�l�oEI�4t-���65L�K�Gr3�F�jv���EhB�ܥ��`3�'5�xQ�����{���ج�/�GZ2�,�P1���i��u���5Z@��wu\
���7�M��Y97@Uv�����zqz�iU���5��j�$�aH��1�ܾQ+մ��-�2��GωpA��V���9y��(T�i��@7���sN�Գ �p���׀��p�6.h�y�gc�e�Xpi��<{�vժ�)��>\��n���S�/�:��z!��Fnlx^�Nsz���Csn�y���Gvt���dx.Ya)�/�}�y��=�c���ѽ�/�{ț�Є�4
�\}4��B	�[��G�E��O)�o�������(�@z��9���������d���$�P�{|;h.�3�]nd98���/�Ѓ�C�ܥª^�;@up�>.��|�#8C15S�j���˺wݣN�_8vfq���vg�Y4��X���b��̼�[��ih��l �>�}DY�usu�!=�/Y6�]a���q��8���z���뱾��n�؜�@��E�]]�&]=Ӂ�@b��0,R����S���)m-�w��4Tyr�f>e;KEe�t��SlZ��
r�=�xS(b��)�*toa��ݸ�_X���γ��@����,�J��V��ye�I�������i/$�/��̬�UJ�3�J��M��)$o�f��I5+)ei���r�YbE���ǂ��pm�Z�lHҖz�qqQ���n�peK7"���q�=x��.~��z�\���"�غN�lk  � Hʧ!tM7���p�T����ʗw���y�D�1��O:��Vi{V��@e��^T�@�A- �R�K�O=Ι�c���x2�ᔦ%+[��	���Ep��vhpg؀��ݓᏢDL5�X]�{�?��:7F���hޑ
Ii�w[;��}X�Y�]5b6��[�^O�f�����8���E�F��>/��`����׹����h��++l�A�I[\>�E ��u"�4�̓.�˼	�����)<C��k% �*ov�ɤ�¯����6�أ]�5�wk"QQv+�чz��]0S��]j�N��@�SE��.s'Q[ٔ~z��=���Wx�Z�!�+Rů��Dm�u�g�O�{$@gn�{�$^@�����r�-��tJ&���я�m2�A�o&vt���Ok(�c.P�{�d����{N���vd*�u��Ts"�])���}Z�s���̈́�g��ͳ�e��}���v�!Ilv�k�S*�f�T�ٌܭ����>Y[
��mE�a�E��}&�+��ql����1V��am� 4f��EѢ��ؾ\zwa������q�;.��fۙ1���o���Q5�f%"c�й6�`
(�p]��-�bQ��n�g�X'[�,�/b��@���Q�,D���zg{�gb�x{u���LR�}|�fnR��x��5m�Ӗ�JM,���;I�:�E��9�i�= C0U�-��B�)qN���2����ߙ��:Ql��e[̏'^���#ek���5"�t���k�����t�
�JbKaB���;]�[-җ�b���o6������U��6���/�سiD����O>̻Q��yB�8�*S�Y�S���I�Fk��6�kk��iQu�$�؋|.m�0먽\凬t N�X�\:���u�/p�v5|r���Uԧd����nx�oN���巖I�����2L�>�\3r��ഁ�e] fff�S\����YI�1V����0��m��6#��S��$v>5���Ĥ˄^Tكi�h<�s2��7j�*�iYX�0I��0&k�V>坠j�GWl���iHb�8�E	��N��\QL�t��/N���c�ZM쾰�E�N͉��}�!�G��eL氵��6X�i>�w�N7������j���oqWr
�LV�=N�	��☰�΁��B���\g(ea�k��Da�h�z),��a7ڀ]8�����G�[aڦ��
��l�_R��ͤ�������۶d��#R!��uP{��h��g����[����:'1���*���������#�+�J�i+�P��Z��S��s�Z+�������]H�ld�uEjm��s&�:d�ڼ�O/xbA�w2EVWV���㮆�j�Lw%ZW�%���=i�1�����lVw\���eA�I�GUFY�/x��v�1K�
�9�7/x�eVҤ�c�T/]&^��@��#.�V�M;8���GR�:є�n<�UKy�U];h t�-�w/��Ky��V�t��� �Ȭ���"�U���;}��b�=���@��kN�q�S���Ǵ���`u�Z���A�oi=��N��}f�����e�%���eu陭�\���[q��=Nn0�6���K�v�ٶ�2�
��)3���uʘ�q��WC��D�A�U�d��o&P��yr\��=�ҾQMgU�Uj�v�*ʛi�L2���r�+/l[qjE�אm[��߷�9״Wk�r�5�iV��e�[Ӯ[�Z*9`j��r�pM{c�emV;53)i��/�%��^��\\RDP�����[ �*2�fs�A%s0������#ל���4��/IkvY5tl�[�P�A��B�����Xn�=����Uh7e�l�[bܒ��W��w!��wx��)���Z�*������8	J����bp�Ưi���.�����5��omjVsΎ�	�n��%.�v*;�Xu�ej �Ϝ�b\Ij���BJ(�k��yY�Ř{�Eʾ��P��w��[�V����U,Zc��SR�1�)�Z��u�[O��n�ܼ��Q��R�[B�mtsM9��ry�4�+��.���@'��@��,���H�:	Q��㢃�N��Z�t>tQ�޴W�]\Q�-�3�]��8jq�cM����
���F��Ð��:��̙rj�����pK�@�	�p�{a�V��#_%V�I��p�3P��k:j-uݹ6�f�E��OrHUɬ�M+Lm�|,#�hS�:̈�(�|���]�#�ˉ�A����;��N�m�����HR�к�>�S+�-��*���E���w	�J����kY�y�F�)�5�������N;�g�'Od��r=(��R�K�՜,���5���*3X�j�-uK�E�V;��A�g絊��fa��ƚz��%2�o;-��t�e6k�ge�+�|�d��Ǡ��5f���X�+�v�/i�`g,T�r�6�wݚ��e7��;k���ڔɔZJo��#'�W��Vk0���2�``�U�Y/{�Ms"�`�UӴ�� �Ԯ���c�i���-�7��`�$�6�sfަFl�u������f�<4����������g��J�u�Y��)����:�+�Юb�sz��h�V�|���&�u������Sa�d[J-"�p�cr�$���|V��GjS�����`�\�tUk��vq�tWU.<�K�rQږ�n�*e����;j4�̰[��ml�zW;MpvS*-�ɡ��w�� e(�j�u�&+;�Z��o^ӼLjk��@�~TjV]������}m^O���u�n���]E	\�Su���h�R� �9������Q��XЕg9{p�k؍��a�Lú� U*�"5�|���=�-J���6�v�v����<9�]\��֦"��mD�M˛����f�H٣;)��wv['X|�a� �T��G'V���U.;��E��N����͋9S�3����-ǔ�񐪎�5yp�u&��M���m��]�u�XEcC�e�l%ʛ�m���ک]y*<q���T�^��i�k�׋s�y�\�lz%���>=h>O�K}�mof[*٢��;2�]
n��d��vU��[5�xrKO2��f��`L�N��e#$�&,����)q'~����8ku� {�YyV�b�i`�d��x���q�E���`�I#WxEb�Rت]�v5[\i���G�7+)�K�Y�	ǷEn �`��y{3�V6����*H-��M�>-V�>�ʴ"�����O�Nx���n�'�8�ܺ��tb,���ڕj�]�rw.fЌR�r�:��կ�pZk�&\�7�&�1z�ګ�Ç���E�'	�(�DE~�H�ɕX0`Tu�ގ:H� ����Y�op�7|9$�zt�t��T8e�Y��F#��o.�r}�۫<�:�VF�ժ���eF�ǚ�ӿ�H���r3��=[���ce7���9B�n�:n餥!� �דk��X@P]V­՘D��˕ �[�v�����axXBNu$�}����+�X��/��O{[\wX�Mk��~Dd<�7O}1SA;\p	��[�1�wU��GC+�*�\ݧ��g��b��� g\�v�sč���J�S�P�(u#X�b8��D�'sPb��1I{S6�1Wm��mft�ҧ���{���׎s��o������TQ_���~�����?B4>���h}����h}a�?Wֿ�>�@�a�:G�Ƣ�\VM�U+ً�{ۣہɲ3���I9c��k��Қ��Zpp�4QY�4VՌ���.���� ����v�\u*;gu�r�d���AΜ��<7e��-p��B��K�M����Q��(�1l�)wk�:�!m�K�������1�w\Z�/]� �p� o*��9�:�	^��`�}r'Zmu�g&�7O���Kk,��.����N������e�7��JT{����I;j���2l�QV��u�������*�7)�=V�*	e㬕��1Q1k�97k*p�2�G �����Ɉ������}Ì͏_�\���������L\�&"N������s~���-�$f�XyW�ϧhg����\)]G��d�90b��_[���i��IM�t#��l�o*���v� ����5�;��+�mY����݅��Y��X�̫�}y�	��=�U�oF�z��8��F/��»���Y�\[jk�E�=җb�u�	�qU�zeB���&�a
#8WO3v�a�T���� �P����j|��+{��W�X���F�_6V��5-��#NP��z�c�m�v5�U�K�2��٣.�:0ulj�q��Q�h��%g3������i�;i�drI�K�WR�:�SWR��>NW}盿`�*���R��5G�SR�KD@-3�w��"Zh����*��IZ
��X ()��i�!�����h�d�4�E}���jJ��b�$�N@E��V�*�������b�i�*(��j�U4xڂ��k�%QO6)� ��������Б�MB�EUEAW�TDDE%1WkQZ�DC���2UQ0LMW-!T��Í5AEAETTUM$ESSQGh�W}��@f(63h��0�D�v�PTsb�����*"i���"�(!���3�b(���bihuT.��R�R�՚���2Vwm����$��w��x�_�=�N^��J:/:�%�a6�#�2;��yǫ���]J�'�U�"�7�>����g9f��إ���������֟?1��}�uD��ጺ�QFszr��s����6�"͸5S/���7S�.���5~���ܞ�i��r�>���u.F{f��L���ޛ��o��`�t$_��׼#�S��.��CR5�=���RWO���{��6���+�F�{�"�l1S��\��ty�}粞��(?z_;S
ŨߎJR�C��B���ׯ7�=�;�M����v�bR}޽�۶��!I�M�}��~|�;3��U�{��������emX���;����ǂ���&�uo�=�T�9�Ыd�9�����v|���b��u�뇞��=����8N����Ľ�4I�����μ���s�o�~��˻�K��x,E2�rS��OY�ra+�-	=�������e�7,"����G����z$(r������Q�|��ϵ���ߖ����<jx��#+)�[+/������4��z�G	��s���A����39	Ri@R9�ڜcKr��;���]���[ɒ�>f�K)Ջ:�B�&�B���2f�}%���O껆�����og�ta7�@�C;�Ͻٽܗ�O�H�3����ನ�pМ�P��Z�M��N�����z�\����k��i���=�O���yUqTo�"h�Ǹ��w8��N=$+N4vn�w��ۛ�8�qbsǚ�h�]h�H�74>ڞsַ˻�'5��;ݽ���mKzz�;�y�O�=����ɻ���g?^��[�C|���=�sޜ�J��J�^��VEF���]tř�wï>'G���v��Td��4b�jx��oNl��w�X��}X�-�Sν�K���~Kv���ŷ�[����Z���<���7%��ؽs��坓|���O/k���#u^�a_Lj��A���
��˕/o���6c
WHb���t'%_��������}�#��X:�ny��W]v���#��v��7��3�5�s7VbWZ	�����[��|:�p��(F��<5Zsss�1�pO���@��
���U��{O�%��,7�Tb��.�h��mt��e��v��LPdi:�0�e.i[
���u���:���Z�ۢt�S��6=Tn�T���y�i=\���<N�g6`�鍻���rپ���a�]��/N���s(�f�{����9������]�����F���H"�o��/V;�|��R�7O���j���[�2���>�y��L�)�/˴�-���X� �C����0�鹌�����v����R��u�'WQ�*�T7�3��Or��W�+f�2�����;9�YH�D)�(���hy�l;c]�q�� �dH3�t}�w���tsA���J���o^����*̋��/N�n����w����	����TA�Cjc�	�\�N�G�����}`'��������kN4�oX�^��>����S|�sdS:]���m<�o�	�ƿugS?w~I̡t��W����G᳼�=ݾQ=y��_W���j-)���f��z{v��GM����&%�}�Xv��8G`���Rя$WfP'ag.�+b�l��5�7���A�/n0�t�/L��k�è���U���(*)hC���9�*w̸X�'W��Λ5��n8��cr�ĺ1OM��y4�J?��^���ܨݗ�s����+��n�*�\U��_��uZ��Y�䪋���M�}���3�6�ܓ����;�����a%�$�''kNLٷx,vC]�n�ݔ�����X.�(w����/���ϱ�C���Y�����.dY�����^������=���{�ݠ�v���������{/ĝ�3f��Sv��!�V5���}���W�L5�%���_�E�zm\>���}�����O�Q��t˞k�;=Ah�KO���O<�)�G˦٧�{Vnm�̱��{��j���������Y�1t�mX�y�9�^��q����B&����o����O��׽��u�װ!��J��=���\^�Oh��sSx��y��>��7c��9�Ƴ(����S�U3�k�8��Ҫ��o3_���L�#�ɀ����o[�5��39���!<�n����E*��W�#�0D4a��w�۵쾁$�p3�: �����8�3�4f�,́ ŻX/=Z3+���l��"J&:��]�V�T�(L�׎PX)vp�-[j#oo�8� !��N���i?��#E^Z�<n�D��3h���V�c�kj�+���l�1oktE�7sq���8�Ňm�["��(�:�>N6dA����z� ��{W�׎޵�2��K�K.@J�F��k_R�Y�:�y�j~r��rL��;~�:��o&U���L�_@=��t�e�K4$0I�8�⮧\�y�G��������X�h@G���6��C_C�j�z��I�[����=��Q̩ӽ沧�X��qU{a��/�ޏ}P�Y������R�_<����f��=�zz�3|k�k���nb�d�M���ӗ����v������LO��5��rݿc��{]O?l���|���%o.Jc#q�����[�+*q���[��-� ���-����Iw�ۖv���Oԇs�s�Z���z��WϤ]�-8�̳�E~�Ω���^��Q�k�3ݷјf��g�{=���7�D湪��g�dh;8�x�oѧ��|���ʭ�;.�:�I�;눻U�$�>�Թd�����pG��C����R�x��S&לk��8��A\芘\�w�!W��y�)+Z�f�bm�4y��;8s��� T��p�9�/���X�YZB]-�+��"�d3m05ܾz���,>l�4���I��x���㻓�������"�^צq�o�q�6�>�㴖W~��B�����.��|w|��ep�q�:��<�x��\��T���^5m<ڽ7���G��/���:$T!�f;n�ݙ���U�L�B����q̪%�+�PO��pq�w��D{G���p�}��m/y����U>r�[�mzg�i����ϻ&n�2[�:}ޞaJ2N������vQ��9���ʿCAt�^��}���D57r���zsp�#ݷ�����N���{*�����{ND,s������xO+��赲,Z��������=��;����+����@-�ͣp,�����z�f�3ʭNo���T�n�3�$^���v�����f惌o�m��ә%���d�#��C�Fw���n{׏�ZW{Ւ��.���R��H���!�/|�0�2�J�洌.�����3�&v��A���z�s��ꜯ���O�um`� 8��i�6��{(C؍�6�S�w�<ܻq]r���Ɩ�ٵ{��1͖tͻL#.�t��3���\�r��<e^s�Uen��g�U�������~�J�'F/F�{>�)��YYˎ޼D�9�j�T�u?}�ϩq�w=�g�6��������'�!�x��u�^+/Tu���K��Oa��frA7tM����ogKP|�J�1<�i��ݡ<���z�I�k���@}W��s������I�b:�Y��rQ�͹�Y�_�vh:K7�5;��~��==�ᓗW�o���n�=@�䁞o�,�J��S�L>�k�׫X�Ϛq`ڞ�ʿ)�Uz�pg1����ӯ�s|'�)д�\p[}D�ͬ/C�s�7B_�ۺ�\����7��n�oEM�;���Q�ʮWv����8�U��o��nP�g���Ϗ��o�@��&���y^+�^��;��'ys��m^��&��B5����'����{ =n���9=�הTĹ��\��^/7%�>�^:X�^4��;��tW��,8|�vC��U�}�Hyp��а_�C��ph��E�%H�dЬ3�D?��)��:���U�]o�Q���*�vAS��b�l�pŔ���l� ���k����"�%j�\�*tOGX�QY1�o������[�,��iI�zZ(dp�\r,W�z���w3��>�5z*�({��~���f��7��om�	���r���v>f|jOeut?4�})��ස�g�I��H��ٵ��o�wz�F/��WW~�
W���?��V�r+�� ��2L�e�,��8fm����Dk�NѽNdh��t���72+l4�)%�m��ay[����:�k�Ջ}qg��`���`׼���y�ꇵ��x��S�۽Q�NW���Q���^8��dk�BD/EG~��|�1Q�v����55�L�t�F��`�w�,�ڳo{ُ<΋�v��0D�vh�7Ç/U��K�Ϥ��J��hfM��.����<��{ C����+y05���1�U[��1���|7I�O3=��=ԛ'ۉ��dv>^��Q�{~/��T�GL{v�V�ʯx����]���pJa��+E�}�ݚ*�\߭�%*Y+=��a���7E4�)ڶLO�F 6��;�;8�����`r�>S+`��"��S�S8�`�m��iO;}
��w@m'�G�,�z�X�*�ݼ��:TcF�V3�)���qP��eڂ=&1�ڃ^��ޞ-��>;���� ���V}����|��ͬf-3"��������yŕ�|��zG���]T�P��~M��,Z�����5�蟑���� �nk��ɉ��o���<�m���p���I���#U�T/cH�ž����'��EϽ.��^�yL�z{���w���x��1�`R���R_��^�X�5�UW��C��ތ.�����ԗ-~ȝxNAx��2���T�V����*���i���X�ڇo�Hh]b���:5���_+�I�j����C�_GT��w7�"o��Mq��'s���o��w#$�X&Ei�3��d<d5�I���MEA%��6��g�8�oݭ�w�^�A=Z�A�>~��,�NE�P<��g�Z��z�>=����Q�����S�o�����>�}E���6v��S���+Tby����u��������k��U��P�|�n��l��_8:m�8��*x����.�4]?W+5�;��T���n=�8-�A��V�bڰ�N�j�to0e���ށ�t��r�,5:7��j���	L껔�B��jݡ�I��EY������4���_
�}8�Z��ţ�]7v�`�;h�/��gXg�s���<u�h!ܖ�{䕃N�BK����u6���O0�:�ܳ�y|�{�Өʈck\y$�<g������@�G�Y��1��S�m;�����	5[�_�e������ɾͯGo��lm�Z��/�֔�����Ln�v�ޔ<�2�$������X�\�w�l��������D�+u��_�k����?g�q��5��ߙ���ؖ�/��{ӧt�����ϯ�}��^[��A��z��}g���j.:�ݱ"rSw���/��t�}�įa(�I�~�/\mgv�� �hV��}z�rm7����8~U�t�8��]�\R�I�p&�Z�����-���^�χL�����|fp��}����@�0�@�0�7�nn�������7��+~9r��+�Rd�����np������Z7�%]H�5,�m����vav~��V��*����X��R\����M˃����9ْ�G�ܻ��5tp�
�MOV���s�f�;p��4���tiq��7�4G`����A�h�+��t	�F��,[��a1X�ط-����0\3��H���͵���wb��>����{v�q�A@�a�m.v��%�/�9Js��R%W.k�B����e>;EѸ$�lV	{i���S�n;��Z��A���zT�j.k���4�)%9��Vru���b�ʎW<�ǯC����6��[]Y�@i�g���NU�x��e�;���ۣ���HQ�έ�9��&�%�B�,i��n�8\z\"g-[��k���+^4��;Y�/@'v�ծ�u9QB�չέ�re[y 4-����M���*]魴P������~{l_W8)v� ��#�]ʙ�Y)`m�ێA�r��t=��Q�EY*�G��lO��]�[o��ݽE:��D&m!��:�>d��o3�E��ˑv�m�M5��i�`�<6K��˷n��͟:�԰��nV�9���6�#�jtyo^t�)�D��ʽ��ϯf:���ٓ�s�|W,����-أr�^b_+�������z���Q�MV�'sDA�V�0���BMW-{�ǲwA��(D�X��u[N�'�VX�ʏQ�:�T�	��pc� ��M��w]^
�:Tv��>��\�6Q�G�z���f�p�Ū�w\�؃��xi�K8*��X�n�MCENhp��b5������y[m���a���F�F�Tn�n�{0
���Wn������4�)Z�u��0j� }�GKw�>�{���[�|�њP<~�ފ8�1�XZ��?Ǽ9��%ދ/���߻^2���; ��^�Wm֓s!!|5���A�,ar���bF��]�!n��� [�p�j���azV� �\�fF�om�J��U|I�AXh�O�(b`L-����{��K��"���K�X	�8�uӷ&��ո�eQ�]�d}�'Hi&U�j��j���L9����;K���Z�l�hɁ�ʃ1n��������Q��3m6bjF:+܉����nP]�mX��i����5�ʴy���W���˙�aTNm��t`�=uQ����-Y9�e�IPUz&��7l'�M��uD���9�ݾ�E�]���8����q0��+���c\�rWa�k\z�Q|���LY����;Gr�g�:r
�#��͸��(s��@E��,A�`�\1p� ��H<ޚ�J98�Rf�w��u����t�{��\�%�J� L%��Q5wMe<��	��A�/�ru�ɩ�9'[ �h�w���\\��Ȯ�-���w���	��=�.��ov��ӹ%R� ܾ9�T�Z�6�Iո)���δ�9��-b V�����כ�~ϿW�~� 
�P]񕢏{Q�C0�5ESG6�tIT�TDy�QAsb")�"�KNљ�)�ք���3DA�T�*&�h������ڒ��i&J(�b"��IA����P�Q�KEUI�rm���h���N�����` �"`��QLs-b	��m�aǉs<�5�
+lQ�D4�Pm�1M%:;sSMD�,���Z4j*�cEţDS�*8cQQ%E1�j���`�(���&.N�:��Zb	��(*b��$���b��1�n�Y�j�84{�EW�;���cp��(��:.y.��Q͊�1bAMclA�cy�)�z�*8mclQ���`�`�h�Ń��F�l[ci�j������ �4Ō���}ĭ����X</�h�J�d�G��5p@XY}�f�Ƀ�ԧQ�s^�F���ʃ1�9;���
�㯻��l,��	f���#YN�]���U&�Uf�"��n׎r������5�z�顉탿�񯱡�{%5	q��vl��k�%䣬�`3����	�4��Uve�v�m~��vC��ȞQ(y�CM~>��t]�7�1��Ϲ�2f�xӴQR���k�E�]�3(����퉜3���������{A��Ь����i�r�q0��ר_)d�U�Y�;Gd�r;�U�y��xM��&�vܢ'�<�8�^�D�c�r�[�Kx=R
y˫�I�C^��Fee�R]wxr�{6d��]4ɻL��K(�ީ�xi��e�.��!�ʟ��A�v�ʋP���4�%�.�R�1�{�_��mx6�LRsϩ�?R)��T�=���,5��"�1��Zx��1'�K��knws*��N\����>���(-r˂���Qi���_P�X�X��Q~��{�7I��vp������|֏(�-e��d^ϊ23q�A�8�Er̶�v���z^��J4�N�dh]��5˺v�;���h�2�f�L�?e�1_oK��� $a����KV��f}���+{��b���bIxF�]޽�M]6LO:��d"tؒ56#j���K��˘��LY��cQ���?z������d�qXE��j��Z�L��Z�����#��	+���\��,�.�O��ql��[���:� ���9�f�w{��9I����?�rd���Lwx�����hK��sԼ��b�O<�r�lG��qKw�B̳܉��[�n̘�	��;�x�"%/P�$Y�eta�tf��T��9{��B�d�`�7Y9-��<:����&�L�>��}ٳ��{^du���Bؙ�*����y�x`�c�ԉR�guS�����׮w�HcƊqڌ�n��B*���,Bf�t�ˮ�I���ȯ9�d�;�����Ϳ�,�������1��\g�e3e����>#BML��F�t�Hq+%x؃���/r�	��������@=���~,{��"R����w.|GP�����,��Za�:M����ŷ'"u���۱8��3$+\5�,�w=1�cWS8^�ҙ������+�g��}	�q"␽�=Bny�3hQk&"�'��U]�q{s�7]=�R��ׯwd�\��7?P־�G�.m%/��A�O�]�X�m�=�p��y��4��_l@Te��e�0��ҹ�:�����ț�u�Q��*�L��N|���V?A��N)���tC;�L���R}R����^�B�q�\�����3U�`�Ы�&̠��;�<2m]��!,sI�R��ZU�"gHK�E�hfu��QrZ,��O=�z�)�����*a���=Ӳ���f͚f��|i� �/�.�[��v�����=QI���(^�*�\]�G���L�U�պݷy��v��`��3�f�Jl�#ˉs�<j�k���QU�&�1�cP��.�8���(�r̡�����ZlZ�
ԉ\ڹ|=� ��r�g���uT6r��^�/�+YK9�'�c���?��@�T6��Xf,��CtR��qC�;��^���l�r!dt�u=��٢����9�˰?N���^ ��	RȩX +; ����d8��jnuS�:M#C�sͦԵ>�2*�a�.(Y�\��FK#�g�J�{g�CV"�!d��K����w^��>pj��ߏt-l�r嗦cS�������qT���6��;��/��r�ܭ^�+ʄgLY\r}�ȵ 1 �	�`~�}Nj��H��-��V�� �/qi����.��U�r�2��֎���,��1��{��8�-�bdx@X}���ОU�NL޸�����lq��{��.�ӣ���^S��O&�@'9OЎ"�T��*�XG��|���i����N�(�\�/T[���K:�z ѕ��2��IL+�1�c�/�iW)�l���me�ȃ�3�ީ��mK0Ar�W�� i�/���Pgohթ�.1JG�o<B�U���f�C.=u�nX�V��`�YmL���I���S���;�҆�D��`����ˏ��h��	��$�]B#�o�D�S����`ּ�ܽAF2�;�ۯWCk����#vKW��P|dXn(��sF��X�'5��ͺ��u�����&��"���[�T����-��������p���a+g�*�����w����u�Fg�1�q����S�\$J�g�R�mnA�D��y+�X�J�Ȱ_9<߰���__���=��?W�����j�L�^P
ˉ�l�ZĨd��!��Z�O���;���=��ַ��ˡU�wt�O���P�v�䨻U)�n�G��r�����)�������@En`;����X/b�,w9U2.sT�uZ��(qw0+�\'诒�ü�����51�H�s�;M�mڹ8dn��oQ/a�Jr��U)���U�R�:�rf���5a(!��z��uu�W��'�p�����/$3"�H[{��N|8���q渾\s@n^-0��(�j��6�^Y�i���٦3A_y�F-5;ڂ�k�~���T#yδ��]�9��r{�����k��g*�8��nt��x����x3��u�Br
��Vkݭn���Nvq@p���r��d��g��1���uw,���`bw�k3N��0!�S�Vf��KW]��u���jY��]|��g�qI/{����*P������<UcA0u�N�\ѯ�O��n��A]�uJ�"b!��
�9 z�������CC�*�q*"�UnoM��t�������ʀ�eV�G���˼m�ɚ�����὞�ʎW^Qţ�aY������ї�>f��&�K\;v�`t��0�ސ���A:��ڣ����E����^����E�Y�OgG�Ew��uE}�Paq�M�؂rq���=R��Mw0�so�kx�T���T>:�&�H&F2��ܣ#��w���G�f]���%ml
�p�l���V܃\Q�"s%��P�qB�7]_ne�w��=M�i��-Ϛ
���r�k��M;K+p:�v=.%q�����+�A��a�SQ�ً�	.]���Fw��2��r�D����<�}�s�^Wޅ�~�k��(J[]�c�hq��MG��bm�hԦ��{F���y�#,��z.Y���qV�u��x����'~�4��H`��Ҳ��]H)��zh�W��1ɻ(�h�˙@��%�"�}a�<m�uG<����np|ύ�b���q�s*M{i�+��ΙR��Kq*Y6F{f�ȱ�hE�����̠U+���.6�\5;���L	�0q��aU	�a�p��Yԍb\����v�Z�,^��d�P�{����ω��IoS��;ǢX�'�B���믪��O�d+�!ݧ�����}1'^�1_:/����u�[
���Qm�����)��zr���c˰ix�c�����s��y�:�\p1*�>	M�㼨_U�ƭ��
ݒG�6��33w�s��X����Y����k=Q��vQG٭�k1Eͽ��}z�C���x��y"˯;@ܜ�`h7@��#�5��z��\����i�de�0���d�OMs�]p�� ��슅^���ü&$��0����kz�D�X����]ьY~��t���^b�ݝ��۔�^�FK-��}�S�W�1��f#A���"@�����/�s�3��(��W΅l_=�U*��1O3�!oO��u�i���H ���DY3G�d����U���(j�g��jct��7[8�fhcu�i�J���{	d��=��N��Q�yQ;���8_���S�HvST�8�=�|3y`%�ۑ��K�%�X�o��
�-h������p�7i֠Ï	�T���@8�t`FE�ԇLU�lc۳��3���q��@��~��5܆�܎L�Ih�C0�i��TU����ە��M�m��̈�n#�
(�:��k�c�5%����g`���YG�+�Ck�l�����k᪹=#�Z�Zz�VpҩP�\�vE��f&T�ﳑ�'}�5�u��Umtlv݉$4<|<�� f )|�ٛsI~�(�;�o�<a�j������DC�!B��`��k���1���ED/BX�c�c_��Cڸ�R�d%u�9Mê�G�TH��y{2.�$��vD����1Cs,�?uR|�r�P��U�¡�9C\�����m%!��(26�Z��L�aC�.�h���9�{���������TE�r�v��4�~�
�sdIϞ\�U�1B��9p����Y�����ꄦ����N�lK8}��^������=ͫ2ך�U6�՜�����޺�$\#�@Ǐѝ�6hJ�P��f��:�O�\sws��X�_(N�z��=B���%�����i_Őn�%�=��U�� ���!����5;Q8`�\#�O���B-it�3��'�e�ؔ�i���̓�K\4�>#���k����nR&���9yT���e�i6��afa1K�*{����(s��P�Q'��Qt����k6���S]��;0�i[�[u�>�MBq4mV����,��s��**��H�����t ��]Y�����	Q�Hs|�4�=�<l�2���<����.��Ц7�Z��(�9���π¶�X�k	��Wh���*r��2�ٴa�	+K]�Nj��U������N�f�Ud$T��c�BIW���!�4SU`�Ʀ�����{��f��:�6��+��k�����K�Q�w�pf*e �j9�?s����qn�X1.��k.K�U���,M�l� �A1�]��cS��E2�E�YoJE�Sϑ&�O+7f��h5���Z�UQ�]�f���2D���Ȩ����=S����f6�uQ�׊������ossVƭ�߯/���xZ�^�[�cϮ��di�?y����@|tS�ދ=�r���Vg��5�f���~�^z`c4�T���	��ш]C#�t��)��\�\�=�Ϲ� ��s��B.�zn�4�4�6�������#\ц��X�Ul%V�
�Q�yy��,i���l��*�jz)�5h�?o[:��9|}C6�	�����[��g8Hn��{�Y��.��W����-1k���`X}
���z����}|��8�3�sWP�Y3~hƫս�b~_��"E0�ʈ~iwưL��,�0c��u�ʲ'����~z/�����g�-�_c]&ojG����*��W���=��)B���'��WjB�%ڠy�r�p?}���)�;]��'FK|f�ݞ �{�����&�=K�����	�RΕ��s3�rm�J�j��_z;�n��K����p���|9~�y<{:T(y������[�((.�td�3�Rf9��=1ZY��{-ٻ��-�3��l��]ЙGj`�Q�m���N���x|�  d����)�f��P���b��S"�4��7��^�Nj�b?Ed�~��ֻ�$�{��dN^���� ֦3#��ݐ��|��'LK���i�\}��k���m�Ԋ�&ЃZ\���~�u]���x��p\}�`/ާ�yu:�?O��a�=%J���9va�D�����NwZ�9�J���>����'�����,�ל��Մ��*�o�g�A��wF#�#_#%8�e;��_F1r�}cU4u���A]�uJ�"~��sf ��q���u��p-���KA�8y�y���-�aӖ൮Q��lsJ�!O���%N�h]E.�������5�;�L�*�{ׯ3���68�ם|MH��[���A���@�zB��C��ݝa��^�r��iq�ν�Z��[v:l�q�]������*�D,�>�4�]��g~�6���Y�\,n�i��l$t_*�mu���a|��7��}Cq-_DP0E!RVa@6��行�od�����~�!3�%���
���dv�i�vf��k�x*�*�����^]�����e��3H��eoR��'�QV-s]�4GA�Si���qqN��G:ߥ��j�a*�>�����߬z�ש"]!�%`�%yusK�Ͷ���x��|o{����ۓ������s]�n���Ug���\ʗc�f�_����W���=vE��9�O8��F=x���Hw��'���{����Y/�Đ���z��*��WI�r���0r�O��t
�_��v�.u1�ƪK(�~W�ǯ��N��槃�zxͤ��s�~�{6�nk�5B� �K'��L���W4�cV���
O��<m�Ͼu.�:��J��sŴ��hg�8����Zm��W>w�����"�Ie���8�͚�sp�ϐ/bB^�9�X�wu\b���1LDz�>������\<z����j3iθ��M�x@�`*�[��Q3Sƽ(���/o��������=��P��c����<�>B�%ֵmǚ޿�:��GY�UT"�Ʉ�f���/��nUnG��U��l����F����(��u���$�b&�szOk2���s?)׽\h-N����w�k�!Z6�x	P�P���P��=��w��_���}+'�r���!��[?��(������R��c¸/��U��7�.�^=�Ӽ���릺�%����#mH���4a̺h/�K�m1����E%t�RH��W������4��<CŬFmN��ټ�C�r���v-BE&g"(-�����"�gR%u�Z�(��N�UA(ۙXi�p6:۷�ΰ�5���ͱ�����^�
��w�Vv`F���ˋH�X��l��,nc9:Ԡ[�4ck]��(;g�����!W���::�%E��6N����fN�j����*SS�geҭ�vۮp�s�blCe�A�)]��������$�j���V ��W��5EȞu����B�Z1Y��|����"P�::�v������6�Y�0{�	G��n]u]��)�o]t����e_ɥy[����_]�vΚ�8��pQ̹P�msޖ����E�	Y"�ړ��әV�f���s1��'a��Y��V��*uӬ���ݒsu�N�}��♈мAE^z�gL׊��]����� �մ�qS��F�9u��[;V���3xI;�;�L�F;�����B�(CQ�9��cz��m�6������5{:�E�5r�oXˣV��͆�����#��I�-FTɊ.�hݭN�x\uʖ�{��r����.i�.������3�(*t��ciqgj��;r���S�7k�Eٻ�K��*6��f�u��]�3F��[N��6�"���M�}�`���	�&�J���.>כ"�#\gN7��ַ�F�f���0�w�cGo�{Ky!GGlR�Z�}�L:�L��̴xc�Z$ulэ'���+���2�hRm@�T����NU��Kgc�f��X�����͸�g�_n��3���>W$�8o  r��s,�����V�07gf��[L	6���`v�JYEY��Λ���}��]]�(%�X�z=�������]�]�;f�7R�m����5�E���fk�b�P)%�.�Z&]bK��
�N��
Tfiq^�wP�EO��XD"����ȭ^����0[�����\n�q�e�ز4D���=�]ng����.�y�v�Gr�^�Q�$�N��Hp݇�ܮ�#w��X�[����^)]W��w3;ITt���� �-*����W	9:භ\ovP���O�ׁ�7�A��q4:��a��n��뒞بl��MB:���������O�� 5KhJ��[�����|�E((��J��z�6��M@�[�ͣfc~����\�ʍ@A�^wU��sʢ�â��]�b���7!��Wc]}n,�غ���N�!�q ����d�ū�v�W��>����I�˭)=0^>T5�rX���hJ밊f�:T�V�ќ�Wq\�8/#��6�՗@J�����d�rA(��*��<�mb`��[b�wg	�вƯ�-�p:�3]��Nqt��+p��.����v��]�́��z����^q�˵@FRـ��a�Ϡ�ȃ�q��1���m�▙h�v��i���3[\���@6�m�$~�´-ˣ�H�E���/a��zY}yA�9���7T��	 	���$T�L
 ����&��-8�c&�9jj�X�Z��j����6"��jq���UTUQ���z�{Ɉ��	�	&���QTS�uTw4lSA14U؈*������l�SF΂6���
�i�������jMÜ���:����`����<c�~Ƙ��墌Z(�Ţj)�����*��b�F�G}����ª�B�剧Z)���(���)��RET�E1����Q��QQUEw6嚠�b��#lTEW����b!�*���

�);�Q6H�J
��j)�&��)�(bn��|�14D�DDR��LTN�|5{>�k�����p�UU4��M��������)�"��Kd��UQL@L�EEx�]���ם����#�˲�ǳ+�v@��Wuq��Ue�L��P���[ϹJ͗)7҂���8�sr=��J�:�#{�=7��ﾯ��a��SX�nPˮ��K�?�=��<��B�lb�g/K6}C��5x�=��}�[�/�v	����᝾�F,)����K��1�<�q����'�(���ZhF�U����rb�����Z��{D���:)=D&�*\��`�]`\}}9���j �����۸�7&"0\����<��4��c�}�WG��T5JX��N+�zBg��l���?0��W6���8�bVe�}ק=	�iS��ȉC=���J�5j���(�B��"~c��#��x�UZ��7��W7�{fzC�n�L�{�9�M��Y2ߪ
�s�N�>8���O*�NU8��{>m���gm��cU�x�/.C���Ph{a��S�,��[���p��>��ZLK�(W�)�LM�����N]"qz�~�~eH���R�� ��T�~�+�;\�SS�;�;|z��:V�;�٠f�P�R9�ś�����%5�G4�2��ڡ�4;����n)���|��ٯTLI��8�=�j�p�c]f!�f�A�{B����3f2�;�U�Z�d�o
E���M̰��Mpqz�����C���<��s=qX~�ږ��Y���sy<&��l^��H�9z\D/�m3��j�^%r��Y%>�Z0|�VVC���Y8rNޝ֖�׳�̜E���8ш������f��-��7i"�D�]w\�R�-���ݳ�<<>o��n�VT>v�ǿ��@<`b�z�.�n�r��z��QJ��1�U�����y#��E�#3ݒGn5L��9)��m?��ն���O��<���Pզ��(�(��l���QL�Gv�s�o��:��`+��dwL3�s��/�'��}�p�	�a)	��ԡ�oy��%��E߽lؖȤ�α�o95�2u�zͪ�2Ys:CĨ�&�����=��;��؊if��	��1�P&S��@�l]�T���ޥ�*,	��|l2Ξ�粚�k6�'�PoM�j�Ds�P3�!8�z��jsb�ly���{��u���i��!�u���{�����Q�C\Y�\H;�k� �2$@X}���{t�dת��O ��R�j&�.�Ʒ�q�h�Bz��tP�=C`���_@��|�/aglc��je],���	������v�}��·��`ށd��3]&��%b��#��C��Wi�����Nlnın_!Bj���Bn��n�4�#�o��R�`��i�>� �0ܰ��t�~��93Nd���B�x�g�NE�\������t���~t��ܞ'9rQQֽ;��RZ<j	W2�o���h)[��i瓙�\sV\����z_c�jd���4x�Ќ�(n��)�c�p��Z��qNp�h��'���<�^>�<<<=�xxd�E�ɿ��?��c�
h��Ut]��Q���;�[��IccoB�%	]����M/�6�c�3����(/n� _��lj��㼨Ji�j�{�:|1-�ôvv9UFs�Z�.(�f��<3�W��l�+]�;���.t��s\J�5�ˮ�6n�_���p�#����ı���{i,�kv�~򴞪J�Eڹ\Ҿ�p0��@��$�|��,B��uGmBn�U7j���h;��9�T��1�bËf���@�O��-h�	�Eګ\|<�h=G*E�9�NXZU)��Um��_�I��:��sW�zR��~�sE^�b������и�g}�d-ޗ��;�I��.�m�b9r��C*����PS�\X� �2W�B����E�3�;k��E�oO���"��W'���삝	�*���^�;�zb�^+��$�9����&4�I��(�2wo}\m�\J#��p�ܪN<�Oq��R�n����i�q�q���Q���0�`&����10� Wu�(�9�ʹz��n�W �r�h`8#?kh�w8�]k���lw�NU��I����ȉа����9��2�I��GQ7�o��K��$^jx=c�q|�����X���2��Eu]gKR#�'w����-E�e�m�ޱ���p�KT�wj7v�N>c�|�<��x{���g��'W�kC}U[X�Usv�Z.�W�¢(��j��(�"�ϢzBT𝇏�f�\8]^�o��s�59G˚�U�cvF�nϙ̮>���Tg���G��>�.,�G�މ�QUl]R�Z~�';�0��Rc��lt�M����E��t��è��:D8��cs蜪7���Ph`��#�Q7�v8���4%������t�x�����֔���.���/�ng�����ւ��5V�K��cqA��{�n�d��W�.��/۸|�'�~j�٨z�Nt}�����_?�#ǳ�Ω�LT�:
�p(�z5�ʏu�i�"	�X�St޼�8S|p�UOrD���^���Z��%�o�F���1E�D����z1�9R/3B[��n�3�:V��k�#�˫�{�wB�ka��yĖs�6��;o'U��Pg！�]z�$�8���������C5��䞐}�q��~j�{Tv-�-<Z1�5��I�Nc��s��%��B����=�fZ���w���8��j[�r�Ƃ��t��a��9C�ſs�5����Q�n'Vk�RQ%p@˝��Gpr��ٶ�7ļ.V�k�S����r��T���YimƤ�)��(�4��w��7����骖��5k�����MÜ噘�y2ՈZ9��)x3���e=�+�u]��r����2NW��*����� �y�� {V�*���5�5�9��Ja���S^�?����ƫ�9�dn�~���ᾣJn����^;�ax�V>�r�y�,�ЪD7qZPv�ή�%W(,4Q�`�7Y�O�Z�{1RlS'e�r��z�Xǹ����+�+ҕ�hh���U��7�u?i1�];>�!���w���W��N�/6 ��cz.SIu��X�ϢЊw���;�`:�yR���Q7�����!��>wC�/产�y�h]��Ra�1O3���g�t)�dC�?�6�Z3DY��|����GP�4���2��<jW�m�U�n��Go���;B2)��u7�iC���^�����zS��<j�A�$M�Y�
��!;]W_H��bw{(o�ܪ�ȭ���<Yv_�&3�H�=V����M�RQ� F(N1�_HL�Y,�NsI�튚����Z5=�Y}J��G�'Џ��~�y*0֘J���φDB�a��p�"�T5_�^mLmn�&|�����]z����6�J�7��k���^��8����o�jx����F1tŏ�����J�`��wS}�f��:���.�I3���C�u�oX�W�Fu� �ђV�1�aR޻���V6�.�;L,�z�(��W�Z�1�Q�M��G>�v�D7/r6�hº@)���u^�n�J*�c{�*�[Yoy�
�)
TD=|�u��v{D�����^�ŵz�m��UCг1����xk�'(>���oO��R'.tj�UN�o�=yW�+�+K�`�Ȥ���Tu���0��JW>A�9��턲�iξ�� f��q�w�z����T+�Dy�x
�_�~�ɷ����oGE��4�&^'���B֘>[��{r��m����7hVc��=ix�����4%6�.$�"��3~w�k�����f|���|�m��� �g���ˍ���Yw#5�nWX��"�܆�V��7�Y��>��2�,�V�Fކ/��	�͞���eX�2��	O�i��&r2+��)R��;;�5I�½UcO۴�p��OΏ�0%0sU�j��3!H��2(wT��XqS�����+��B�ƘK;��v7�e=�܈r��77�֗^x��R�p[����7ɤU&�8�Jy�$d�8�y�{�^�\e�Y��r���5eamb(�d��õ1�Й��xVO�7�B���q��P�=�%�2��E���x�ld��;�/=7+W�|V�LQ��&cS��
uQ�E����_�7��G�IR�7��9����d����F�ǽ*��WA�|�nk����Zk�#�{�^'	�!wd�YW� �z���Z�W���)f �S*��3��;�1�Z�r����1�Мh����q;RW|���ҷvBmGF��� V��d�ͦ�jqw��H{���o��=��y��{����l�B�}��f������J�:�8k���r �J�qG�oHRC"`,>ܿip����i�[�Z�9yXZ�"��M.���Q�xtP�=[ ��0�"��(D���?pډMݧf�媗@K����mӸh{Z� g��xY�{��>J�5�hu^�X�*{w"$k�Bq�T#3��1Ӵ��n�D�98С5s�z�/�ҏn�4��Z-��Jm�<ud����X��S�����&)0����$����m��^�E�]�rn�^�>�G�w�U�������cj'���>�U�B�#YMK���ؙ�1|�*_
^��]p�%������a�e�5�]� �f��߽�οC=��w�D�[�R*����#U%fB^>2��mp9��2&HJ[����E����^��8����SL���V~��w��<�P��+I�&�%�xzZ��3X�|�pǳ�k�2�K�!��נls�a#��c�䪙s�QM��+P*/&^4Rz��n�z$�<9���sV���Q�N�L��	k��WD�,-*��ؕ[u,���*�!�S9۞��D��Z�W���7��,y����:9D�R'B��]��f�^��7�~�ۦ[������V���sn3��V��}Nj�"[�t�P��ʵ�l%b}��[YRv�pO���w4�ˇq���aVA�e��L 
c�ۨw�{�=����y��ET~R(P"���T���Mr�'��A�v֩���@M�����6���Ғ����7��s����%���7��%����l
�*>�"�_N�Ŵ.$��]#���<8�rd�f�z'�fCM��1�Y�>�?f��.O�R����ڞ  Y�z�zTi	&sn�NQ�ՅJ�>ۇ1�x=�u6��cy���[�4�ȸq�^J9C`�P�in�R\o+ʺ��4v^KD ��8j�|n�B��4�8�5��8�Xq�z��L��Xk�ܣ�t�Q� ��]���Pg39�>��aWB`��j�d�w�L����o�:Da��q�hr�<i�c�ṋ�b�Y]��o�:��qL�����F��)���`��{.�
44j�����T���a����֯]A����hY�%F�fL�q��8�h����w{%�~��/�o�y�f�3����~�&�A�7�܂虆�T��~J�^���/lj����Ǥg�i�CWR���a��x��Id7��MN�J�����(��_����9/e\�=t#	tR@}��?�wM�w��]L�g;�:���4�6����a61�t���,d�z��w��,n(�uؕ(���9\ƩqV��0�mf�h��p��yg�����1���|�Y�Y�4Y��Q$�^�x�[!�)����Pf�xxx}*��*Ҡ4 �u��:�ɱZ�=/V�Íc^Ԧ�^8���T�8���~�6���q舝T��T+��n�޹�α'�oB�"�r`r}˫���%���0Y�8��y��8�͚�1���9_B��1c�ݟ*���Q0|�^4���N�r`�t������`q�N�����9P��×R��ƷaFw#k1�{+�]K�f�;����ʒ���r�46�b�a=
Qqc�U.z�Vs�)��7;j#]fteZ�}�WQ�a�z���?�ςQdH�f~��-ez4�ͤQ�$%�$=d�Q�\e�lwz�t�}��yտH�ޡ���"����+��T�P���7+���.�ηK��(��t١��|�+�����T9�P�@�6XE�O$wx����9�[q��ӾO��u"S�(�|d��9r�Kߒ2Yn3�A��/���֮���عt,J��F��������M�!��|�T�|����{�EQ�V�v�mN�c�Z�xQ�	��|��Oc66�ٚ/۪yA_=�Ɉ�`㊐W5ƥ��~T���P�h^�}Bΐ1�6�����Uw
[3�vUd���'�+G��M0��j�ظ��04���
�L�w��f.T��z�|��8P� �e�1HF��"L�%����wp��
�c� ��������fL;AdzZ��:]��y�bfR�Ѝ� ����UU��J-�J��P�@�	B�Ju�o��^�<ݾ>6�����uK�Ü��"n>+5"m�6Hu�hd{���X��0Mi�t���^k����/��)�Ffˊ,L�5JY�����R<达��H�q�\�>��'e�'_�����tN�r�rT7��C7�0�j���@�R�Ȏ�־�YW4�./�ձ�j��^��;�l/��QfO2��L�O��[����$����NLE�����W7�G���Q���Ⱥ�:��/X⚅��	g��w�fcC�A��R%��NC���]�D^�B���ǎ�g_m�Ju�%��sd�%���F�)ޟm�v���H�=�ŕ^��)���g;o�c"ػc��S��F��d{���b�����[�PS�f]kvC�me5}��>�X�]���{���cN���.srEm%X\]ꬹj֨��?Fw�٩\���ZO��4�)�]�U���&�no�>��(L�9��{��=�߽#3]�J�X��!]�\�Z��&'���H��a�jԆ��2���"�<B.��c�s�O����F�f.���ހ0 �0�cF��+���5��}�l5q>T��&[��e�\ks�|�pҜ��h+Ǧ6�)eSN�	k��-Z4�<�D�Y�G	3���W��n��}ؚ��FΥѧV���g#��sb�f�����G;�h
lҰ=�:�V�c8mq��p�A��$�{:n��#��q���qLϵ�.Y�-�蘪ʂ �M5�h�RrP��(uh�
���-�N��u0h���Zz�R�,��g@��aT+n�\}�I5RWZ����9XP�Jvt��[gh�4�u���1vT�)�I�+��jr����#mlnv�u��\�>kV�zG�N���GF�Z���i1s8B��,E���FD��HrvZ5�)kЭ
ٸ�-�}(6t��٫�fŝ?b���@�fڱ���qؔ�2�Щ9%J����h�Z��Ց\��;z]�-��i��ي�ř�DKw�.k=�"{�*0�n)�����V�1ʲ]%��o���M��녜�لc�t-��j��K[[�{m����i֛��dVAQM��e]�֔-�\o��	׍8���r�S�[[S[�G��ksr)�"WJ��W\�7� �?��ۦh4�8�&z��G���ұY���**�ة������Lj8�I����;x�⇤��1F�^k�Q��?��m�(�u�J���&]]�2���r�jq�5�*��E��pUZ���׸�cV7D�{��a��Q��=zV`��$%����c��Lk3&�+����d��7>��#طZ�M����;�yn�dt���z��ܷ��!N�B������t��g!k^�]5C{!��g^.PȬ�W)v�'s�	:r�)J�Vh��J�2�@Y��_Ԫ� c��c�2fS|J�e@&ꏞ���+/�V�A�f�Z�x6pVw�i�i푝���ۅ�P陣K!�.�n3n�Yb�\B�NQ-��v�,��t��f�W={�u����&?�ŨKTs���N�5}����V�Q�{[M�+a��/*\���-VE �u��͹��M�.��u<�����Yc�ӹ��������}fSm 4�ә��^&�᰷6�����J>�_a��N���w�MrK���3{|�X����n�G!��T�Wk�ls�9����粻�}�x�Zk�ER�2������[�D#���eEn�f�Ճ=�m�7(�C�F��`��gb�a0��ɺ̬�!΢�[�X9�̢� �Q�o�0��=����,�N������*���1#H1|�G]b\���"E����,�S8����|H�'��yKi�"���ɻX�����-�Z˹n>���7w�m��^�N8�����*u�
�a_��	�''v���v9�73M�8%e�o���L�KF�^����:�	A��t�-R��$��z����%���2�^�"9�ɗ��>D�I�i�u_�v���b(���j�F��QM1R��h���"��)i���y:��.l&�17ch��Fä#gUF6j�KIE{�#{�Rw�AA[`������f���'#E�
��cESACAUE!TU)E%p�T�@PDT�@R�RUT!�U3SM�DMSA�4PU%	AE-@RRPD�-�L%�RS�iZ�@i"ZB����)������9D4!C]�ĭ%,E-]̚��*�)�&�K�@�QQ4�W���j����7�J�R��!/���K2	<ס��Z��Ճn�Ϗ.�N�^ʹ��L��h*|�)	\�4J�c��nI��$�h�v��^.^��{��=�7�Ъ�E
PF���F�)B!P�D�h�iB��������9��~�_���Ϟ����S�Ť=�L8�Ŧ�8�жt�p�
��X-n�����۲��G��)q�*ژw�S�}ɤU5�,Ҟa^K���^��T�\��`��wnU��=�♶��t+;�%�LBc��G�۽��o:p�(Sp�\���Z����w
��<�/���B��ft�"����	��f�1�w�(�g�V횟�씷]����^�e��R�C�4�S������r���@�b�R�8X0`�D�?hz��Җ��_�=c�\�
ɦ�5�&����q�q�h_��^K�x?[�cκ��UVF��x��cue�|��/��ӈB��^��b�D��vr�aԇa[��ⷐ�6�S5�R>0���d��xo����"w0��R���X<�;"|:1� Mܽ^�! ]ܸT7a�yx8�Wό�����\�.}�u�[��îH,74b��<!�i9o*�������+ȫ뒓m�M�Y���+���n�����/��?H��3��=ޤD��F��Q&�樫��i���=��d\�
L��བ��U)2��Y�s7�i���tM���tk���J�oX4�{�PH�����@܉�c��P(�3r�s��t'k��U��Ts�.V�q��j�b�p��j}�'��f�kӯQ���Kk�9"�a�us0i�;%�JI���￯��� � �ii�(P�h�JAJA
T(�"����t��57���%��*	�L���
��?c�>���T{�՚���i�Q�;=n�9���k{�.�}��slJ�����u�om�,]��x{lwz����o�,�B�o.6';u��NU�WW!���j�#>ޙg��n��]cT�u,��T^L�pJ�iͶ+�����6��y�>l3&��צcϚ�6���<��X��B{a�*��ؕ[u�/KΕ畓g՗~5�+�OT��:(�S���k�nQ�S����3��B��iҢ����]�gn���;�U/�[����e7_�,~j���_`�;ǌ�_�=x��D?��i�/uhY<�=SC�X�ŧ�m�#uc^+VZ���0H)�R�HI3���Ö�i�Qgy��r�΅m(���ׄ���p1tPn4�-qvj�����vB�gQ�fCyٔ3��{iv�bT��r�鿣6h�޺���󯉩��Z[%�ц�UR�&�yW*Zm��\�Zܐ���bQ�|��Y�vFvi��3��z �H��S^�|�jT�4�~�z����Χ����b�ؼ[>��t�z1��)o�.6)�Y�����z ׽^���d�+�����}-�36�p��E�ĵ%�n��VJ�^;����R�������
��4��V��6��^ۗ=���{n-M�TX�����T���������\*���n����}_W�R E�(Ei��|o>�>�q3,�F�>Y�DA9�!��r_*����~9/�8�i{my[^N���-�r���:����`�I�PM�����/�P��o�nP�=t�&qӉd����ܩ̦��[!����-Ϛ�f�R��%��PdK�j��Y녷���4�F�o�����q_�y��i��pO�i�{�!O��P֙KT��i�Id���U��Q^c��^��ߝG��6k.�q��Z���FK6�%sX�j�K?rĭ���zq����2�J:�Y#�:i��Ԃ�r���4����fE8���>������>��B�X�P�c%6*:h�wt�	g�E��w���#*!S�] �&R2���ؓ����%�آ���s�|h��ׄ�ܣ��ͽ�������ވv��u��^,�/~Dk���=|��s�E�C	�U�Ր�M�tTY~84�o'kPe�?��=���g�:Y_F���tbyT��n�&�t�h���ei�D�<E5y`7C�PX��X�t!�xk􌚈�|:�y�u���}>� q�ʂ7Q}7��:��y��/0���v�n�8Ú��:���ig`�N��8�d�Fq,�N�Xq�[�U������9wK�<���
�T:V�!�����ٜ���Kq]ܻ�z����GK�ݸ�W}���(|H�P� ҁ�^:������](m��65f4;f�5,MB.�x�#n�>��RP
�,�F0x:�(�,�Z�����5	x<��y�&�D���E5z�ɇ��M%ב��s>�hE;�g�%E�e���t�y��$a-�dHл�Z�+�X��|8��rȷnt�Tl�/��&	8��uҷ_bL�a���P�"�@����G�͑��^׽��=�Y�a�#���N���+����Sq��H:I'�
�H��rZ���42=�g�w�#�]�U(lẀ�V��Qu�7<��c������p^�G>}�RΥ �-dFG�F��'J����g����ϥ{/���������g�}�D�����_���YT���c3)���S*4��B#"�!�=����j ��q�P�q�⯟�e�T!��&���B��Y��}�|�P�<��ޑq���mE�k�A�����:���(`��\�7W!��yzT�^�Y.�{Um��"~��8J-;i~�}󫴧��g�ULQm���}�D���ܛ�������g�}���&�����R5bWK�U�/M����o\�kn�mS=�n���1��h�N�b�OXs;+f%�����hY�5n����pgQZ 51�^�#�$�?�(Ƿ�nd����
=MU�r��v͜۞���}� ����7�����V��;�+~�a- ,�xy��]�~�Ò
�_HQ�MS���9�ꓹҟlN���bb����Y��Y�,��R~�r+7��b��3���c���;�l���,�b��-Wo8�g�u�_hT������4Z�bes�x��㊅c���>����B�$$�Wr<��Scn�k�^n�
�^NS2�(0d��u˥�fM3�.}��>�r�����+�S[c[��j#��u^|���j#�<w��\꯭J{���¼MJb�<�e��y���S����\�Ѹ��q>��jGE�J@LQ�%_��\_a��<5�:?�k��^��(Y�\��ֲ��u�C�y�؜��ן��rȐ��çD�v�,����>z����6����/�K�_,�{c�wj�q�����A��-X9�� `�V�L'���UF��
�)�9ԓF���U�0�2~Wٻ�ln8��y�2(�8��8G���Y�C��Aސ�x�C��b��(90U��ɧC,�钫�meS���&/\WƷ�	�hǃ0[P�cY����q0�4v5�
�g5�;��em->�d����aփ,+�;�t��ڝ©
�{��
�:RU�����IÆi�$*v��v�א�T���e0�p�Y��>��*�����Γ$��b3�����ݽ�3� ��4��OviY�5
o�����<7���u�`߶S���"g�kԣ��������#P�+x�ZWr'[�gr��S���9������IX���a�H��8\W��J}f����R��r��_8��?iJoM��eC��l����l���^D��`nT�'C"��.8���[�=�Vj����c���<;F�0���w���O�=��r��"m��W��l$o���+���BP�^���9;X1Dl��x���MHiUMͅM[��Po�*מ�U����>��Pf��0�Ǐ��(fwCW�T=��TNaAR����kwB�c�T�~�b�O׊q����d�>ݲ��p�����fG'A�/|�U���c��ø�V�7W#��<���W��,�[uE���>;Nw��NRr������&�[P��a�R7n.y��d�Хs�9�NXX	T����-3����{�{�r��j^�+\ߤ�G׍@��>��R�u��_;����4�����-�8�5Ȭ�%t���Ƚ�\�"�i�{5ds��L4:
���V>�U�?{�8��&iCn=�	�M:'״?!blp.��E��u�����mu�|����Β
���:���xz�m"�<�[��#��aN崨��]�.$Z(=�ekƖԢ�)xrRS�Z��s'n��ƴa�+K݉�uz��V�Ϣ���oyL7����_2�Y���x�!��?���꯫>�2��v�紭z@�\��A.�ӡ��VV��% ���C��Q�]�_-���^�*y+pw�~�<�Ug6h׹��C�'�:�\u�����'6T��z�[=�q���8�]ɉS���'�f׎�E���x�ם|MI5Z�Ų]�;�2nn�ČLk���mhqI�P;ʥWʅ�jb�hi�[��������;���j�9�̽�����2�ݨ)a`pG�NGǣ��Y}�8�VM���Ch�H��(�"��,xwȩ�ᶫg�ۺz���4^���`��"�(|M����x�҅���l�)f���m�&�XB4gt��z�Ԏ4�|dp���4t�CZa,$�2���^��2�#8��BL}���"=x��i���h�ʩj��T�T��^��fC�)
u���2�<�@�[u�#�t��3cR�GD�!,������ώcŰ��IU~��<JR���W4�av�0�QqS8-�͓W��i�����|��"�ђ)�_�AO>˫�lwD�{�2j�,盺��	x�:rhR¶m�(����K�b�\���^��~�cn�C�1{]-�nX�)^��˞���ì��(�o��[({`S
�8VJ�'>X��u�3.CD���c���K�ڵ���N����q��7�- ��'<_��&���$Gg}�{�/�|6�䘆����;�CCܙ0GC��-.�D��|L��i]k�SOUTѫPdm�=S�y,lnT�{���I��n׏�����4�����}-�9B�A���t�G�4^l��Q�>2����A��;O5Mf��W���-V0֠NNK�;ˠ�Ä��Ã�sZ�[���{�!z�xvմK�t�3�7�Ð|�E5�m��U�:L0#�V��	/�.�/P�����9����P#�dyA�Pٔo5��r���>�a�Z�r�\����_��jVP1�˥19�!�
�FT�z�ƭ��1|�[X�Mܦ�{�,��y��q�Aչ�S~��7Z�@2�N���RE��	դTto(1���J�/n�`<�0�Q��9����=�Q�b�vۍ�E-��|}�W��B��Gf���.��~���Mx��o�$�TF��ވu
C��w���wr�:w�<��.�Sj�Mg܈:`$M�+5#![�5!;\�����.�S���͊���}X������P�cN��d��36\P1b`�s˼��d���!���@#���rwVtXQ���9�]�j׋�����v=��y~\�__����NvjY>0]�Ļ6j�׳D��{�2r�<��P�E���NJ��F���K�!k6D�S�>��df�K6�lH�m��P��|����K�3D��v�8Z���諾<_���~��=���f�2ݯH�3�o�(�%_oJ6���]�V�K;h!��oEN}�HF:��Ȉ1�.&,�/X��}[SqPs�C��m=+����J�;`�ٍŘ�Fz�+�c�K�����
aP�p=7����~��[��� ��6��������Q��~�(_�y�%�8J���R_���Y3֪3��G>��|En^����e�����N��R^g{gp��M�V���Ь���(������V�ǈ�Yߏ��E���2�����S�KT(�mk&.{���a[c;�8��o\�
�vG�h��i��;�"��ʉ��������l���p٧׳����&�X�I�F����+^|�����}�>��}���(0�r��B�mj
	��.C��h�C4�)E�.�|���|_.k��/���7�z*Z�2e�No�X��վ���u��LߑJ�:{V��wUZ��{�Bυ��'���j�*W:��Ј�ɷQ�j:�;���5-j@��!B6�N)�R��*���V�T���*��q��F:G��t�T�f���=��u���{�>j���]b�2�gaέ��xbz%d�R�d��o.�2�:oB���;]+�a�&m�TE�ŪWu6�Us��*���t�X�=�hGNbux��֋R�-'v�D6SWc:�O>Nt��m&�w1Zo3D��� �5��%�d��������ȱ�a�<����U���`���b����VϹ�T�O1\�<wp����5ĬÎ���W5�P���9
M��_r �J��ZA1�q����ڠ�D�TKT����q�^[_vKy'�¤�Ez�p1�����ׂ�_���F��i�c����]��8E�5���	����.i��������9�ɞh��0X�b���TNX��qy�r�;	��:�Dt[Y����>;yn���/��r�|U�ɫ�G��Y>�5�V���v�Ra]tIX�D}��2��
j��dBE�8S���4�]�̸�A�4V�E����իK�ZG	���#��Bz0���&5���N�ϾUuN��S�j�;��YH�ex��^��^��vQmƗ
�tp9�@�=�Bu����l�7ԢM�sV�# ��Ls�Ӿ��;U�[eձ~F����-JAeI]
ǰ�^EPŕ�6N��������ن���qnk0������7�5��Ư����#V��[{
��D-���@� X``{K���#A�J�ŘѶ�xSm�n�Pz@����x0���Eɼ���(�^B���Y���E��
��r���bS8�T�F�l�l`���yR�������[b�n�@5�)¶��ڻd�5�M�/��ݦ��̭��bu]�d�xYˇ��zV(r�3��E�d�f������u�/�[�B��]X���F�<T�G7�G+�+xuխ�[@ga��3�������lh\F�1��+5�ڊui��j:��ϣ}�gQ�2�g�H��cKhP�zK�
L�
��`��*�ܝ �F@ݴ���n�{�i��%��>���戳�NpGi׹h3����e��[��u���X@c:c��A��QrL'f�>8������Tr4hӱ�%�
b�_� ܵ�cOku%VT��d�K,tx��+�%���٭m}�� vZ�O8𽋂�D��[��q�[G`�lM��Ү��۬`ڽj��p�LN��[3�FT��_'{;\V�K���Mn��?v�G^��l���0���u�s��ʻ��*��n텴�M��Vʲ��� [t����[�c��A���u�E�*#ս�v��w>�+ K�S��r�0�L:xڸݣ�F�p�u�V�^��j�By����#�
��ں�W )�KuK��jnD�I�8{vAP�i�]��Z1R���Gjj��7��]��V��:��TT'(A��'0��+���|�s�ӥ�TZ�]i��\6ˌ�W��3,!����ڧ���ח[�NS�;���SF}u/#��:��Ǆ$u�_��nn��:��n ��7fY��I� �upN�S���zL�h�+��Zzn��Ls��N��/+6�96�ۋ���f��)fؒ�[V٢JĹ�mo۲�����@�`M͂WH^���	=���v�*<L��=��6��9a��(d��>w����u3���tI"���|���T����:X���ۗqU����Yɫ&�4�힫!�ȀD,y��}']	��\�Ӱ��|��1
�x8%�tJ�!L�Y[q���4r��(�2ѻN��{�8��v�ܩ�P�eī�k��s�1��K�.��eXd�Z��*�-��WGS�<p9�oR����S�J�j��j�x��m���p��fcd��q��Ρ4���ڙ`2��[-�n�5sBֶ�sW��N��M�sW�|�
���՝��Kqoc	2�Sy\[իn��!�v�r��f�����K]���u�r1:��[	������ږ�����v�Ӊ�`���_4z�7u���D,OM
y�]wN� ݗxS�'3j>t��)t=ĵY��/�#�%ܧ0���b��\~鯩b��Ÿ���-P�dXr&����U����*J��	w���q��3m���C6)�N=�>�zΌ⊯��d�䰫�X8&�aڹ}��-ړc:��*eɼ��cn"��W%��ݜ�Eq�pN����҂��������.[�L;l�Α��g�:��B�+�Ѫ�\{�k������QUT���D�FçN��(�&����i�Ji)(���*X�4�IKJЗk�#AA@QIKA@UQ@rMPSHЕTS�ETPR�rPJR��+Q%-U�i�(J�h
��b��U�@L������$�"&
A�b�F����JF&�JꐭН������&�a4�Gx5TU
��9+�j�
�Ji()(iN�a(��<����2�`�r{Hhn`ҳ�x3���
oe���]	
]8���\,q��&V�'�i7:��E4C�(���ҸN�}g��"�\ґv�xls��۾�` ������+���?�Y6>��U����s��XH�2��%T˜��6�d�l�zfkߋ[� ����yLj�ִ�;ҍ��d|�U����"�>^J�3Shh�<�r��+S,ש��z�5m�Ob�N�Y�^4�%Fs�l��v�h�-!���L1�p�7������<�@�Fj�U�Ɯn�;.AR����k;�x��C�yA���_z7�CJô������"�S��:���:��qej��)?���u]n�Q.Z�\;lS�v�ꕬDKfة����>>��41to�Ɲy8���G+`hG媭�]�ʏ3�{����lX-y�S��|�J�L�Ҥ������kl=�1t�F���;&c3�t�\���s�eʂSFm|m��FC`O���|�Z��F�4������,��ZoP�P��f��;6�cu5���JL�ЎO�:��9 ��$B��!��h���t7�I�m�M�1�]�Zw�wsj~��8�"�*�	ĵ}@��7���->Y�\YQ�(�Þ�v;�r�µ�kN�R%���%g��e����K�t9�!��Z�����v�ɑ�n�j�TL{o�9�kzm�1b�/�rԽxy.�:���݂$a4�Wu_0���f�r��6�h٧���׌ s�[7e+n���;�����=��}���_E�������j�&���f��9��ZE�Ϛ
�MT5_j���J�^�j��*wZ�FY1N��}9KP�MF�e���^eT��R�Q���0Ɵ.���7N<����S���F�9W�z�Nv��ϰ)�FƧ�5UW�X��(�P��<N'�t�A�LwL��QMw;��c��5I<U
�����#�Re���׹0t��,���·i]��v�ǳ%�Ջc�+��9
�z�����e��v��6]-�lGD��m�b��'%U��ꅶ��QI���"�P�u����\/ZE՘�yR^>�Sm{6x5���f�Ʌ�EԼv������C��C�*V�����B���m����Y���g�#SO��Y�,p�6\��>��o�����&=�H� n�E����
"���EXE�j��r-��U�'�>������O�O/sߵ{8�J��BV���f�L���l�ޗ�`O�b�tkbG(:�H�ܘ��L�U����c�&
dq-�w*����T��P%�_0�*I~H��LU�$��ۃ�����^�h�
ť�k���!�I�/��a]�vM.�X�R������4�#2������/*J�����t�  ���L�\��6'D���ȸ�Xʾ�]ֳ�t��7�8�d��X��q��`��Ѿ;�tþS��S;��wW���d�d9RY1��������=?D`'V�B:7�J�O��l_=G@v�i�f�����W:���ŧ���z��i��
��t#�f"���ZU�q�(m�W֩�\6�ޭ�Q�U4͐ۖ��љ��/1���R2-���B2��U��@��r 逑6jF���kqa�s�D�xtUb�(=������N�涇�N�L��3e��0_�'|%��h�wV�:@��3W�o�Q�7(~�yfW��y�s؀|�� ���-�3�I��*���Y�wh*�WJN_�@�Rd��=8B�㼮lG� ]��U��!��:fǔZ6��LjZ�A�����>{G����s�_��h�.�2.2
}��qm@^��w?�V���]�F[����
�}*�21Xk���9����te]ҽ�iK�k��-�W=�p$���-�<7��I}��Z����SY��g��E�B��E�Jұ�g�h���'V�b^�3ܯJ�1Ť��Wѹ4���^jZ��_]g���=�u��37?|Ta�apм̳��ߝzb�3;�Ҭ��a�t����+����n� ��V����H^�y�J6��d�(�n<�YZ	V�`ie�Sg5�R}��`K�:J�H\b�"͚ޘ1iR8y���a���Z��:HipG��w.)�7#�\����[\l�񯪠�;r���3�o�/��-�5�ZkY7D<�L���)��~°g=�\��re�D�����^TU�̜�\� �H��Z��hkj�p>ހN���˦_'mE2��J}��\;�W	v�8�Ų棪8h���ވb64쪀���K� �;����g����0�5Y��i��U߮/q뢳_������Za+"��舳�$�����.�T��fEbC����E<I<z��C����$g���ϓ�"~�^+�EXHY0ь;@��L�C=Mע�l���@×,φ������a�K	�6��Az#��%\PznV��A�(`�V�L��k��Df[ql���N��<�L���DwQoP���2��<�<Ҫ~uTl�/՜�;޾qJvu�g��r��͎���4."��}q,��g�\��q�c�߼g��O��<r%W�����V)ֽ��'٪ 83�����:�ENM�(��M؋;j5��3����Ϸ�4tZ����1P�r��[K}Uf�&��V.��� г�EK�hW�W/W�B��ʀ�톾?Ez��x|�g	�K3q�����Rʝ���&:����9Z.fQ@��������l�ވ�@x붎Ԭ��q�e&n���M7��o	�s��mrb�c��]k��}bS\�OH8�r��*�+��-�[�b��vf}�+ʚ��_���p?��p9O���dk�0�l���DI��F���&�7�޴��c�M��Eĥ��ͯz�j�k�P�
�P�$NSڸAH��'f�dI���k�?	��L1�w��gSZ�xaM*���o���,K1^r�ߨU��@��u�U%g`x9+u�k�QB��Z�m��l[H�p=ׇ@+w&�[z�W�R����]`b�om�,Y �Z�u)Q7U�X�v�C���:2D�B�x諫�)ˮU���S������^��#��v�?8u��O�wVC�Q��c���F�^-��E��R7)��c�9�k<�9&�3�4�4?Y�y`�U:�|��NGc�1Mr���x�Kƅ	�H���z�g��"�&�����0�/3�|��S�{W5a�W->cNW9x��\��l
�*>�Xw��l��>��X+,r��k|��/��C�C��On��]��w>�� ~ m�u��&�eH��ó��	��+���S���D��v~�ƺ���A3��4���-�싎�2J9ޕ?!粃��a��8�R�T��GLo�;���kw��n���0�U���j��",�ERX5m��r��7��w�+k<���bW`��ڂ�N�;$�h�e5uvQ�{������#k��Q�Q�>����j�o}8��]��3��}�Cσ}�z^y�P��֟�궱��Yc�t�W�`�Y/Pzec�ͩꙥ,�l�n�=" a��!@9��GVr�TԈ��5��y�B,���o��ǚ.2�uFc/V3�2#+�����w��ggs!��"ae�
���Y6��xI������+�}�{!�@�:����y#CESI��P0D�2!��A7�2%��NKf��Q�ըw���E��7�7/,A��7�PU���L
�s悡�UP܊����m�k-OӾK�g�R~�e��sQe߅��`z�M��F(s�k�am��@Ժ|�1�����;\�K*w�OK�2-��E�j<n�{5��9�����-�&��4m�3zs[ʷ7;�c��O�|�}��I;�	\n��W�
�}�)�W�AO e��'�N�a�1^�|k����ի,�y��65�s-���k�S�����.��z����S��S����R�?9����Hu��3|�]��S�q1�)��M����{���J��E��O�������hv�%����pon�ۢ�m��_���sWnIS�� ��m4;dZ3cc퓬�s�
�����Wj$ \��S�;��G,X�J��N��D���t���-wc�St�}��X�j���N���a �N)ҥ��MPǺ�m��m�e�nBW^��]E2<�O�͚%I�����a/�$������sڨ_U���}��m���x(D�~�k��G���K?bw��/��W�=,��t�3{θ�t@EE�I�s�*��X��*�LtWV�u껆{�z��`�rBP��_LR���i�go]I���|�+�{�N_.�""Bu&��Wt-���`bJVF�GT��Pa���m��5�=
������A�Ӄ�w&�=�j3�ka�A���&^�$���ǅZ�w�������q��<&�S��_��w��w��5N�~�S�4d++��B8�b,�9T�z�R��D�k	؝W.��יӓ�!��c��ak�+�S�#%	U<��n<
j�t�H���R9޸��(�.��iY欕L���uYÜ�si�{c��m��3�2�36\�_<9��MW[���{�c��3V
i������j�����'<��/n�Z[`�rS�(�-�1�-N�~}��|��?|Y;�TU=,�&u��Dŷ'����y�R�����(�d��\F�vƔc{��ߦh�Q�
���P����A&V�eL��Mm��P���t��Wapb�����������a�L�yHËF��w�v�J͕v�S�ww]���-�]��K���2�m�[]�-�Jh�*)���tv��3w�;SP��'��s�cNE�{��s�w�?Vٱ�K��M����Cμ��S�S��^�Ʊ�$���w	�/f\Nd��vpz���0��u���f�)��uiA������)��@�oo/n9�EĠ���i2�̵l��>A�9��o�e
���A�ʅ?mB/h�rWy|bh��b��r��d^��x��ԁ�~�=�xM�D�e�cR~�YB��U���[P�E�;j\ed�c�w0^GF��F+oVcF1냉��f��ZŮ:M�be�J�+ˎj�|�fP���yl�mצ�*Y�I"�3É�>9��/|�=C��`��_�/�R��0��O˟�^J��e-�v���ר��X�{{�9����
"����P�������zmq�Z��:xxq��td�\/�5�/U8{XQ�'��B�r�%8�ԏ�E����A��֧V3���n�#'v������L�q"���9,�9�a+a�G����g�u�/�~�9��<5���M(銻;�m��uV�/��6-*T8�%j~Y�y�^���&;a�rA������V��y�3����������\ƹ:�����D�8甃Ow���Oc�<�,���W,�r+G_lH_R��>|5�*ǣX���eR�T&�i�g��;��	��g:�]�Զ0zҒ���#�iPs�����xz��zKzf��:B�X��N���z���{�`���"����u�>��M��qX�I|����L�k`��]�MpT�����{78�ru@\�)=i]�L~r��N���S���e׽ZnTWq������m�{<��سr����A׎A)��&| N����VD�㳶���n�n3"��7ǻӱ�E�΁d�ͪ�C���u�%b��#�o�D˛�+髞k؎*2�4�s2����[�ȏ��N�w�?.��0�8|`xXmՐk�)�0�=���`�A"K	�@.#��W;�/Q��ݚ��I��z�v���=��®p��X�6�}>{��0���k��g���1�{��/D^vm�TV���j�f�X�ꎟ}|ĳp�o�_m=�r��B�#wy���.73ۯ��^<d�S�>�GS=�0
�2�X�)��J�O��SL��V7��0Rml疋U3�2��:]�¬�^=u�yZ]���%G�Wҹ�ujG>{ Ў�,(�L���-�w<ϑ8��y*|��-`8����i�z`W���V`�J7S���~����&GoǍM������=:���krcZ��f�ɼnĺ���^z�֊o����jmN��]!��͎�']�a�W�S�C��4��m4���|�+{qy�{�̊���u5S��<����Q�$�4��NV���
�RYj�t���ud%�Y�7���1�:���O���
���SMҮN>���d��x�s�p�~�,�:}��Q�W>�5۷�c�p�Y�܆�S�j�DSX|�4�x+_�ĨC�8���"̅ʷ��l��Ձ�Xݮ1Hڷq%���H���R#7�k^	�r{a9��k_N��Z�Ub��W���o�s�^�v��ω©x�$DF�ٹ��nxѡ������ᵧ�A�(-���]�tu�В��:K�v�a��� �r�`0l� ��R�S4%I³6h��s�m���.K�ឫ�)��6��������}��C����D0��)��>U(�Uj����]O5��>E��܌Y���ėĔ����t��55�&��Z�>�� “q�����y�f*�A�<�L�e�ɥ�{I�G�."�UϨ`�sMWG��d��u�l�Ahk�l����?ȉ훈�Z_(�vl�h;G�8�vp[gĴ�>qM}5P��R��Z\�v�P��6?7 ��B�y��n��/ˍĐ��4�⤆�P����u�q�@� @�< ��1���R":�.����D_���oO���V��R�u&	1dX�z��X�M�k5�c嚣�Ѫ��p��L��K�֠kNs�M��oۚ��ZM���"�z���z��%�w\y7�h�Z���:b�Hvn-�k���J���a%�K�vu�7-���U����	÷��̶�wA;	���D'M�I��k&,��b�"�o\3�����k�!wA��֜<�_.���3�:.�3�h)��Z��4����Pa�Lڥ�4���@h�s�^�\�hL�=�9�
Ϥ�bՂnm
�z�2m�;ͭTf�a�G�z�U�����f^���Um���������5����]C��l1[A�(4;.�e9����u���]d�.�4)4�[yS;Z�*�I���vJM�ܗ,��'��6����RK�Z��'��K9��(�9ř8-�qG�-GxE��c��n�8��N�ޮ��PNbd���s3+e陴v�B��+7��e.��=%-���^�!���5L�aoD���^ �Û�noVlI�ŨF�����y;[��oc���A�o`�4v�"��X$Nq��w5N�8��J�'J�4(��I��~����MNM��K�ʾ���z#�O��W:.��5V�m���a>3ɭFj�[�Xq���6;�n���|�����yT�:�`C^V�Z'� ��4�iR�Θ+8���;�D�
c�N9l�]��pgZ���`b{kr3&'��w\D�{���@�f��+s.w��7+'���SI���_V,���4�sއc�t�2�1����a�w�F��JھcyF�_s���=����p]��z�m�J۰^g##.5��fIN�@�oH��޵�omC���f�
in�8��,Sډf�{����|m�Y�\���۶��tj6�rC�g(7B�V]�Y�R���t�!�0��n[i����cʑ���,���� ��kW"�-|YǛsN공2X���>�w����r��&��qe^����چr�����ӷ��g
�ȡy.�w��(�W�qkX�i���,�9O�4��'fҽډGi^((.��V5�}P��'D�X���gc���#xJ�V�ZyGlm��Y��N;B2�f�V�gsy�.���v��=\�f���L��+�yV�ok�Q�'��ۡMX2��n��S�[�1�[��Y���a�dFf
g�j3]���ʉ��Em�NR5sv�_b'Q��v+�8z*&��WL�F;��	e
MG\�L1�t�:;ՉM���{���C6���JI�P��!o�(v�B#Ueb�3�L�����wi��t�*
�`�JOy-��Jvj�R[�.�J:`��n����ԩݎ�=�0]�f���@�����F�^�nP���JK�\دkF^�T�ƣ�C���TP�M�����(h���
x:�� Ĕ��WKO%M%=��\��I@hQJ�@�7$�BD�̦��NJj������it��@
9�J)���!�=�A�҆�D���h{�$h(J䆖�����(�P�(@��H�#@SB���PP�$JR!�̭<�)t��@R�(t�BP�S�e�!�$5�y ���rh
�CIK�Х#����9.��:��������@��PX��S^�"o�f+hXXc9�AFT�O;�uӋ|�/� �{��\�C6�P��F9vrv��� k��k���|x��8=�ճl;vR�����3'�5��=)�Űz�.�6 N�0�gE�D�ӽ�����H���L�`��̼�y�c����y}����Nt��mX���1n�����z�~��"��T�`A'��V1��� �3����wb�޺������o��^��ׯq�NS����b�M����Ng�E�D}(���`�3���p�n(� so�F�3��t�w�\��B�\XxS���������z�cj���KWʪc�{�(���th���/�/Hq�g��2���\�1��E�v��H"���|)H%ϭ-�ϲB7
�ё��;����҄�Ŕ��^=z\�����0��_������Gٝe6A[-uW���ƛ����hr[`��wh���}� t����[��H�R=�E���y���//,]7[g����t���p.��يJ��IK��H�q��T�|�)V��N�$��Ӧ�PM��9�U��%I��)�r��>��f����?���ٹ�L�GAk�<}xd:��j���R��ǯ	/j%3��a[Adз����dX�HLU�2����
��'L6F.�\gjL��[�8v5�=�������lख़�[	�ܺ�s5q�^���o�y���|;��s[���Ӄp�#�>��c��T�ŧ�41�i�ޕ5�@%�ׇ"�H��;��X���g���=�~�N�	�u\}}7��O.�����\	�a�͗�D�ҦRk���qxy���Kd�q?���ڽ�d.<��U�������7�%��BOo-�Q��������VS��qb�R�:E=.�|�7��O�j���?�L�l^��3��t���غ��;�a �]Gb�l~��^w�
���N���#�/t�P���J�B��܆��/�nb�~�c+8:]Ӧܥ��Ba�,�@�ob�'�IA���.��T��f�`x&e��'[0�p����y�l7\۫0�t=Z�O��D�u�Q��*������7q�iM !�e��^<�5��
�R��֯��c�SkY0�s�(��x���R����]��^a[�v�ț�z}�k�s/��3~�x͚��W�O�8��<hF����	>ߒ�"o���|T���<&"�9hǴO��m�d���$(�Wr$C�V�J�^���p1���|���/� K��K��V��'�AY&"��>ق��E_f_�$�J4T�)�ޘ��4�����L�z�m�hT���������M
�uk�EJ}�5����!*f��^Y� ��:���9g	�\�>
h+��Xx�]7��z�]Vs1CwcF1��	c+�$�ݥ�WN�流�̒MY�wϥ��>\k�Z3�`9�1�Z�舲�/U�\���j~��*	Kᣪ^L	"T�cJ�l�g{f�0Gju�v�{�l����4�S�ȫT�,�}*���O!�kzB�:U�{�f�.�QN���UY�0�ڮae-�<�y�Ĩ�7��PL \a�ѐg���σV���/�u��Zs~��8Ъ�����8�q�����B��3���A�Ӈ����z�n�k�0p*�&��LƗ7�e>��-��qXҌ�����u�ݍp7S.P���}_D�ވpbSh�y?(&�)!�"��Mz�5���8���J�`�5�����tj��{�bOT��" ��`�"qPO�Dd_!��-a�xG��9���v��o�]"�ڻך���*�މ�xrL7TΩ�	�q%b�d o�D�s|�M�4TQ���D��G"s�z#����V����:9��	0rC�#��> ��4a�م��D��n8���W1�ݱn���⽨
j7�/��:����M�c7j�p���X�7A�\ �k�A=�(� K��SDS���u�JF����L�ҫ��*G >�N��xi�s)��E3�{�w���7����x_eYwtkn�!'a�)˫:V�"˽�|{'��{7���7Nt�!��𩆋�i�J]��4�́N�`���1�K�S�_:;�we�����u�Nؽ�-X�=t#*Y�A��+*�_kꓧ�1�y��T���Z�+�0�a��p7Z���퍇�T�	x����|hA�^�9��W�wl��ҡ��SL���~�yy�S�繚��[� �2��ͭ���}��zV���xJ���܎��M��ad��{En�>�f�n�3,y�8ͷ,ɲ'�{f�'Q�Y��J7_L^��sX��qY�����J+���B���ħ,-*����ۨ,�<����A��^���#�b{�4KC�����};��-'|���0�OjtS�jÈ�����ͥB���%@0�/�6�W�
0U���6��O�='߳��=��ʝ� _�"�⫓�u���w>��TײB�n�G��Ś�s]��!��P��L�I�و7�c�>>�n�ը�(%݊2��w;Go���ϓ�r#�O��';���[��Ѽ�Ʀ`��+7�}��kj���ە�ƍ����{ɧ�1��L����gҎ� ��N�_b0�P3��P�� O^��O���|�T��̱y�cuL� ����ҹd�)�t��V�V�c���A�&%l����^+���^.��"��;�;G@���IVJw��<&�1��h`�Nm]텛�J*i�iq�=�,u������V����CDjķ���#�s��8-�c�d��b���3�K5�3�7	f5o�3��{{�E�T���w����\	�	x\q/�<X�C�����#�lZ�O������#�&F2���ފ44T*���b*��"3��1^��PVڜc�|��~0b�0�(_8�M����g\��$._H-�	i'�M������������א���>ٳ�̞�0}���?ʈ�9y>�ݪ����0�IR�*��`�Ç/}^N<�{N?�[?Q�[0�i^"�W�ǣZ�5o��5do�75� qK�#��c�=VOC*�ȵl���8~�kB�yD��d��H����R�;�v�{���.�WA�"o����V@M�6�U�,�B�$�M`�2m����Y8գ~z�rd�+�V̑}^9���49h5Oi)�v.c+V��_�yC+�ؗk��Mv�jZ��܊9C�ݯ{��,5y��c廧euD{�U�z���S����ܣ��$4�1�$?j�,�+^ҋNN��~�t����?s���N��=,��ɂ����~Z�Y~�&=�H�;��}�B*1='ʹ��<	Lh�r�B��wE�4]��a�{��Y�vÔ���կp�"_*TV[�sk��a倭��}@�GnP��q��f�<=���
@.w��H3rpƄ�v�>�v�t�<�VV���OSE�v%Z��񓜈p����A�l�YV�޺V�y�;@���;� ���Hshl��7м�F�����R�0��M~��jv����7(��a挡��o5OT��܇.Z��#��`s��g��<�d���%�?"y�	c�c�f�����UD���kW�nu���#%��s>���ⴑ̈�c��H����N���5w��Zb���)�j�=�fE �i�fƜ�N�~��Ϣ���e}��[b"ɀr4����o����E�~G���Z��({�cI|�_q�$ŧWH��妄m	U\�TgtB
��[��+ފM�^Y�;�]�x�^���G���G�w�N�M�t�@oN�ʎ�aP�ɕJd�m�{�6p�^L�D����	j�U<�=;����~�ķܢ�!����Z��,ml��<�����_��lӈ�������_�ʛ<Q��9YG�L���͉��$�v��=��{1���(1�N*�Y-��^}>I�����qt
��O�^�ŷn
k
Jsd��ɻ��n~�B��U^�1�I�m�(��NC��	AΌ�먿�*��O���[�bw�׭���+���/�{�Z'G����5`dx�O��֯/�S����Y-��]X��x)d��o%�m���6*�4��_����Q���t(���"J�h�l�v��o`�DP�{(�Wn�M�|퍒�Fs]k.oM-�Z�(xUl�3����� ��&�|��C7͹~���]��
=ҹ�� �}��x�g��XE.T)P�4�X�ޘ�UL�����{jf��<:ʼ_pL��57�;���e��m}6��ڶ���[�/�7:�;=0�f+op�n�tv��g&��+��!���.%�k���-�����*|���`���υ+ǹo��փ�?O�m{����6�Ą�w�9ʵBW��G��	��/�@�{���3��*=c�
غ�ͨ������O�C3�默��M�W�"�h�����yKG�F69`*4��ŸaS�E[Ƶ�{�Jb�T�G�E��-q>�a)W��E�����n*�C�F���v&`�6���y�Y�"��чiO0�~����#@w
��C���!d�e�B�Y�fa�NC�f�C�o�i���<��G��ػU(q� -���s���|+~�-`�硴M��R��M�a��֞����/��
�¸�U3�xTQs�e�J�Tk�+Q�p���]
ӃoE�Զ�i�Ӿ�����U�=wW<��`��
A�dL��C�E���ZOtV!��m��ժ���,��EӆtT#��a ���7�
΋����"��R��R��*8z����+��/�Ơ���zR�J���/\X���f�K�I�b]�s\FS��{6�rCSc��L�'o�i,�o�}.���K����<ٿt�p�Kj��|�g7��s�T�^��E�c~Kc�E��l�k�3iwfנ�3�|�����e�6u�e�R#ԍ�74_ϦC¶�ʐ����q�I�tĕ���<􈟥��	d�}�a	����oWE���qjfA�>�L�w/~Q6������SF�cjT&��^�gb~�w������M�	�.]zm�X���f{���,a�!�{��9K�!���u.*�Ђz;YO:;ܽ�q���Q'����:X$��������uGO��bY�r�o�*�G��=��ޡ\iy^Q�>�E7u��V|��-�F�T���3*�Z��`J�/�5[*8���
3rb^b����{�*������ƫ�WjBT]��Sh�}r8��;*F\�ߝ�X[���İC�c�⪙9`j���n��5W1������j�qg�\�+,�`�v"�5��|�4#{B�w�����rU)���m�I�����{49��G��F����e����#��-�e�MA댢⁊U���͗�mi�p�����(+�g!�V��s�x���y޵�Tr���`�¨��=zL�}�WЍ�S�CnQ�:�ϔL:s���;l�QFw4���s�yP�jLo2�"mp!f�uAi�c*j�sDk#�]Y��/ �{�+�T �3��
��ch#!�Dl�pk2���-]=c���|��wd^������eP���k��e7<���8��8����	u��Gs��i.�N#��?E��3�,���kPv	 ��:���$�g7�2rnuYll�r�CRq���j�	�M�1X����~�d�=�i��ҎWײ	[9 P�4P�}����t���9�W<LWM���O��Oc�%�,��|�64�kP%�]�x��35���C�l"��GU���_An�Ҩ�x�z���!܋j�����>�g�t��5�&��P���@ؖxAaY3��}Yi��Ċ�5Bѵ����=�0�E�4��p#�p@�Si��"�C	�me6�ڽaH�w%N8��9�O?���J��wO�3U�n�r�6�]#���y�q�a7�����ڊ�Vv�kf�BxL�+22"Ly��jmL�Y�����0/2�Z��v�J�޾v����~ܿq"�u(	��R�?
K|�O��$Ћ�OBj=�B�kv��{<�]SnYmi/����cn�u�K4���gIŮ�O�=ʂ$[�DD�T��P��M@�BK�
�S�rb&�lL�X����9�/ُ�l�T�;�ԓX��n$u�UZ�_$s"�ϻ�5���n���
��/�]K�7W��+��!����Ό�@�el�a[���M'��Hَ�(N.�/T*g�P��b�A�]t"�:F���w,�U4����*�N*<�� �M/���ч��������S��籆d�j%�m��ݷg���w�rP���ɂ:GY��U.ޠ+ks�+cj%ݩc�M7�#�ގ�8���7.��j3i�l	m����E�Cϯ!�Ѝ�0r��<�� m�T=Smbc~�����}j��K6б�CH�RXS�$�������T��`NK�#�9�Z����雨w/OgJ�t�e�<c	�Z}>a���f����(������ʚ����u7Vo�>t:*��3�o[�n��lIʆ�tm�C��P�WҸ2<��?Vi�g/]IŃ1f�!u�rXt�_tWMn|}�m�<Q� ���;ʎ�7���g����]y�q���K۫�Kgf�����������^�F%�bt�9�'3�X�N�C"�G$D`0�i	��ψ�IΏW�osv[r;��žB��ȃƅ߸�L7��J�A�O���:s��(���"���CV�6^�۬�V����
�\�.�zO>�ަ��r�s0�e����l-4#jUW=��:{���ñ�YC�q}��%�*d,$M�����K4$.�42=�}��w=�-�C�1��z&K��H ��X8>���9�)B�G�()��A�Y���7O��4�5:Ns�9a�8:CmnV�p���M��3�6DNk��n�y�#-�j4@Ys~���7��y]ӳ���˻曒��K^U��B+�qw���@��4TK[��������Y�p�`�In�ʗ�_&��2P�����b]	��2����ܽ�X]�b�P���|�����W�^]M2�}��5n���=6,]��\y�o��u=��o.m�ǌ�wa��5�uN܅�
�:'Kk[զ�·X�+.�yr��O�;���[�D<��.�if�ͻ&��V��ZD����ێV-LM����#�q `���B�|�gPq�Zuk�D��sFba�<�u
�w�w-�t��y,
�+�j�K�9(i��r5&ʕ�Y�t�L�M<Fʏ�[Yz���v^�"Ӹpf�5�ߴRK��,��)/5�\�z��q#*���9���]�벛�k��l�4�4=GS�Ո�l�ںV��tW:˓]��5%���%aNu�A7��&@����v�	zs�4Eo�U��(u�*�B��뢳kn�Z�15p�8��qzl�W����N����S��Z%��9<1�W��^J��b���4�FnC~��\��X�wh#an��|�1�b����f�Z�y��k��9).Lj�Jr|�V��u��DЦ\�Q[y���v*�2ݳ�����W��C�Ӳr̓H��{���[��7W�P���խ�.Å-M,��ZF6VIE�
;�������x�E�ϗe.fĬY�0J���6֮����J�i�4*��BP�A�:�>6D��\2g�U�������	2Y������LpT����/kpj��4v!m��6�����E1%� v٫`f5�l�c�f�[G�ݾa�Ժf��:���;lA�-Y[�.�f�S=��c��Sܦ�LM�A�k;&�K��>j�@��#۳h�o��x�9�2�뼨a��J�ҙ}�t����q�YAE�I%���s��ݑ�zgvv�&F��q��&��:�\�B[.�эNn�c�(Azx���B�M�33�VG�n�=��im^;�m�\�/V�^ͮ�&)ݨҫE�f�kN��O��;ã&3Fѕ��]��]jd�ё�ܱ�P|鋿��P���)����|��uc��%���R怗׀ad�l��z�Z�(���f"�E�p�-��B����	k��5���H�ԉ�(�Y�-�u}���%��:�m��a��X�f�g���M��R��ơ��61�*��s� L����|Q�E3z]��t�:KL��۱>�n����0�	����+,�+*lg�V��B���c�N2�pc`R�T�9+`ՕM�aƸ��D�;k�S&�69�0�Z�g@�tG�	YJBUvT&�	����moL�[�K�]���������E����z{��7�U���^���%	I�}��IwJ=�ѧ����Ɋ�G �p��q�u�%u_��i�nHk�VUF�VQ0*��Ơ]�� H�� �]=�JP:t�A�Z
iy �$

i(B�@:P)JH����"J����B�F��B�҆�H҆�� �#�d4�КZ����Ph�:T�Z5��C@����4�-- Z���ӤM�ZF���:Q�ҕ��ҚMrCB'!�i��iR�(iн�K�`)Z;T�"�M
V�H��4P�- ���b;; ��;{��!��(�V��Q���z�)PB���W%o"�Gs.��M��n�8��s{�tM5�Vd�RK�tr/
�߈@�G���k#x�Nu�D!�A�?mV��x��E��r�����{w�kv}�k]���l��.���e�)Wq����9�OzQh27�<k�(�U�R�*��F�g�'O碝&�����.���b�R���0�z�T2��Z�(#�^��d7ꂧ��|����
qt
��nJ{z�����sPݵ��j�q�hom^���q`�-��\�7A��% >�%F�+\����	�s���z+�{&�I�}�HK���j��υ����k��@�*����[o�'+]Yi�ʉF�+���J:��lfu��g}A`�a���d�)�2�[�C�lj�0����QI�Ȭ��5��L�ۃ/�xu�;���`�Y΅���X>�A�'����/g���9������܁'�[�_G�򦗻9�^���cQ��|�?c��<#��U)���G��	�߳<���V��f5iu�����2�8�l�9c=����WڴߑJϡ2�T�}����0��k���A���go��,�0Vei���1��b�o�ܼB��%ʄL�#�2�r��愭����_.=�oIU.Zin"u�.��̢BW�n��چ|ʴ.[U�6'_����+���SD�{�Β̵�5�.f�&�=����\��۠��BYkl�cH����Q[1w5��n���������[�zH���!0��7΋�׻?Ñ����m~Yo}���ۿ&6cױ佤�&����y֑ϣ��ui��XdV�lR|������=���33��$yY�E7�S��sNtT{��Ь�C�����~��N�+T�j"��s�m�_�5���@pH%pY�~��uTS)�E�I�C8�/��úζ2Ɖ���ۻ[
��c����g"���!O�!�?@X}�=4Y�u֕�������"o+5��Z�`7|��Ly`���]&j�,�(�1�"F�R�d5v����%*UW���'wWH[tr�|Uo�~�d�o��tT�N�ĳ��l2#s�1�vc^*\]��7"D^��s(9����#�z����-Ls,�\�s���h�U�h����[��%��¸[w�ߵ���Ȳwt��73cZ��uK;J_Ҙ��Y,���p�YGOOG�;�ʥ�rr�u��Zp~��#�T2�W��Ԡ�2�{��:�A�b0�9��^���Y��	;t��1��Z�*�vTC�K�3553q�m���S=��˚�j�t����*����R'�ۤb$-����u����3� (zP��ߤ��Ñ�̛ߟ�`𤧊ɶVy� ��s�M��<��,��$�4�ح�.��l�΅f�R�����|�(�"��MpM��C��� �V�N��(�+�k�;w6xۓ]��1z=ݿa�oo�b�ے��j�z�|�ڟ���T�e]Z���\�7�t��9t�ו��jk�s�ZG��2��m����Ց_s�\����0%f3�.�i-�~�r������x>mU�-v�c��}�A�G*E���Jr�ҩM݁x���zc������\cwl��_�Yp�>	�ܔtԱr��f={Ƃ��|�}�N���k��ӕ�9x����%՝���f4{.�\q	�*>s�����Y�E�oH�%�E{��On���k6�w{��j��J�ǪU1T>Z�Y\���`�Wj@J�"b!��
����[E�J�5��	�Oh}����@�B&q��B�ҵ�]��@f������!��jg~�'�����s�CVK�J��\�a}K��b��񙳣x�Q�=?D1�ސ�'��%u�AF�.q8�oi�W��m1�CN�E�g݌��MzI�gr��Έ@j����X��Ҏ}��_�(��U���]��{���&F2�̓:]�#"��i�@�xv:ڿB��\]B�	c��NX��}(�j�;YB�뤷*�Q��sg�&��\/�f
��66�|��Z^�Æ'&]�`��h;i��ꛩ�|̔�.�qy�4�R=�-Z���q	�a���ief�A���B��ܐZ�'u��&�O��|#�O�s�?Zt���Y���v��Ҹ�������,Ԯ��篔������PO�5Qj�JXd�܂���L�/�o'+�ӗ�X׼e�W��I��e��9	�퓋+Um�_X>|�g7�G��T�	_]R��Q�P?�/�m���w�X��LRj� ca6�gz��{p�3�p{֘�Wݶ�:ϔI:�d�n���EȢ����6-�l��5��F��􋡻�OV�Y�>����٬�%�J�>��y�H���V�����w}�n��%�U$]�ϫ�CZ��pފi�ƥ���C�|������QZg�f�u*��C}��L4o��褼j{e6�G��<�����Tu�%��T=�i��������õ]dq`7sr��}鰄Y�2c�%���}��n�\}�󍱼m"��s��_C�ح�J������O�������6�(�C�����>�x2:�A/�̀�]D�]��ET�kʌ.P	�ܺ.:5��H�適(��#�2G|wU�a��^�������<I]p�Mፙ���G^�2T��T3���Ɩp��1�ʗQ|�ț6��`���U�P�h�a�;�W��(��g��c����u�ë���`4��-ͧ>J�l^�ü���7f��)\���<�?/?a���>��z8Y��?��m�޴�_��҇�H��g���˔�^�����1�BƊux��q+�"��y��>�f�ެ]���/bt�T����rȾ�J�N�}H�sW���?������rMM&�Bw�V�z�k��/㱥M�\��}�MO����bg���C���
ga��z�4\��;�AR��A�"l�k�1m���͟i���4�����۾i�4T�.��^wt��U�Ǣ+�H�#�և)i�����G���j�!3ήI����W���co�P�"TF��݃��/=Qz�ҍ�!�K5�a��T����
5��&-�9�c�7�V&n!���#�/:���_:A�N���\b��R�}�߶>8�D)�}�+EWt����܇��gZ��g�/M@���>��ph{��Ш7�r$�|��RO��>��#�Ͳ��i�Hj��w��#ؽg̪ETFҁ�P��3.���WPc~/)���lr�aMQ�ӫP�5������_��?�E�0䕞_H]�WG4��8v�lK6}���qMi��م��k&vH�_����V��ǚU;vv�ڏ��\���D��n1��=�^[�NS�BXVD����t��_�}��^��8��4p��a�lk벫�v��\��e��Bu�������Vo��f�`�f��+X�]�����Hy-š�����V닿omC	��#��\_�����4��~T��x�5
���7 �^s�m-������T����c赙Clr��z��)���$H��Z�\��������?,&�4c͈���<d��3(���L��(�p�X�=7s5i�*�8k�	���.�N�'��ex����=� �+1���H^���gZ���_�7���B�ƘJVE۴��c��he��6,����E��	x,aƱ/�c�=�h�ƌ8�,ڮae�����$<����t�t���y�띜��gò
$q,�x�LG-1�
��/�غ��*�8��u=,���CwFt���_�h���a���D	����Y�\�h��B��>+H$���3�xTQS��e�d⡕�GsvcWR���{�mzK���އ!G�j�᯵Ř�Y�A]"b;��D�����i�k�Q��'�m��ݾs���,;��+v,�V�i�Q�ltP��::��:�_H��|��ȇ�h?�d��}{������m��PDj�lP+���L���EI��rh�.���@:k}!Pzf2َf_�W���R�k��m_-MP��`S�B�0�tW6�;�t���oj��_-޼���P���i���M��dH2�r��o�Y7]��8��a�7���p-ư�,^���ٗY����^ĶW��5δer���&J�﷧��G��vl��Md��5�\@������.^q��E��>�4a�o�$e<ꅣ�]�ҹr��v4���`W���E�ƷP�ꦆ�/��C�*m� E�tѲe<Zō;Fv���%�&����ԣW4SM+>��S����VU[u�J���aBSF��~�T�eb��]�,Y��8��dU��!^�J̄�|N���'��@*F\׋_Y�hn��v(����ޭ��ٶ^��d�~�4˱M��J���������i=G�ұH�jA��oOOV^���b�s����`bbK
&e7qS,���Sm��X���W�ꢂVO�[�F��S��y;�ʦ��LǠ1�h���>�������ɹm�����щ��*;n�)�m_�g&,�1dd�t�<w=��񐳺_!��iO+/���F�mJs�~!y��F�/5qb\�?F�����k�`���Lhb�oM�/B+�w�[�62��$�#]ٺ�V9�P�L[���$���J�"~�o�d�c�>?���^������ʏ�������m��5��G��c��}|��l�㢔�o���H���~^g�Xs���b�c�s�ɴ��2Zݮ�¦��[�a�ZS�|ތ�\�)�]��vd����SS���Պn�u��^��زQ�C�E�9�1^LI��G�6�r ֿx�6g�َ1�|2X���cT�etm�
vB����R�S*�es�~�J�ۣM�٧ZA�W��<�al�E�Y^�S�3������:zD@�oHOw˫X�.EϮ������+���Z�7�hg�Oʮ��p��W��?�{�|+B8�տ>���sȼ������pɑ�l��
�х�f��~���_"|�����P��V׸������u�W8�ԑ�0��3��x��<I�h��gw����8剣�3�rm�n(�7��Օ߿)���M�����:qA�/|n��ɏ�S7d��U�p&�BH�~�K^�e�#m�����a >�&�j����@�R��_�]������Ի̻y�X��z�8[���aK�T׫��/5�3k�W4o�r���n"+�%mP�v���G���=��qԧ�Ś��s/�ᷩ�Pbŝ�f�,�c~+kZ�T�<5�mKje�d{�S�;��{�����f����q��`q�S��GZ�R�b`c�k|����K���Md_C2(��bS���ڲ�t���L��y4:��*1�WX��Ү�y��(����Ƃ�����7������n��x��Q��9c�]�\ݝWE�nӗ-���]oo9��Che>�IrbQ�����#n�_3�.���c 3�ܛ�x���ez����$e�iV|�_V6��ע�H�}_��O�+aۮ�G���6�bR�n��C)��t����:\�/s�5�`�uCfg�v,jξ�&�ڐ4�,�F�����)��X@���K��$��m��j:66���n���j$�U��{`J7� �S=�φa�O�����Ke�2k�2U�͗諶b7�㺎��_��%#�Py�lmy������)O�C%��Z�������lTn�K����Gue�(�&���=���������ͪ�K�B1|&#�Ϻ�����0�2.��zBֶ���l_I��c}O-=k���_C�-��.�C�*��<�,q�|��W(��g�+�3���g;̠d3�G3�FfE�23�H.k6��)�qv'&�o(����kͱ�v��6d��3��g�0$����R����:헖��3CF��!�[�k	��X�M��T�GCi��x�b��z�6Sm$�M��Ɲ���k�yYhJ )JS�����_�"������"�Z`����_*�k_
/��-.Gt4v�0��v�3��ʜ��v����r��[����(+-���-8��,���U�}]Y-��]W���6f�����ʿ?�W19���62_�D��.F3����2�z�m(�j�1|bw{�goc�	�y��˸��r��$��.��c�ygpNZ����o�6o�1'���pҝO�*]PT�֤���)8I�Ɇ����r')����1*���<c��*����HNT���}�}�-���Ԛ�JB܍��v������$������m�	�.�i!�D����R���NۚO��vq丯l�	U�\�"|/Զd)�`��љ��e�����g�Ɯ�������\���l��������{�]9{��Ckq�9�;�4���E��\���|�H�	�.���<�*���>�V��<�j�f���s��U]S�E!�)U3VQz���WrK��sh�{���}*��ѻLF�`�f�a+��C-��>􈄍I��j���K5��@�(@@`��Q��X���|��6�+rd�#�\��Hy�����o;�_��8����g;	}
�,��oRy�&l����r�\se����.+z�=�&���Ҟyt�� �����	�ò;�y;�����
�����
fёA�w��n�WW+a�6��*�M4q,۽Y�C�q.�R�
Lհ��oY��U�/2� ř|�m�4�� D�ķ0n�>4\�q��[�5�J�$�n�m}����W>Tᗜ8еE�XbTmCD�ovTx��j���:y��Z̭��g3:ɠn��������c�����*�g+�p�t�en�PfCX1���w)05滎�(��8˟��p*�ݹ�S��V.ͫEN��nvM��(2ݻ0Q,k@i�Ð�9Zn��x\���;I+�P�{.����WN��ޮ�X����3/>���cG*m<YӶ��Ls �����V"����R6nf��
�D5Ih�됼�˻oih�=����]�����,��&��'�j\�@3.�����1,�:.��KK����C�ro:�Kn�=kl_ic+ա�C��J�!t���pd�ǻ��hB�,d�j��ܥ%����P��[�4>�uٔ���*Nںl5X� �	��%� �vf�&�r�Ag`�Y�s��"X�bww����`���F�a��.���_n����h')�v0gEx�.WZky.���"��QS͜1���J�����|#y����̂���_T��S)��vL�7��y�c��>S���8A�)�+��z��*A�űV��Uܮ�j�J�$��)���b�R�quX���fh0Ǥ8����o���S�!P���ʏ\��κGRv�i<��)K{L��:S�uG�J��0�fMNWi@.�;{F�J�+mQ��Î�β��;�u��Z�8P�%8(��� �G��rw�7�D�)��28�,w��Q\%u;4�gN�fŤťr��f4Z�=��S��ep�)�L�v���:t;B
.�{�u�����"G��֦k��,^`8�����(�1�ov;L-�6�A<W4��e)������d��ʳ5�L{f%��^��o.�Y��;�m�gV�Zi-|\�)vJ��m�l}z��F
oSՙ�f�ý�6Aۻ����=�Y�|%��iWW�P��7�#LhCoY4e�>��u���"R5��w����q���(%���}VY�.k����V�b���9�k@YG������	�k�mE�[W �[IjBn���=�|��]�A��E�k)nΎH��(+�v�/ݜ����q��r/w��IN��d]b��.�3(}u�#%�6���*g\��.3��n��u�!WF����t/5��*jOkk`U�n����y��Ȼå�֔�5�e�g\el�I����j�WҤsV��J�f䁤�6�5�Q���o�+�D��;3���uj
�.��u=X&թ}�d��#8��8���߼xo�
�@�@R����(B��:��GII�t kES�P9 P�K�(R�ҺJ�)B4�P:%.�EPP�IAG�O.�T��R!�ց)�M"Wy�r)H�@�K��C�MiZ�;H��(��C͔)i�Ҝ�A�Z9��JW�rP�9���%#j��NHR�A��G@��$(E ��J�C��W�i҇�aR��M
R���q/y��ЩZ�������v޽z����Ayi�̝u���m,�;I1,Ζ�i�"�#.ww8�z`V����bb�jU�:��rU#�+ob/���w������1���ojn�����v�<��zDF�^*sI����bv����ݛ�ڽ�Z�Z��sy\�,0���ؔ��I.&S�it�'p�����rF�e�v�D�_ݓ^�E�����d8���I������f�Kw�KkԪ�Ӟ��>��n�:�(��R� ��RCaq�-8��9�^w�K��\��O7ŕ�OM�~☦�|5��4�+G(L�nqʌ=�*oz=*;��ʋ��sڏ�{���/��=
Au�;uwK���۔O6���ب>=n���u�ر� +�-��A5"��V9F�<g4��:��u�=��6��З��ڍFj�����o���T�﩮�*�E=�M��ti��ו�֊�$�
�Rv���fV+wʶ[-w7���S����yq:��^j�w���,�����~\.5�걊�A��^Jo"�)ր�'~x��f��7U�]yyTq*f��̥�Zj�g�J͍�:��t�	�u*������}Z:Xp�B8� ���Jx�d'�W�Yy���ll��opHU�櫙�:�>�d`$��.)'>���w��ř�2��8����]V����*���������[�k��<�q���7^w��1�7�
�t�<�7Y4���0Q�c�$n�x�ݝ~�� ���g�y������oYG�h\h��(���fP�[7nt��TqM.~&���P����3FS�Upc�Ɍ���v�ͳ����n�h��5�v�����]�Ζw݄�z �酝1:��}���.��_��v]�2��Ⱦ�0��V���r��,jl����l
���w�_����|�y�yC�
���G1U.8��=p6���gg�S���;�|;I����D���i��>kސ m��_�um�=��9�A��&��#�N�Ǭ�!�FHӂv����,����͛�f�n�XX�Bq��2C�F9S��f���_}�B|��ZZ�~�p���f4{��n&ʢ,k�`��LWf�����2�b�3���HȗS�ؤ<d5�ǐ�Jbl�3�t-��rݨy��ŏ����@�΋s[��o��o{X��F����I���dl��Q9�Ϥĭ��Cnn�]WYVL=���׼.RȒ��]��s�2��hrIĻ�kx+��,@u!��{b�@EL�X�(��J�s��ʘ�*M4����WN�'��ս^�0߽�tg�$m��|�ݑ�W�ؤ������?��Y Y�瘷�N~����S�6�0M�������r��}���O?�N??B^��5�W����W�p�mS����J�c�We�Q�+R�����]�Â�BTx�Tڑ�w~�z�Xf����6U��M'�"֑��'/a-�,�5�*�c���b���/�����w�7�7��,�M5��"�V�8���������+��C˚���3ޟy��kd�1>;���a�k�!l��=��49�}�l�L/l��WG=Q��͋Q��m.�E'�msJ���fl�#KX7�.M�3$�����@����f>�މ�x�uگ�ۓ�u-�l�Zf�/�׵����t:���;���qEժ_�땉.�m�,jl�n0�m��n=�O��_�>k*c��F#��Mo"����U�֋���#�+y��u�̝���F�Ί:&ݶ�-����C)�t�>�o:)B�]��5Ʀ]έ��{�9��Q췚	-e�:������{�gB�(w O<sp�Q9�fP���z�IW���Ul+��G��s}�ы���yt�mO��t��1��[j�κ5�i]t��^L�{�xgo��-l��E�F�ga�Bn�:|�j뎬;�V6)�ه2y��}���EE�?E��n#���Ko0�o��p�.�n��~�9����W�S-�E�bt���>5��":�uH[��XB�m,�����z/n/.-��f��i�ܯ�!���[�y<�agCi��Yz���oDR�ꊼiw]�M�$"s���^NPSt�ع��[�}�\
�S����a�X�Q�VZϚ�ϣ0ȉ�Uz�+�=/6�Y</4��]�ڊ�{�����Do`�Ήv~��.�oM�W^����ŉi�H���M�L�S���bz�we��]��5?Z��:9�s��~��o����]gR��z��a�&��Y����b�i)]VV^�.g�m��#����m�}6Y���ny���c��ׄ����k��^�	r�x�f��r���c-&k�+y�."o��7�T��c����w���8�m�����^��%���e8��r�k�q�z~SK��R/<�${Γ�����Z�5'EF�ln��T�^��G�CڰmC٪��SV�m���ܔ�t)N��I�L��=Z�����SΫ�C~�z�ܴԂͰ��������Z~����8���\~<�V�N�+z�ͯh��%��Wi��k��6r��}ޭ;:C�=Qú�X�,��|�i#`'�����GkO.��2,����i��'���u�tq��`#�@����tO<�����ԠF�!�q�U�\r���|��-l�0/�؃��!f��X��n���m\�;[j;�#z�x���c��ڲ�V��ۧ��6$� 3N>�2�"����D�˹���Iggm�H��hΙ��#���Z�lI��܇����D�˹cwO���FI�����|�x崂K܁O4�&�~Cr�mvq�*�1UvccC���VG빁��Y�z�|(?A���;��%*\`'�>�=��ޫ�k��ލQ~�&�S���h���`μ�S��2�d�X�6�.��g�^�t���?�~�ߡ�3�QkE�6n�s�we�ռz }'M�'˫���Ɋ�^�Ǥ ����w�Jk9L�Re��nq]�A˓;����L�Sw���(i��H^Μɧ˾
�_Sukv[��!5K7u��HK9�e=��4���o����.pd\�/���>Zo/�]J�P�^�ۑP[��w�<M�;�.�/E|B.}�nѽO������1U>r_�/��k	Yx�V�UJ̾��U����rhjƙ-��'���=�:��o���H�}�d߸�n�@��Jjԝ�6��Y�C������w���b��-���g��˿QJ�ۡ�gvg��t%Ԕ�ا4x�ڠ���~Y���I|�3tݢ��-�xX����.]Cq\y�>������*[֕k�]�@���#s��>��'UԀ�q�I�c���/8�O��<��m��6�����/���A%�B0�ݷ!����ħ���_���4�5=�|�5��ڰ�Y���]ϯ0�{�p��±��<��m��ȇ�"!oz�q��B�;�4��#�W�;���<�u��.�,jl��StH���;�^�ؘ�x/�����X��"�T�G�oz�,�s^ͧ�Q�8�=}��b=i9�m��H�銢�ˀx��6(� >�>q�Whk*^c��y��؝7�fb�V�6^���<���1C���+�@�ܚ������c�yOgA]2���)�L��K��+xН�Wb��r}�$�Ș�m��'���J��%�9���>�Geɡ���o��������`�X����[\{q�sޙ�����5�1�0o���uE��t��h����[�D=�lY�{����6�4��,�[�)�_���ӯ!���?O�ɍ�Xf+
��}ٌ�P��{혽e�:��m�5���>>�>�� ەڠ|�'���!�d�F�g����T�n��u:�ɉ�H:D^i
�S��L���Τ\���	�=�3[���&�ӽ�������_N*I�^8���o�%3km֭�x-f��;��@�"�s�vU�5]K���ʚ=��}|�UjVג��fP��\���S69��|=�fOD�-K��uǃ���f;��8hÝ��}�y�K�ۣiveW��|��3!��k�AM���j�ܑ�tv`T��[}�b���ƻ{����	��;�ty�>M��'C|'�>�VP�CT�fޥ���G�;��T�'m��`��0�J�Y]�f�F�|��L=+����G|�|_��s���Q�o� �7Wj՜��b���l���|��}��V+�FS�=�c�����h��.�}*�b��]z��h��:��a�|���sM�M����^bk9��lͽM�'�*�OKr�=��]x�& �fC>nAn�?��V�t-�ݦ{g�n�sl*��O�Ը�/K�6��#z�]����Ĩ�p�}vX���d��!�k��߻�y�Nh���yҶ�����M^˗O��(j�7�c���+Vo\�}�k����n�"���^���J�ۜ��SY.��҆O�ۏ��"I��|���~9Do4 ���hd�~��=k%�$��N���ݛw�f�jGx���:Ҡ�{ڠ8�����g���:�Y��P�XV�-��-�W�	z��P���F�ِ^C���S$�|���[�%S1;9�;v[�gY�W�Ί�݀1t�VA��]��5]6�a"�q�V�tS�J}eV��f�Eo� ���g�	*��4��&��=7���r�2m��Gt�Z鉾��M�/\�>�H�T�1S���ݗdY�ӫ���(�fmq�����q�Z��^B��-�u]*��џm;���M�|�宙@=�=��ObU�7/z)���;R��[�m8�a�2��/R�ǘ�M�����;�Y�"*�9R��1�X��a��S�M�,
��:������[��$��P�vC3��^K�pR�j�z�]]^�Id�r�w�������fnN����̣�nz�=��n3�-���=ZV�|�!�W�$�q�������ySu����$^"��J������U�.2x^2�wcM�H��-&M��nU���v�u��/�<�@qH��f��mO�,�~̫I�;&��v��g|���l"(n͑[e7%�1�U���ĺ%��w|��9s�g;��6n�;��t�i�J|M.V^J�ݱ4-E�9��}�!����fs ﾪ_i
���p�d��hdt�MT�y�t�M�,eT����&��R;�b�k���R��xn�f�`��C阂�	=�j���>��������B�Wvw�Uۻ�`��� >�l�@e�1�Nٚg��^-M�ۛ�^��Jݲ�T�[O#�2w�A�i���l��U*֥*�r�	q;��z@��=[�/�E��liv�g���yP�}���m'�����s)QK��gs��ك ��2�p6�K๸��aQ���h7yb�[i��z�֌��9�WR��A�%�.�٣w0����Eɗ���%�󫬌Ͼ�.��?V9L|9�=ȃ&|9�?O����bΓ9O���y�
��%O
k���k���]�g���c���ޑK9�̴�uP1i�1ӯ`1 �E�X3��H�)��bV��c�Ǯ�9���6�ݥ�uh��z����|��L�0���fgO���9����]Q��5�'�'�/�qi��
���I�&�~Qp[5>�[�7T��I��x��ճ]�Ϊ��gl�_���K+lv\ϖ[<l�����S�����E5��ާ�-�m�����Y@�c­u����K߶� U�)�1��QX�����te�e���$YR�׆�q&#�������U����u@=��/�oLl�VE��w��تΦ���A�n��Ի��-F��J�y3v�������/z�;<1v��<�g���6����Ś7�1�� 0��4��sx���k��!wg�O��[�2g�T��j0���VJ1N!���{�)ٰ3�
a���z�c4�fbJ��n�W�h��W��8��Un���)'�'���}�n8Yn�ږ���L1Ce:	L�`[H-<�tҞo\� ��Ҙ}�'��z��S]-�ݜ�uf��g`hg_���9D�AuNN>Y�;2;��79�:�{��EO;:Q���,]�<�w��Sj�J��m	\2biU���wZ�rZ�Z�4|ؾξ�Cz���Enn�x�Za洆ޅ���nS0�S�ys��~�y��d����'��Օ}�]�v	t��ۃh���b���s���C�H��Zt��j���b�]-���(�)rg
�v)!��YZ�e�.;���-�W�-t^�\�P]�^@�Ṉ��G��Y���Y�d%:])�ig�S�Cl(��̧�ݳ(�l�s���V���!���·������y����t����/U����z��ɼ���jKc���F�������N�[�T�Y��ntN]�vF����	q6�+gt>֔``+���u�F5w�Ĝ��_Gf��_R����Q.��nf����y�`앙�AH.�nn`��S�ͺ��	 �;-r��Y�|u n�#]4֬�O��DI2D�sg_fh�]���kv��<���k^e���g��8;y�Z͍�S�tх�;����gjpm����k�N���:苻�]���e�_*J��c*�u�֞p�@�3Zr�`X�Z��4�N�WB�^P0@!}E|C��d�xe����&��b�u5�?���m�'D
fV*ms��fJ}�5u���r����^ܸ��.6F��7t�3Bܹoe
@1)ѣA؆��@B��"b�;�4
��KTNT�5���U��V�Zr���v������y>�c_��8�����Ł��8&���r�r��,ar���9w�5q���Md��1��e��P>����[y�:Umv�v���q�բ� �;���%l���%�EL��ެF�#��gw1�j)���y���(�-���B�%Y�{h��^���
�(x���Z2��ܾ<� �^˾�б���w-��Qyu�WN8/v<�,.{5>@�r*(�l�`�Mu��������H�ѻ`N�b,��}rL�´�v.Ɓ��-�Y�щ��P�Y`q.�Ztf7����9T�z ���X�Ly0��9����9+.�H��y�3._�o�)^�|�Y�,5�p!��δ�3�v��e�ۈ�k�%vE\�o$�R���]u@r�S�f��n�v]h��w�em�*�P�D��	ȳM|�b-�Ύ�v�����i8��ocs����.��m����ו����Q��ޖC�)�����,8q��7]�`U}�4��\ܓ)�<(,YD2<�@��%{�|Д�(y�!H�
@������
Q�
�i|@��l/$(R��V���J��)����hG�4���J.�D�	@�x�@<����d5B�#�E rP��n��i{@h�#�C��4�I���P�q4h	�t�4���"�h
S@��)Eiy<����J)i���A��hy(h9&���$(t��)�*���Bb���
X�э�KJѡ�IH��#AA�5�t� �G~��������֤o�X�`�ǔ���������YW�mL}u(fՋcm�;���c:�XB��	㻙�Owky ��4s0P�o X�7�_qh�_��iJ�D"a�7V�=��[ G鼒m��Of����11�t�oj�zrt�9�
��<�7D��0�M�[3�:�$DM^����q������9|Kɵ�h�����F��c�ej��G���@>[Ȯ�}��ص����6�sz�qŔkܛO\cs�S�VC\�l�>6���w�}�C��)���df�[7ṟǶځ�j�j��-ã^jei�2�R@����!�2#p��l3�a�8�7k���=�m��ʊ7�a���R��oM|��;錾t,\�EGhfؕ
h�&4�ݪ��89�49�fz%9�6ʱ�W�ǵ5�+F�gDvo7��x�]C7���k<������}h�:W�m��7=[9p��6겞N���V����W^�ժ�(2��+IJb��mԭ�y�5:�k��6�/�G���`K��?x�Z����>L�珫�E%�{�z���J�L���D��h��97BVv���U/&:v���ν��]ʌQ�gnP�5��
�oH��R�|�n�}�2�%P��8om��Δ��&i�����������iͩ���r訫��c�d�~C��d%r\N��Px}����؞��$�w��t����d.Qwky����j#���ǲ�N�'��.��[D�QQq�2�O�{L��B��΂�v�#����~w��m$P����}7���f�A�[\�"Aݩl�)���� ��!�l�!c����`}�Be�u�EPO#����R*#�5�
]�ͯ2i{ҍp8~u���LH�>�0)s4�3�0�.�G��9q�T�����*�I�˥} R�ڶ}�}����Ԫ�	�2����X������l��a��ThK[i�݃��pއHȝz�5Cy��䊷�N��H�����A�q���ni֫k��*�}~��c��Y���O#�	�H�v�M��N�ounr�9ψSҕ��!h��u� ��'b'j`�?�^�|Ex��h��o�k��@��j�ơ'�o*N�Ǜb��zL^=�&����{׻NVu']l^�ȫ.��"=�z���JC;:m��9+Z��s�{a�p���kis�8XuݺũT3%5�xN�٦�m��GSEǴ4�N�p9�pI'�d��ϟ�G�^pA�w�>�q��Q��wl��'�����@��˂��8��ڼ�ͣ}�s'�/b�te��u����`��U
�6��>�D(j=s���RoqϚ��.Ԉ�Ӄ#.�G�x�Q)3B�T6b�f�M�]*��jI9��{���@)�e�a�G�Ҙ��W�ޮP�<���w���޺�*�A��̳�kl��x:m����!� 1U>{5":`eMmxpԣgU���v�'�/��}!�ח?h�S��9ϞY[(��c����)�8�hBݟV�3�e�8�����#�e�R]V�*�$wT�u"�Hk�K.L3u��˅txNu��V�e��Wn�s��[d���*���9V�����0m��d@}�V���V��=T�vE��{ɫܑ�0��]+v����R9�v@c#��<������s�������[�Q��Uśw� �EXO+x�fۧ������h띧'<O��'	ܚ`�9~ٽ����͒u����@�f-SOշg6ۦu����A�a@��qC��7y)�7��0�w��_C�u���ڜ��٭�YG�c,��D+���b=�Uf���d����!�������l����H�[�n�Q���Q��t��`��ij�3�А�{���y��P�%v ���\��r&Y�͹V���Ƽ޾ު��8Iy7��ُ��s�Gl��#�C��U���/�x�3KE�׋ Dd�¯��(�k�#۳s��C��8Y���aL�5>��Z�׻wSX��9x:vd@7�r`>���������y����[E��[fyۺ��h�M��PnP�S�̈�}>ձ��=���=�xU�m��t�8�H}kk� ����z�'�Xg�e=��x����~�����m��;����W�_Q��:���m�P����mG�|=�Ӛ64�s�)�ZH:^^0���>+"Fo!z?����H-�`C��<��b���'�b���Ys�o8��|�:����jW9CV4�o=SNd}�UM�3�߿
7�`.���RIb0�2�����P$��̭���
.���9ҥ����D�Y"dv<��74��ԫ��b�*t~b����x:&�h��״bα�Nkr�	�;Zk'T
�E�陵0.Y9F�Q�����eޛ�ut�[P:r�u_T��	ޗ��6M��<���SD��=��	��]�n�wB�%4��x����2ջ��;�wb��]s�c�6�g��������Zz���#�eJҋ�g���%��f���m�1L�iq�y{�蜂�S�l��FN7����g٧�n�ُ*˽U1ugǫdW^wUE�Sl�@9M�,���怒���8�Y�!���%gi�gZ��1Է�vρK:�"�[�d3�>[|5k�`��jx�u�6����}}���y�P	��7e�%c���nǙl��}�N:9`���x�W^�y�S+zf�s���{�˰�d�E�x�595�3���ΣϷY���n�oϼ��;�:��,��5��M1�3�zFBy<P�9\�}OZ6ǢZ�׌���$��":��R�Ӳ�VXz��<r�;��b�	���i����L�ΰ˽���s�8�n�դ	L��)�]<)7�g!�2r:Ѩ��ל�렑����b̆���G�H�8��r���hb�Kn�3_5Ea���U�_[��m�(.6I�-圮v��j��e9����o�\Ɔ}x&%�R)�R���r�]��V�n"���zU��������o���#s�Rg�C���gO�c�g��9|���A�
��3w�4�O����r=@qk�)/.���@x�|����8DE�˧��	��'.O��^ե�&$n��y�+J��T�xb�0��z�����:�k�M{�_�>-�����h�����P�*:B�uF��쬎��p�͎�ܼ�+�N܅H���K$�u�n%y|�+P�泺 ='i�l����VvO~����w���*��A�3-k�<�en˲L5z��>�/ǻh8`�:����_)��Y�Ecճ�<���s>�����Y�\)mR�+�.�7�?K:7�H�Y��v��\��2��wL<I�KX�Æ���&Þ��x8����ܗг5,�]x�Hz;Cwc(��S��'U�[A��;:v�H�ϣ�:��f�m��ޅǁt��u��r}z�^���L-�����Q>;��ooЬ��#�:oL�T�%����-l��s�ڈ VLZ\턐�+:+�Ap��#�7u���n����}��n�wW_|ơ�&D�n�'%L��_'�D���}HY��R�J��ʻ�-�Tk,Mċ�o��;���8|kو��s��}-�x�����T��d��hEq�q�+R��&�3�I+[:��;N�D�s&!+�;S�}�Z�$!���6���r�M�tU��E`��V��
ͥ���x���;�] Vq֦��p��,s�{B6�\2Β���"��w����{��7���'Vu�-/�
zBT�F���i愯GO�>V,��ns����8�a��͑��wi��2^C���d4\e@�|�L�h���7#4�J(GWLQB�-�[��-@̈́L��t�?L]F_�U�C�WL�^��Y�7��#mLM�.콍�GP)E�SI�|�L�g�^�]�v��W��#�����u��jȪ�^-���k�;���&���}�s�G?e�P��NPӎ�	����>s��S\: NMm�"�*q�JoL�r����Q��^��&��ڕ��å�M*�@�5 (��/Rt#���D�jk�vi��5x�)��
�ze����	W���&u���UG�~ւ��T�ɨ�s�����_��u����A�e ��MkwQ���W�P՗���a,�����%��3zZ{��v#�3v}� s����F2��/�`w|�b����Ww�v��]�wv�vEC`2����8D�L{6�Nlnz鈿>aVn:���]zJD߆*��܁����F5�,f��Q�n���z65���x���g���UW�����R7�-�o�<�q7�ȫ��GUāu0
�O{��j����%D�*�T��f��8y���uZϦt�a�#��i�v�ܩw��"��{qy_| ]�̀ɿ�_`8]R��!+���<�}kv�W#��v$��R\�(���bY�&6G��^����p�ê��)ct�wmX	i��m�C#�~��~[Z����5����"�b6<������(��!=ї��	����݆��O���,��@l� @�3yI>^�n��;Mu�@�2�i�m��$]5���ټ���l2h*|�fF	o2�Cd^��{��1��)D^5��ر�r�_���ᨴ�-�k1v�ywbaI�]n
ۜW>���7��N�(i}X V�2�!P�
�����(Wn�؆%���ͺ|���2,O:��ДĤҙ�(8W7 ׹����HP��n��(r���������qP�a�رa���p�-������|����}f�a� 1/��YSl���D[��k�������V��I�ݐ5��i�N���T/��_{⧯���W����5��{;��r�u�{͌��zR03�<�}aD�?*5U{P󨘼ͥOs�\!�]���1\�?%z�:p�@9L���C���h}������'ZSs�o���ˮ*.��[D��R��M���(�ݞ𽷡~m�'��|�#W�j�o��l�J.���q.�yG��5��:pc�k���T�z�V�l��3>f�-S���*�uK�#�nNH=�������pn�ܔ�J�S��Us�ٓF��j�d�V��/�c�A������[2y��ٯ4���Nu%̆��g�0��vU;GiT�n^0^��Cy���#���nq�.�O�����khv�o��r�ڙ�n��B|����x��u�8y&�,��g3)���*�]2��wZM�klp��õ_�ϋƩ�y���z�bG���n��.��;�7̧j���@��hW)ʻ0PI���U���/I����u���VX�e,}��zʸ���,5�zc��~t���F{B��DX�u1��.�O=xqNO�'�Y��W�18��)G�K��^#�zs'�ڛ%� �a����J�v��Pη@4�'O7lD��a����ͻ똚�֖7�n�Zg���6́r�>��n�I�]O�gt��~�g�E0��~��P��	�ǽ�X]�#p��Ґ���dS�s`�솰_v�87R�p1�i	O��F�=�GCa�dt}5ʩ�[Yך��B��C�or1�h��ڱ�|�N�[� n���S��nB���w��M���]�1�=���":��ׅ��ɉ��J#4�y�۔�f�p��"(UU���{\�«Z�S���ZT�8��	!����W�O�w�F�mIE�{��ʐ/�Um;�5�~����U�\@�cTT8���=+7o��1QrIʡ�� ��!���j�L�Qt����  ��4%ڰOU��4�=�M�\Lmn�/	q=��p��>8��]ڊ�����[.ȾX���뤈�A0��R���f�k�}�������Vܻl,3X�[�t�]�is����[Wt�����؅_^A���x4�tF��c��Ӝ�&����L�&�v���w\Ʃ�m����l�slN��A�*�\�����$K�·E�VJ��=��jV���z�j�Y�z��#�]����;[�_:��� =���50��l�lY#�\d�t�!�L�,�^�X��I��r�0��ŽY�9d[���s�ӭ> ��e�:��Ru�e�YD���{/+2a�k�q.��s���+5i�����@��7��[Y��0E��@)�WH���U:��b�%����4R��3K�"�s[s3(sK����`yFqqak��S���N����b�=�"+���巤D�'��E J��wMv2�[�����_1[R���Ǚt%�JNɗ7��J�W�|�Ǧ���B��R�����;fX�ءÙ��U�D��`�!�;�����*}����;���S���JT�����C&�u�+#1;]9tI��'8���	Ȧ�4�L�gd=u�$�o];�z��h1[��Mu"�q�ruG5����e���m2)!�ұ(�]/�W[{�)p(��L걧�ͤFpE��[K%��4��ΪC1L������XJwjkk��o9H1C���ơZ�k�kFJrV�lO��tvc��B<L�ū���K�z�n�K~TP:��3���\;�)���Zv�f���d�l��k�j��j��n;ޕ��Z���(s�s$|�t����\�7��X�Z�ӵ7�ں�P��Nu��@&����s�M]\X�Ne%B8��Xsz��Dk�����}�&�wi	E��b���fQ1M�K����n���$���P�O3"*pcܬ:�:�4�ij�)儩��1uj���]�)#��ǖ��ܺx�p|��,�*�b.���Di�G�W\�C�ʞ��dCN��ڽ�X��3/-��.�����63�12M�:��J�{���6)m�a����;X���e��.5ٷ��N�xf��S��[y �/��d	1f��H�/>�{�\�N�o�֞�x�+�8��F��2�&4��2�����qM9{�� |�]ʱ�nU'�"f�ݵ���_Hq�ܳmN62���Jy��29a�E:b��,wd�4)��b-�WV��Q�I�NRV̖�^�5��=2���3&�J̆��D�vu����z�imo�,�3z>�qm��j�[]�)zƑ��1�����n�&���3���77}I�*$I���n>َ�L�l9���箺��c�i�^f��Kh�К��O�z��.ĝ����U�1Mj� �`_p�UȎgtT����*M��WW&�;7c�{�k��;irG�I��Ǵ=��T�T[#T�������4tKHS�4TCm�� �)��h:�G-#JU��KHm�iZ��S�b(&
�A��(i�JhF���h��I@W#@D�U����(���h*�"(t8����%�J)���yM!2�h45E�IM�!������"Ř=�$E
S0�4Dǌ��<l!ESKA�l��"i(*'lU��b�*�h�KZeu�(�h�R��Z������"�����**)"]&dP P�|*�mU��4��偭oosW(�5�U��s�4����8��t�ԃ�cE�����Z{:���x�߱1�&���������k��;<A}%��K������*����V�mØ�Ms4"�l˜�}渼OZ�A���:�H�&Ax]�RޯY��v��+|;�������F�D�ܺ�1�����V���X���*��V�W�����]:��߈���Y���*�	��K���䩾���[�и�.�V����YCo$#�wں:r�����..����dC�>�حJ�݄�F����9�K������0s����G[/ی���l��� �S�W�\PoZ�ވ3A�ɬ:*6^�`��ݫWw:�+ݺ�Iֶ���X��+�½<�Q-(���;��xS���Or�ϳx�_��Zr8B����{V8��o2<�Yێ�S~��n�5�rK��5kM{W@c����GvsGyfR���(>���^V����/����<A�q��
F@�=���i؀�����(vٿby>��r}[�J�TLU����l�2��~�]���'׆�q�m��/;�)�tqdЬ�ּ�Wg ��Z�W�{��L�Kם\��]����;��Pm�N�SN��o�vu���y��3f�-���ܼ�߿��y&��'�����ސ��i�Cx��|�f��7�t��X�c���4(�f;kj��`>���ɦ�Sjg��Y��UxD�U��޿r�}��'v��f�>U�
�U�r��ђ������Y�� 1U!���N,"+|����SToA�=���.����{#���8��[��:[E_��r��`Ԕ�acM�}q�şe��4��c�w[����*�J�o$%wUfrn۫4�S(�Ɖ��(�3�4���et���^Tc�l�v�-�dR�xkT��U�}�5OVp�l��=��q��Sf@t[��!�[ŤwbD2;�d�=ٻj"Kvu���۽�Ԩ�^����,�`qY1�t�OD�@���y��]�h��z�H����yݡ����y�s��$�c�ˎ����9��bޥ+/;2gMx���Ç�/W>�:�-��Y��	��k�C-TY����k�����9{Ccߖd��B:�:�:�*���P�d��x*�r�x�ix����w�]"��Cǳ}�W�jv�O�6���R�]8kHٜo[�;L#�U���k���	��}\5����y�E�g,�uը������:U/��אּ��)Ӗ��?l�U\�y�,n�wVXKJ��#y�k��@�C��w�w�}�;�����~��|���8���Ԅ�Fo+���k V��5���{t�i5c1�g�~��,w8�Y��i�ꋃ�wr�cr,E����ڍ�?;V4T0�|���K�v&<�e³B�oV�wa��N��S����果j�7\�Wxh�9������|��ȼB�",�������6���2�f�6!�Q����o]�&�H�N����|��B*b�~W\V�ۉ��������w�dϒ �6��Hf��i� �N��e��x���n�f�G�jF3N��v��]�n}j�+�iS"�y%-��sU��gW�ݗ�C������[bNn6��M�r���wJ��0A8���[��i���C63�=\�w[�P톪�2��<�&�JÛ�]��F�'קn�L�� ��G=tjL.ʒ�cahӵ�r��ƭ>9�iy�uF�n������8"�[X���Y}[��V1�UuZ7ti$��m�茾SoEfԴ�*[U�5�-�c*m�pMw[u��8b��)�/�Jϱ뼨���n.�;��d͗��'mx�)J���K���T���m
R�������O��Y��e�F��y��YT����W��q#�Ԇ{���?������D�Z�;�x���7�݃Sޯ�OZ��iJ�@�\��F�/.��2nў��w��e[��Jw7���|�	�?e�+��2^�R�j��F�d�����Y�|ۻ C�ޡ1�+Tȭ\�eAo3�ӛ�1u	��Jڝ��نp�y��pǣ�x�F����޻����f�,����y���Fgg�??�����O�!�!����f�h}ӷ���b޵�X�,k�����{g����6�k����ً}"��Y��G��}������[�۰}Ǜ�N^�	�>�=����K��ʮ�uq{_�q�|'U�B��s�ã�8�f��1����+iYF仪�Cd?�1�_���[��AR��fCf.�����G�һ���#K,����vel�c&�Ҡ}z�hN��2��8����C'�a��n�%j�˓��3���w"S�!E̻�XRw��Co�*4�>[t�S`��L��g�utWշ�5hm�Ĺϱ���_`	X���;��LH�-p��O��n��Y�32�9fo;Mw=s�#W�ȉ�wS�f&�ׯs�n%F��;g�!�u�J(�����wUe�6�}��륝_�R��K不{�}�LM��eY�3�v��4a�]�X��em��J]�L������t4�s��|���Ѷ�2�s��_.����,�ڲ�k�fUx�x���Q>�%��e����ɣz�9���j'�xG-#�@Y��v��+Ȑwk��i��b�%��s������	�� {���Fc{�o��j^g�w��t^�-#p�Th�յó3\c-rb!|�x=�Ƹ�`V�07���{���9���O��K����4�w%/5���6���j_�P�U"����1�{�ӹ�֦fs4��������f��Y#��Lf��Ѹ�b&"��7����^1 Y��,�8#
�j� ��r��r��\�`%�k�P���y42b����Co��-b����O9��t> ��ds�^,ө*U��¯7T�H���\��;9��ǅ�4�1��<����/��<��ͪq뷪sխm�8���h�x9�Q/WH�?j�rU��s���[l�����b�ZZn���ڨ��jsPͮ�?-=���ygXZ_]G%,{ý������qc�7�x�6�9ˁ3gM�wi��d�5���2!ν��W��Z���@�Q�~:���x��G��k�ו7��3v�2��r��Z&1�p��(�jm�5��V^/��������2f/`iv�s[&�<uHӯ��Qt+u�vЎ�c#Sj����`/6��|=V����yJ-\�(�ұDVh�l�� oV��. Ҥחc�i�t5��@UO�٨y��t"���:3�^��R�w-�(�R9 ����PŐGKh�zum�Tj����d�sB@>KW7,�ݕ�R�-JV�ʪ��Zt:'T²c����nfd3'���Z*9>�['�Ejӏ�d{�e�R&�*��u�����}ݖF��<,T��s�>����t�z����U����t�Wm����4�Δ�sX,�hf�VlӲ���	,=u�n;��/J�mɀ��3:��z.��2���;�q�˵\�'	A�>;�pH�Z�.���wv�7�u��q4��������۝���N�����KC��Dh��4��at̚S8"�`����+I�����ɍ�$��Q9��9�����t�N+�0�
�2�g\�Od�6;+y�yO2���C�`�ܕ��X�nj���?w�����`�g�Ef�rsq� ���YO������ޥ����W�M"zGh�n�޹��h�R�ޓw���m�n����p����XCs�*�h�{o�N�?J�	�B��,֗���t�(�k�R��NK>��׮���u�]�;��[����E�6$�o�\��O{��{��Y���>	���K�+��v�;dvHs"�3��}��Y�b�=z����X�[�ESM]����+״ҏ`��H/!�]��?`E�az+�I5��C����%�����Np�P&Sn�NF� x�HP��M��%u1��g���- ���r�#Χ-OU�q��\�z@���]��82��*`�{R�9��o1F�X���0Zջ����}��p�KD³'�Y��clfkYav톲�n���l��Q�j녌��K�kQ������4&��ִn�=�PA���넌\:�E��\�i+�0�ء͌�����F3�9&�ώh�?M��+��T~���1���[6���9�]�����"wFm�A��\]����oc��,T�[�kT�rJhXdв�JiA��<��CED=sn���[��z}t��� �;N�F�r<�g��d�5%nX�+6�gNDɺG�m-2z��I7i+���U"�If��o���a���}:�K�xv����+J���U������Sl��0�/��՝Bfr�6mcnqm�:@̐�ݝM���x��b�� �{Py���4��i��W�,�^��o��j�ȍ=O��;9z���zٺ�������M�G-���p��:8��b����X�;�1�W��ֻ'��4�u�m��u7��M."�!qg��숲0�c%6�M�x�F���93j�[������Ț�>��+Z�>3q�Z�دW�~ˉS�Þ�W�����U�m��E�*�G)<�kn��7��A�7Mz �Q%uk��vA�s0V�`�x +M�NN9��ҋ��1��/,=�2�μ�ܜk�%��g�%39.W�#��ʝZ���'����&���l?d�hb���a�f���ח�W:{�������n��d��gg��3����[�2����o-mvC-��vk����������Q���3Ͻ!��ꠞ#zG��jE$=Q���e���f���\V[���Ӎ��Ow��	麈�sL[��#���p�՚X`��/<c�L��g��&'ۤ��Df���������oC��.����v$�܁�:�
SQ|�&���Gc���5L^r�1��֣�����
Cz2w<_u�k�R �
�]����j�A��)�эq}�G�/�H��UZ����dϭ[�{S.��pơ�z&1;���%�m
�=�%{�vC�J�]�(�5eV�K2��z�[�S��
��`D�:ب��O=ݹ�(�h�&s�o� ���K����exo,�@�iTlnV�n�`Z��g�[���m�դ�{%���K�OΎ&���S��s��Xy�M����Z���O9�T�<��-d�÷����Рo��[9^���;��%[��`��i��܀�}�����E^�*[��P�7,N�����@�s��@h\%��޷'�LT��#B�¶�X�O��*��ݴ���ުo��^���]��� ��;"�?i�*�&�DpΑ�p*3I����l<륋*ԉ��'���ڴ����e����l,�u��:�:����ԩ_^��g��y�z�:�������cSf�5��f�-�(�|�8*��Cp�n��YS[:4���4[��!sU�tg-jm�`wE�~ϲ�ڲn��b3gV{^����G2㝴�<���L􄭏{U��yEz}�;���ؾv5�X��Y��5��)$�OC7���n~�f�h���ڷ���J���3�����3��_�>�٭���߽�y�����d�Qj�f>Kgoprɽe1�턇oil��Vf&�P��v\�2��F���e	�9{�����wp��� q�e�al2(uq�EV����ߟ��bP� ߭A����e@V���Nc�q;����8;x⪼`    �( ��p;
�� �T �A� ��@ �D � �T �P �E � ��� � � �@ �  �@ � 	 @ 	 v�� $ ! $@!@$ !U`�  �  �  �� ����� *�@��  A  A��8" � � � ��
��2��+���A
� �*�H�B�s�8�++++�A� p!pH0H0i2�!���v�&|_W�T�EH$R(��zM�~�����})����O�|~���߱����N���O���7����뿃���W���eUW��_�?���~��E��Ȃ���K���	�0���ү����R��+�ξ��E;?�7��CȜ
7�?7�����>���븛��'�f�y�X�UV�@! � "Q � 
 �Y � ) � "P � `@� $�@ ` 	 � !@  � ����LH ���ؙ�����E?'��j��� � � � �~���}+�'o��~����S�&��?��$�/�����O΢�o� �w��~O��{����ß��O���|���� TW��)�W�?������=H�����UE���)�2�������`ADW��O�uA 
�����H��n��'���I������@q؃�����Q[�����?�� ��z�0����~_O�O��NzO�?X�	�������@E|z~�����D��@��
4�� �@"Ҋ4"� �� �J Ј4-(@��"4��*#B�(��� �H"� � � �B"�"4�(�H��*4���@�Ъ4!@ % R��" R�4��
�J ��-@�Ђ��R��H �-
P4�-*#@�Ҫ4�@����(�J��H4�R���R"Ѝ��-*�KH%(�H(}xQO��9���J_������%�����O�~3����<�I���� 
��O1Ds������Н����'���>����>P�_���w	8��(���}�����)����/�����)��ز� �8/�9,����������0d���� T��%@
E"�Q@��%T%H��t�T�5PJ�J�+�&��r��BJ���J��R�����)w���x�+��ke*�m����Tِ��[.�E%������+��٪ٜ�ͳ��Ҧ�6�[�sCRV�����mۺ�٢��[���0��%�Rd���q��)wx��j�F��6���]m�%R���uݩ:�J���w���kUMb��[Hͻm��Sa��-��7x{ʪtވú̫X��ݻ��[k[]�"�IAn�-ޮ��u��Vs���ɗC��g .`�$������ P  � 6����R"�m��]��hd m��  ���  :A
U:��h � ��i����\յ���-�:�r�^     T�4mJ�(�A�i��F#F�� �x�%)T=HтbS44442@�	 M	��i�j<��dl)�"������       �&MLL`��jy *P�44�@�@h�  �xwvxW~w�UM]f�tED���x�AN����\AU{�-\?0�L��y~��?�i����G�"A@(����?*PD�-"�1L�P�(�&�{��v�-i����W�˳z
&�CYf�@�R@����ki���%�n��i((�>����WV��鄂�T&��n伆/rC<
�T�[y��zAM�7i�\
�Ihfk�leLR�N�,�y�ܺ[�p��(*�^��5.�.ۍ-�U�.��J��)Gn�8��X+E��͛��MZ��a^ީw����Y�3%k����,#Y���6e���-TuU�Y���G�������Dmͥ/T��Z7t�`i�1�ݰ���C%��7H�� ل�2&@f�ש���:cA�i��/-�O�P����(` �wz�yLT�#V.��@#�:�+kC�M�8���u��Hn���m)14%�аa+"S".�;ߦ���ݙz�&�������m4����'�4���L�xP��lތ:�bn9���b�
f,��R�Ǵ��#8P��3fS��9X(e!�4�X)cX��;Ū)Y�npӷ*n�����X ¨BʻGn��m���6�÷�-}CN2p9b��W#Qd���;�Re�0ɨ�2ӭ�s"T�� � ��xi������c�ŨɻS�*6�7h6�ɶ&<����fRR��F�⺳jXǣZ��ؒ.�e	L&l�B(U�6��Z�yu�TRJ ���E3J�G��#&��yz�Y��m�שiy��n�^*�o],@T�-�Z�yV�I���r���u".l+�GM,�0���n�ˠv;JL:u׵��p6$Dp�:ӻ�Q\8�|:�"�G�t�y�%��;r�.����EIY�I��T��F$�3���J7Cw{i[ývy�y��:E @ôu�YYCO,:�"�lW7A�؟a���ݥ���̭�)f�Lq��N��m�4$<����5��e%e�z+YDa�xn�;"Z�Y�{A"6�GsB�J2͹dK�ŧ"�5`l�Q���:�ʬǤaf�^�Rm6U��Y�d��]��-A��j�8[�����I� Yd�����˵�=ȣe��k�>���7qХf�S�S]�%�f#�e���jXV���m�¶�Xev��(���W����OE�V��:�,12���!rхљ�漧4
h���A�6l�)��[2���54�o����̴ko��XP��Q�<�[�n����@��V�+VM�B2����_0ܺcc�/)�b�p|��͗v�q� (��]f�^Z-�[�����e�uln���Y0^@�����V���V��7�ܷ���4+(��at�hY�O��+�'�F�yz��o�im�S6�Y��C����/�㩗x��5��[�1�Q�qk��MS �`bRady�j������ò�-B��we���'�eb;����`���"������V�`�`m�@�Ծ%�̛r�a*���#�䱗��C f(~%b�V�:�J�5�S��: �\�X�-�Y�4�J��j�"���_�l2��]��Z�DU��ln:Vn0Iɨ�&�A�.G��ˠF�/.��n�o-Z˷Ya�!%�1��J�M�36�0��S@�_+�inܱ��&�r�ǡ[ʐ�;�����62�����V��2a3Q*��!��bi�w4�y{��.�&86�kfR��B+/#��Y�e]��o2C	;!з��4��bx���)��#�o0P�s.����YeV��L��/7qYO�bM�o ͔�]�;2��b�[4�L
��{1]aca�7����=a�
�x��ai 6��̍I��a�(�a��Xv�%dZaˠ򙗷��Hnn�wU@�L�F�CDX��3h<X�yG.Y�����;Y#�f%ku�#ҭ ��:�Ҏ�l�Ki[g��8��n�W�Tl=u�3�B�Ԗ^	Z6�n�ֆ��;�7��%�N4��z�\�mfݜ�+{f�0~U����hk�n�Ј��m�9B�*�)U���{.��@�`��;�M��嗯.�v������0Jb����;tw$N�nU����A����*�yʅ��W5�#wL)1�;C�f]�Jw��M}g�Y�����[*,�p;_i�5Ooe�,��Xksk�����d�����nŃ��QW����bH]-X�U�SX�͒}S�ش��A9���ٻ�h��׏�j,�$�Z�o7&��fF��(��t��S��",^�x��J�h+ox|���i���H}�j́Kk1�Mz�����{zf�u��c0�e+X��R�V5�sXcd4�:��N�i�u6���SM�ʀ5Nĉ�.�\��Be.�P�:��ѥ[�;�`����ڵRȭfLh�R���R(�ws:)��N�����{���hK#4L����N����B'��,�Y�R���!��d�0X��mkܛ��NV噢����5"Q��IV�yb*�H�;	A�pր���R��*9�.��Z謣kUӴM�]����Ǘ��Ut�� �߅�y�q�$B^��E>�����.�����ۖ���;A��鐺$b��h	�
��[w���qO`��'����1➭p�k��BS}�a��"�;8!0X��p[�eN��J��9R��L�ѝg�Q��WwtNqڹ
�q�L����4�7�Lig�T����Xa�Xbղă��	-T3S�ُ�nԍQ�WɢLw��YZ�)5�\3�fWY�Z5�f�Ѯ�݇Ǧ�oL/K�-�%�{|:E���5�;ZF,�]��(*%;��X���N�L���՛}��P��"!�ws7��B!�1X:R-X��"�p��0�h�p�miR��֬�؝Om�BV�Q�vM����-U��4��d�fo3����h4�:ڦm^�۾�*�m$N�i��+_R6VTe����U����̱�po+�
��U���Gr�m��{܉�X�P2�)oj��`�|E˻���m�Y��|9��Z��J�SH�Q�����K/on�y�c
kJ��l:6�Lf�7/��t���Y;q�K��ْ0pAv�w]� 3�x�%�ܰ��C�*F��FF�fE'K�� }>(�6��$]���D�&h�
V�U��3�;�{z�
:V8�6��M;�ܧ��F�3YjZ;QI�⢷]<u�����-�c\7�:U�ѭ�g؏�v�pW ��F]��zd���[q'vȷJx�uۺ�^�̐DH:�y��6|�͞��ځ�Am\�f�'CB�&�s1ٛSş]�K�e��S�m���k�t��'��i2tb�xd[x�EF/l��!�=M���Ԡ��Y��.��u��Wt�z�:*ێ_V m��3�`9�A2�hca�)rKU��h(�2L`"*ee,FN�٨��H���edͷJ�їZe�T�Tt���k1�x�NH�}	�eښ�fM"�<�I�&�ufwk��m���]^w7vja5��QV�EK�|^����XU��u���nݶ:!>ю-�*���y��^ȁ|j�b���zn��F�������j�]�q��j�*�'���Yt�,iΨn<�6	w�U�Of��os@PU�]D��:F4���}�0e��z�J`��e�N��c�����\uF��Y`��C��2b��MS)���r�5�7��b��U��Z�"ۜ*F{/�ݔ2�c/��X�~#B$���10TNY$��78f�$� ���j��y��s��cn*��1�/�uq��a��K�ښ�GsM�g�s�b�:{r��e;��݁%�v郂�t����-�.��U�����LKoy��+�)�,#�*��@�x4�S��@��<U���n��&�[b@�2�/�ô-���ep��w�������pg���N2j��z��6���7sd�H�cWF���^�!����&V�;D�BήZe��C1+��l�{եv.���L�X���Oy�2�������V���j�{R�/*R�����_Y��uS#瓬ʾ�f��;�`�Q�K%Y�±L"��[�+�(͗qRl;����2Os�t��և�u�:��#��<k���A*�a���e'��p�+^̤��:�l�t�Н .� �¹�ل��;[x�E��c$�;�d�¶����s�,c�[��J�H2뗛K��ׁP!Ԅ�j�.7g"���M�^S�4Ū=t3��<{k���-� �P��ד��X���ژ�z��|�Yۮ�l���R�,�ڼ�P�TY u��t��y�s V]2���n��U��1	Έ>ķn�I�2�/ �3T�I�*�.�:R�U/lZ�?)
vKe5���¼x�bĒh�Y,�������l�����8�ǐZ �Dƪ�j�\/>6[�Q$c�e+��I�x�Ã�q�+��j���F��V�hd�b@�j�6�p��7�v�.����lWNw4R}�\4u�A	X:�mJ��d�J���앁bb��fV:ܣ��Y�d��V��o�i�bGԝ�R���zt��fG�0��'P4=ݠ���p�j��v-�V��hw]�>m�j��LMw�'"�Dd��	�D�PEê~"�ǲ3�����-[}�S���r㔻WH���0*^��p��yX� 5�                       6 h����  5�X�������B�Ux�d�MuW����ёvM��vK�zgU�,�8A��Ҧ�
���J�r���P-�ޕ% if��i�5�AO�|���-e�p��^����p�u��b�S+j��RQv�qAS���
��]�5��=R��m-�S{](r�[*nT�EgtVp�n��-j������,��1�wJa�����ؔ��La�y��W��k��)[b������P�0fy�EU��1��o��ۉ��ӕur�ޯ������kW��DN�j�Sл����"w�$x�����}���'o�7�s��!���#u.�{�#��Bv%��Y��-�"�ƶ��w^:ң���P3v�i��*]��9��`���>��>�,�Ð"(�JB����^KX�vU]��N�.Ȭ�F����,Se��SW���.�4PdRQ�W�*�r��y�|�p��_��:��F�Q,����2��PP��I��ѡ�4��:�q^��\�5�j�o��-���{�a��r��^�#`'�vNnWy��P��X�VM�z2�R��Y�L�7��؂�~�E�� yK��@�Rn5��� {���*ьݧrR[f�hGq
��z���^g�5���ʎ���y�u]LW2����ˆ��ѡ��r����5ev�����]�B�-�ϱ�!�C�v�U�bЂ����*.�b�r�ּ��,�N9K"cN�՜�N�Yƭ��N������=���?�_h��j��VVmK<�b�ӣR�-#t&�lRH�h�[�S���7�*��MCIɨ�Y�s&<�v�Ƹ4AF�[���'�=�v��7y�%t`�p�TKgV�ʾ'Z�����ݐ��5�����И�s7i��d���w����y2͡������.�S��3��K���Fs�a�L�(��=Xl���xb���+0SIJV�:�r�7FD��\ݠ��;כy"g�i�DH7���a*$QۣhSJ���0`*������(�fjCn[�x]��iΤur޻�j#8�]L�<�[��R���NN[��F���֦�:�/��U�}��<މڋ�9�L�q�R�Y�%��R�V�Y��[��5U�:��7�a,t��Y�ce,���!ӻ����kB,�Э�)�U8-� +.r�]5)�ɋS$�yˤ�1m ��w�-vWQ���1Kx�=����������.^��j���`ټ����	�r* ��)��s�:��VSf^����ecQ-��/c� �F�Zή�y���S��ئHk`�IO�]�]�m�`�j�Vɯ�k:O�{� �-]��u.�L5,TХ��MR}f�II�l!�,'��Մ_\��0ңz
��1ْ��n<����u�Q��]��d�����a�;�^��s^@��a�5O��]T9V���x
��������V��k� �5Z�ڗ8((�˦ϩ|U�m�d�{l�Yㆈ�Lx\7Xl��B2�����X�Q[O�栭BD5�m��]��x��Ӡ���R�1|�<s0��K��s�Z�ɻ�Iqg,���GFU���{R����������[�UF��yGc�J�DC����m�ŽbIyM�%�ٖXb�Zv[�v��8'����u��}��^;�ѷW��ٝKۛIlՠ���b3e�]v�h�����F�Mq�"ц�\�,tWvE�"��â8�ӂ�7\�-�y�Q�v��rZ�δ�X2��V�	����.资Ȇ�CK�]B�l��������7U٢��NeR����!vj%�ܪb��:��֌�H�j����u���e�tJ�Ҥ�����;�E@��d�j��k��+�L��W֚j�I{�u��s��C	��1��=CE\�C5VE�01w->!��WoKW����$~n�+w^Ff���\���<��6]EG���!�c82���-�4�n�Im	�\�#�G@�e��`��b`ӌ�t�6> �n�S/7o���� z�(5��ޜ�<4ᱦ�j�&���7CVߵdX6��P
g��V���=����ER��]��H�*��ٹN���Tj9[l��j�_.�8�����HιL?������~﯁Ԯ��&��F���*Ӕ�����n��W0��0|�]�ɭ�R�&%H�7}���y���R<�n���i`q�Q���']yvM"�m�f�����/6�Qb�����P�9E�%6]�uR�1%Y����Le���s��ճ�ڥ^�w��aQ$���z\��mń���
T��`g.a{�n������L��7���x�U�J_^J`�U��+U@�Ҙ_&��OG��}d&��d�m�U/m�i˂S���Ie���z�[g��"VY�T�+\��c�i�x�۱��KH1WB�Z`ۅ��K"+��u{�Kd%�!q�о.�uS��:gn���3��Z��t�p�[��+�-R��p���j��0/������hoh�jH�=�r�y׎�+����9�gNޤ���{�Z'Ht��s�,;�`ه��i�E�X��T�`��M%
�c�Yu���J�NDI.7�mmj�ͱ�m�rY��5���ǽ���m�t�V�3
�2͎9�F�N�V]]���P.��56L]�� a�4�6��>x�� xH�	'�M)!2��ʨ�s�{m~5�G��;9�.1%bX){T�],��S��8S�@���Y�iB��K	y��1����W�%�蓥�,����b��Yah�X��X���w28!j�aV06�a��y��z�ql����*e�M�iQ����O0�XV�39Pͳ�-RE&��y������h���xs�,,;d�   .�FՊ�9���n���E�����}:��b	�̉��!˃�|X ��fLA�]�>$�t�� Y1 D/O���7����%:A*�-���d�$�P*HUS
��,Ir�����J	$�)J$�*�m.��DڪꍣP���%F]�T����Da�L���J.^QDAx��$��@D��&`İ^cQ2�*GWI�2�ʚ*��Q�I�/n���]P�/E
�����7����ouS�]����Wϳ�^Չ��p���0��r/�_o���p��E�n�/z�{�+�}��l/l�׻iP`�W����wg����X&�ΰL4;A�sys6XQ�UY^ah'N���\ ��H��,���g�^��v�ˋ�zm ��5��w��AL�k��r{<U�üƣ�|vmm�a/?I���sǤ��u�]$��rBIDz2|mkg!em�*#��gC�&��j�1�ao��j��@M_Of�ϣ%R�lW�`*�^/ <C{z�XQL���_mw�֗i���K���e��m$|��oʟ��f��r���_޽]蛷�e��e�Df��w�g�W�R��(���g��KG�F��Nyf�s�.r�M���
Ҥ�rQ��9�Qe+� ���]9\L�X�9yy�˨�C�Q�(%/W�����^�z򯴎��oR���]9z��ۍ�K�9yׄ�%o�l3;7��=��$ׅq��|��x�(����?v)���W���G��'jP�2�Xg�7������Go|,��y^M�M�Q�j��ɱ��Z}�Z|���m/镱h�2��*ni��Y��9$f����f���˸.'@�n#�K�G���P�+�I0�ϱ��^�@�Ζr��Z;���:YACM�[��V-�ޏT�1&4��g���I��piYe�K*Þ��R��,SӰ���^j�U���E�F࿥�L�l��y�#�9�E����Q�(x�{\|��^>)�`>u·̑)`�:,��4����
TS����K��Y�5|�,8lWX��Zcǎu�z�g4X�3h��������$���]5�h��,����9����N6�<l=�s�4�<0�o��=�H�7�g�֪I�9.c����}��콪���+�.�S�/��j��O](����/�L��gw��~	�Ѽ�&���� �y�E�B&�sE���H*�	�ʝO����¯�zm$m.�gX�����^��^�q���_�ud4������͂�]z���T�`�s���ɱ�����Z�#���MՋ^����t MD¼���=E����`�9����4�z���=7i�ǘ��sdy���$k;l�$�b=+��	�����
��n��އ2$��%Nu��;���� �㪀b-Q\���g��_��Xc���H��*�ct�čL��b�Ǧ�U��<r'"�����8v�C�+{�Ϗɧ��\ �����ȡϓ�7���3���,�jX���x��
qj�YW<������c�/�-�.�ߺ��f���c��l�fun�2��(b����˛C=z�o2�=/�(݂όHu�-�PT�z�=�6����l��|deOj��ҝ����<택G��DWZY�H�V��]���=�9�HW@�=��l�x�[r����J(�Ɋ+�,���I�d�|��]g��gc�>P��:�\g�M�T���߂�	��	<�
��Ƹ.EO;�W^�;��x<�KxJ�G�i�z�4�<���QO�M��Z��&�������h�x�W���N�i\>��<����Lm�[�f+�mT�(���Z�	�MZ,��9���PS��x�"TGsG-��ʷ f�K���<��q�v\��}R���G�Ъ-�o�y�ڞ&��9�y!��>Ϗ��ٻC(�1����<��z}�$���k�V�Po,E�Y\��58�Z��O�pWw���>J2	ۥ09��s��u����m�7!�U;/�8N�b��r�WL����T,-������yą�����&�9K�Wjj�i��8Kܑ6wx����A#ڿH4n�LW�N��L�g��C�_�%�9�~�{���E�c������TlM��>�Vu�qV�\�z�{{��}z�yeb��2�=���T�ǘL?5dh3�m?rJ�����{�R�z��p2sm�\O�P��=�YY׵��I��Oϑ]��Wf*���ᑀ�` ���3&���ղ.���;������Uj,d��m�r�w\T]���g$]C(����r֪#X9��FQ��n��J�� p��j���W�r��}�K7`Ȱٕp�J�r�w\�6>�[۹
�+�e�1>6-\�ձ@��eK��f�Z]�,�b����ȉb��YT��;�0fTt5VQF;����E4�w$��Z�����a;'%g+��5���գ�Au�RAj�{j�D�u�g$�!�g�8��s��ꇶw�{���E�J2��t64�+�1�^m��嚬e�5��2�KV���JZ����3�R��;�횻�5�
@Ĭȩ�b�����R)�L�͹�_Hl,��*�7����w\�C9V��K4Y��Ad��d��U�*] �׵wc8�ޑ������ub�*��^[m�CJ�2ut��^j9h��������Lt�갺�v�>�Vl����T��3t��O�@��c���*#���Wv҈6�J̭���i4�   eY{���x�-�}��fY��c|�߃Y����'�|�@@�|�$jUSP��FT(.����MF��U$	��S.��$$���uf��ID5!q�!"H��*B�H�UBHK���z��T�	.��\*Q(�T*J^ �H � #^ʝ����x���<C^E���'�vu$�=̛Y���up��i�	��Z�"�+�tg�w^��si,y�|t�{�\�yy�DYVs�VF)O�^�W�jq֥�9��N]R���ӯ1�{އ;��Ƃ�u��
�G�/����{X���C���^�h����{]fx�F{��W�-����fo:ٝ)�3"��ܾ#r GU�8U	��֡,O�pk��o�`��Z��v���u�RW��[���~�i@}z���L�j�Є���E�t߻ma�����`�52xC�|�g���$l�� ۶I�~o�5�SȾ{H�۰4K*�㾝�}�b�D~�ٳy�7�نg�njq�l��L��a?X��ž�2�
��z�\!
��6�Rw�L�l���"+ ����GLs��^xӫە2�7�,5�۲Ҟ� j�o�6�cm�2(�5�����y��g{ȝ�\�/�I���fVR]����J�E����R1W�:�P���>~�\�(1!���z�#�������c�'	��}K�\��E�>O/^�å� +�&/8�m'�/%��=���(�G����h���tɛ�U�k׻�޴�Y�J:^���� �6�]-/��M���kk/�eΩ�z���Q�nH�foZ��\�.#1���B;������A]�N{@U)R����0�j
]��eV��t�����ߩ��m���:�좉���#<l���y8n���Zul�Z�tZ�3�^�.����rK1V�x�5x������3h�g6�Hnn���$j�{�el�w�>xm(!��/s�h��2�a��)t�����נ�PgKm���Y�m�i�E�-h��z����^��g�I=��IPh�2��-���<��Q�r72{qt��τ��8F;B�QSzo�Qzc~V�ԑ�H����d>�6�)�7���v�r�O��2��SYB�p<���x��o�J��7��n��b5#5W3�Z���\�f���im�?`~ZM�2��Î��eҠ���e�0C5m}��T����k/^N�f^�e�Ly�z�I�gڻD�ᴿ���3�~���F7�~A*�Y���E}vF��ɺ�0
�K�7�v�w1h4��m|c���jP͒SY\�^�k�Dz�m}}�����Uhk�p1(��ߕJ��h���Æ�����^���;Uw�'�4Z�+O\�w|i^�{�Ц�ZH�W�����K�3�U{��fdz�R=�kw���t��������=��v=Gʼ&�q������ׁ�[��V��\^�c�������-`-�Y^��hกn�7��Dy�Va����<�Y����D�O}V��#��B�}_+	Ŕ��Grr�I�8r�A�uk��@���P�ƀ�M��	E��v<3!A�s:E�y`�j^�����7^R�]���ġ����}f��k��Z�q`􇥃|�?�W�ğo�xoߟ�d;A��͜H��&wF-�Y�^Q��v�{���y����[6�^1X+6��8���ϩ���#�T"�ZS��=z��erg��T���I�d];y<���V<�=x�``���L��{
�!����#�eNp>U5V��!Tx_�]޵�3��˼3Mn���αc�X��S����?s�qΫ�����\���0O���n���c�����by��h��A��W��ߪ'Bi�0V����W�W��h�c6�����o"{��7]�fq�sO���3�
�o����M���3����=�龋N�c���3j��Ȑ�xż�w<W�e_������ONN�ҩ��K�C0��,��m��,f��kg��{��pYK\s�E+R���<�$my� ���Q��j���ɏ��PHM\^����^�yk�bK���Ult_$7�;Z�M:�z��Ԡ<�j��!�b�\���H�P�g@�w�|������졞h�=+�{�G<���y�^�Vx 륑�%�@Ys�Ո��]����3nU���Rl�+M��E��|I
>O��+�x���[���p�7|�	���:��C-�$&4/��c��������[̰ڥWo�
f�c�ł�]v}�o�j����k9�q<�ubޕt�w<F5�u����.��{;s�C�j�S��)I��2�j��q�Je�m�W��3j�ޘ��`�� h��q�����jʟ]�ojQ$:��Za��{z9���Ԡ;I�x�=�����QM.wה-��s���eY�{��Kh���]aݑ[{�����3�"U���э�wUed�ͥ]������`�s�@���Z��f��iv;�)�i�n�*�����dV��]`&���㲥��f�rs�ڤm�$]�m�o>�e6��N���VG�W��-�W�j�	��	m6E�*=��!V/eJS�e�R���Ie�F��D7��-�n�Ø��M���0�7Q��P�˥N�{�֓�^��Gp�Oh��mY�jX����E�՛��%�E�����    
,X9�1�>���`�:\�\?Q���[�'9D�'	F@9�@��5�@��VC!��2H�2\�T
�aUP�5�PrK��* ��@*&A�.����$�L��2�$r.A2F)q2�3!�G� �7 0���=X�94�2��uK�ׯ��� �����w�'�LL��}��&o�3�|Ȭժ���G��(��;���`�O��0�~o�ooN��<��ﷺ�Ĵ����^�8W��r�@�ʼk^��J�4�g�A] +EL�T(���TF��%N��ĳa�{��^W��#OMzQ���Y�F��=�w�~4?nYaݜ��5�(=�;���N;M��zM��J��V����Ϟ��;:��)�yyݖ�F�攮�P�1%�u=��~f!΄ѓ�9^������Bvz�ls�y�!}��{:AJ��u�y�r�2G�~�]�O��ͧu�[�U;�g�wj��ge�X��Zx�
�)^�/F�����^�R��(��|�]k#��f�R���-���^LB�`���s2xsNՍ�&��2+����{��Al��6[C��^F���!�'֮��9�e��� WH�K[~�ɮ5�d�4Mr'��G�C�������vz�pd9��f��A��^:�<�9���6�6=/�"�H���K+��Y�h�%�O�s��q�t�uӓ���t���ȯ`���X�x�����o�/sYp����b�"|#L��A��8D�S�W�_W׮�国ζt@��˭CM�Ume:�Z�:l8�Ѱ�������غ"rJOq3;����}V_��+?H�	����,��s!)�-v�vxԓho�쓞=^*���[���vz�
 S�����������wUԸ��J��},�,q˺�k���縢_���cʭ�E=�����
�V׽u�62�jݾ��KP�{8�7|n�k��W�}�Q�K��;5��LýUu�C�uC;�E��}�Bdm�b�n�����x,�ok���wvȤ��1{��,��ێJ�)<��N��'�U��)W��K��ڟ+w/�JUhr��;�^�V�.O=��pkz�ޏ�?	ē�U�;������vl�PKg�T�yRT&�6�q�YL<|��|Kܬ��=d#(lg��wm��Q=ܤ��_]��i�j�kfSwZ�}���u�˿h^�f�y7=vR�u�ܧ��-FLyXŧ�}���ǌ�8oB��N'�֘;帗x��f��'j��Ą5�|<}<���A�I>���G��]�L���΃��O�y?��f�lz(�j���-Ѯ���-�s¹pfLLM\���{�=�	�wlC/����>�s�Gl���v�|�s����u%�Mrûmg?y{�[͠(���'���^�~�s5��p?{t(��^�Ԫ�3���W��bf�"��u���w=hկ}�2NǓ������jy�R`Kf�o�kE3)(HH�y���"L(/*y�t��zl�:��ۮx��/,�1�sr�� =�2��x;-��U<�n7j�0Ʊ��e��d��/)�{��� �ַ���9`��^
.҉~��dc��rC�Sq����=-#J��I��Y�GNլoԼD�����k�ٞ�q}yn�Tc`�1���!L�h�5�^+tv��7��l\^Wי��Cʉ�kd� +(�II��rQ؎��Z�ʐ��8�Dɯ2���.�y�������K�UsdE=5X��L ��*f��ñ����$L��n�|T��������y뉃J-����W�jW�аEn�f6+4���g�ʕQev��Y+�3�|�8;��{��g1��+6b�+O�F�߼�����þa/a|�/5��rRުWE���ߙ=Dyav��ɴ8���A�dű��XY$ b��S����&4�+M?6wM]�|���w�9�\Tu���b��ʅ^�z�(K��Mt{��7���'#)Z���A�PG̅ǜ�黜 ����aqh��~~�u��ޚj��Ig�
��W��L�s/՜�D�]��A}����VU�@�������Z�
��n%N]ulv_�����qo7@z4Fg�B���>S�0+��N��b1Y�2��˨��z�H#d�z�SW��>�p`�:���g,�ΛV�.3~"�2��!�o����-Cg,L�V��Ej,�~�{��c{��b� �,�,J�j���A>"LaQ��u��2��%v��nL�8��2˩έm[`m��7�u�\�&.��+$m�#�=Y���V��9a�Qۭ���n�;��U��Ǣ"��Y��-豭xVN�Uw��I�;@�+������
�w��hG6�&(ژg[��A���y\,.v`]� J:8�4us^���2����g1�R�S���d���������UI	wAM+E�U��n_$�b��׋��:B�Cs"��Ʋʓ��88�"ge�Z������<T�KˏhmՁA]n	�� ��[W�J�@	�Z%e �-e���`XϢ�]�R5�   E�F�]Vk��ŶE;�g1���,�6G�$y��e!��&Dh�P��*#Q���*T/)2H��J�H� H�*(� � � ��|����G�b1�<�Z��]�YjS�̬*��k����{����5���Xbb��vP�ک�yS���_a���L�#����e�����;;��)�{'�zc�z=*ǡ���'?ߜЭ����e[�Th=����';�lQ�����ٴ�nw�z8���=]^l���>G�[^���k}^��}�D*���ZU9�^łV�Y�X�z;/�{ȑ�k��=@?w藷�7S�)����Qc6���	e�n~���y���f[
����DP�����j�RY��z�AvG��������@N�M���(�a����fn���*_��w���;��eٴKՊ:I�:ZQ��j�� ��k`Hs=����8 ��wyr{��-z3�=\�pp��wAwfcW�NZe��UcV�e���k��j^��1gy��9����ݣQ��1wb�b%�'���6DS��D�&�˼�V�O�'��N�)�V"����e�.�k���<���꜊��{��IV}5lk���~�Z�xo�<Qe-"�$1/l`8�ff�l�{"�%������c�]����5+ȩ�X{���I�:67����gv�ŗ�{ކ���)Mӫ0��W���CS�n�&o���~��<N����k ���Ԩ���(C���*���UU��������X�R w��҆��'�Ē�xG5>���(T�ǵ-5(1�0w�=F���b���ԿW��gvL���_x�E��yT�]��[k^g���%^N�3����S:�GF�z��F��*��v��V7�J��T܉o+\�0։z��'�mTPM1��yVי��	3�S�3/H}m�ׯ�ݔ�f~@(��<�N�vV�֟X�P��������W?y*#Lc���J!%zP�E����9w�w�=ٷ�ț5e��69��Wd���yv�9�n�O��b��:��Y�tf6=sݷu�~B }�-���Cާ�I_��>Э�w�f]k��NA�������	����rR>��|Toȕ���f�'�וﰨ���f�h���en��#&s������^~�G�H��=:E��랰tn{��-o���~@V�佾ݳ=���X�"������L{lל�L�h�}^w��c��v7�%��w��u��}�����"f	�ȫ0V��&2�kW�Ͷ(���x�tݝg�:�o�V
���r�µ����z��W3�~��G~���� �?qm�'V�t4)h�� �0��թ\{"��úob"\���`�?Sfx� a5�+��%�X/̗蔆GS{<�=`����X��凲�45�����i��<��'k��y���
�˩IT˓��K�=�Nz���]ad@
W^�7Պ�T�*�W�M*I�9�����x'ȉ�=��'��2��lHv�̝��Q�\����o�rwL^�&��(+���=�7�{I:G(��jy��+ Q&Ĩ,���N�l1&L�4:N��=��h�cz�X�S�E�u��Q?phf�p�4����1\�����E��{��n^=�������1���ىM���2�5���2�2���"�2r!������r���մ��3�� �A?W搣�?�\nͽ�{}�ϼke��Y���"vIO�#�h��E^ۉN�������ͮ}�z_���ɓ�@H�>7Xj�ѣٗ���|��S}��+c뀦�b��=7Z�'����
�g�>��RkE�j�缩 NVY+�jw{��[�G̩���^�E��ۺ��)�엜�TP���� �H�V��i�̺���.ɳ�zә��}i/d/�>���m{��<b�\'�#������z���u��<y��@�+缼��q�t'�+º���jss-|�5�O���S�[�W��n�xa���J�������[�mK��^L/��{�n�=^#[��W�����Z���4��� /"=���OA-C�Lh7pmsʔzע���n��}7f�d�w��(����0�j��a�ۦ*�nR��j집[�X���Y��v����Q�CהG,jV�\*.jQ���U��r�:8�l�P��퍹�|U���5Ƶ+Տ8R�G\��gd�w�p�)kV���$��^�Rw:��<���P�wJ�c�7�sHm0I�xva�[L;��S��Ӛ��yX��:��z�[T�'�����T쩍�dGqJl�6�-ef�k��Yj�;j�lVh�T�7��eCӯ0<�鵞U�E��k2����yMv�%�pq�t��������{�B����)AHbs��<�ݘ� ���=��;�M��]	G�(���������r�j���&�#6,C.��i�)�J�q|��A�g�j��4 �V֊�(�;�"��	�[�h��Q�z!�'X˥ƍ�[r"��9]d���j��h���Er�
v����u�F�iթ�yJo�%�C�����Qm]*4�5��"ݘP�i��[  �F�f\ֶ]�z��,�/-�#$1�D> #ix�	�cq��,��2
H H7��*�-��%AdFȋ"�PF�Dn)��� ����<wq�lm��Ӊ��م����Q����� _�nW욬߈��bk_��k��My���)D�Ҝ��J(8���W*_�iX��5���D�ZGt>S5Õ3�d)��cJ/-�&�s�扫_����k�^W��a�g��0��4j4}2<�^�\�-QJZۖ��o_e�����n	�}����^���:c�Y�]�J��/z�#���3�y�44�밭S5~�CƟ�A3�Ό��P�7���[��p�e��w�g-\�}t��]lt�2k򵾅I��e8��8������V�:<�h7�t��i���߄�����vX}�Y1��Ί�Dw-����z��O����JU�������C&Wh<��#��<+&ҷ���;.�`4D��U b
�jS�9t�Z�wJz�5���m�;��K͸�#�%���M[]���+��<������`mgA��eC���fzFA����^=��{��I��l�>̕wGV��W{�<��\���s
E�U�<\�B�z.��L�S6��F�5o�p�Z�۹Vr�qA.}<>W�ն�����gQ����-:�0� �A��u�3ub���\�s�o����-R�����w ���KsK�Om8{I�lѷ�V��h!#�'�%c��ZᎽ��AKK�ws�-3����=�~��GTeV�T��c��{�b	^;���z��vY��Ą���H��$��z�c� m>��1�T�G,��n�S˸��:=Q{a9���5�J=<��d`�ꚐwWh#W�p lZ�Z&���sbwٴ��.�um��aKT2~�F�?݀~�n�K�ϑ�w��R���Q
��V�I�{ �kW��aCz���3�^�h���X�:�J)�t+r��E��.G1V�5~UE�МO�KW��	�{r��t�����!����0���ކث^W�-�.�w���
�ح�w�gO^���+P�ې��9�:�q���-
]ja��t�Ӻ${��~��[`^�ҷ@��y6����`&�~�{����2��Y�?QC���˗�Op�����ǝ�(�su���n����}S^	w/����W�{������F,�h��Ω�*x]VOs0��˥g�%_��r���%V�_�2�'=2����y��u�{/Ia	¶UFH�׭n(���-5�7��Ͳ�[���mg.�&�	idV�!��g-t4qO��� ��U��k�� O�jZbx�''n�Wv"���NzR�^�^��Vmy$>^qD��lÞxa�[�ĭ����lB���+ZMd�L�ݚ���k+����oa����G\�N������V�מt�R�p����
sύ�U�$ҧx^f���������bŜw��xT�����ڊL+��m�^����zc�֬s���?W�(Ӈ�2%W���[Ӆ*U+:���2�����:�^�	^~�o�Q����!h�<���
z��v�e�NS�_u�q��3�3Q�D�{�gG�P�I��ĭ�|8�y�uB�o=^���y���6�>^̮����;�Gs�ك��Cd���۴H��'.�]H�I����R������D]����SB߯�>U_.��?����I�w���-1;��X���@Vr��r��4�c��|������[�N:e���hF�fWw
��9�kU�O/�Y�)�{)�����L���<��9S���Gנ���W��Ǔ�=�?:�5�`��}ݵ�!��=���o�M*�'���ԬB�����7�2���E�������%L<M]�{��>����W\K	��E�7�~Vu�M���Tg}�Z�l�J0��>]�[�q׭��5��<�~�>�_b���)d��ʃHd�u�s�:�r�bkʺE����Oۻ��
&�ѽ[�n�uC���Y�6�f�/4Գ�-�/���WBp�ĝqH2���d�mmt�E�DW��B�ɶ���	j�o�9	�Z��[��L<���Rv�GVXSz�f�έ�!P�:�*��P����(n���CL�J4��.pqdo����!�{+%���Y�<!j�g��Oܬ�ӥ�L��ԧtR���j5�M���c���Z�����E��n��c�&�����n�D`��AC�׭zL�,J�l�+�6�X˴���GC��<}�^�orodU�6l�����Y�*������J��.� �4��Ů�rG`�Y�;Si+�1ڳ��0*���v��i]r�l��ܲ�u�B��[C�!إ.��8Q{��^R�EI5[n�sh�޺'sl)�B
a��]%���۰�C�wU��v���Z q$PR��N�/��|����7d����h�Vݰ )c*����S4/+*rȼTN�2�t  �I��3.]���7brM\�e�ɯ��A�����D5����r$�H
\�q$I��H!"\A�d��"D� \J��	�$�@	�Iq�##r��#q�[N;p�����^�]Bd�[�a�����56����/���{4�/r�p���2�Y5�<���~�Nѡ5�\�S����vPg9��Ֆ̂�W�S��'/�Kٔ���lc�g��m�j���yW���bn۾�묡\0ǖ�A�}���ȽO��f����1dM�9&G��N��2r�
�.@�y�;�(u��ƻ��W,��sz�"tGvLsf.�L���Vro�1���7B�����L!V������Jƻ��"�:zb�����~rzM����<�^�t�~��s��ˬ``�F�n:�˭]i�v�,`��^$��Z�U7�����%D^�4�zML>N&��ˁ>YSk �<��#��ae_f�����+�%K̷W6'M��4�=�`1z������n�YBA6�11����w�]�K�ix[w�������V����=��d>�3��cu�vv�I�e���Ʀ�-m.J{����^�D�ѡ¯��3���9)^��l�zϏ���\�Wk�Bx�^f͇�*���.5�������yl���� �c�j�-�`ky�W�q`�q���Q�����TF���G(-y�f�gu
1;�6b]��\vQ�f�]܄�BN�g=�U�"5C�m2l����I�SP-1;R/$���to��K�7�mze'[yD�*�M��<�K�e�^��8�㲱)�G���s��A'n[�m�ugC��`�
�XX0;i15�Sņ��q��v����yz)S�J�����G��5�]lX!z|sl7$���[�.�FwN	4�1�V���ѱ��k(�����
wի���'�UĬ[[6�(Kς�^�E�عm�7��X�����(�^L��:�#>����2T�k;����_� �N=�ˤ��t�t5�L�F���^�1ѥ�v�l`�S�N���0�0�����v�dMD}3���u�� FV{(z���觔��U,��R鳦e<�~i�.�'7tf�JV�
�i�n��T�7M��� [b&7��B-w-�1�xxc�����*�b�G��>`����jaq{�[,��X��O.2��4F�x/=DY���-�{ӷ	�f�M�+7����g5` ���5ﻡ(�;}Rؚ(c�����q�0Y��� ���7�����W�6����T��~�3��ӿl���O���
�dn�4z���^c �=��bv�'"�[6:H���$>��<p�1�	�
t+�X���<����;�kzD���TVY�Fi #�O�v鬮���b�6]*!WG̺��\�O�]����؅#r�$�]�Y�.�������b[�K�z�ܟ�Y��<�>>��LhP�s=�e��5lz�9R��r����O�<Vgp�	����~(u����/��P]*=ɋ0�'�۶����f�8���+�h��~�)&�6�V$\u��A�~��Y��i��gT��������;�;��
�~�[QJ=`�U2��O=�7�/����jo��=��0�g=�*��n�ߤN������k�~�O�e��n4=�aÚÄ�z�1�7\Yb��R�?{A��$������,<��ŀ#!���ɱ�77�迕U��H>�?>������Bn1�~;T�=~�r�vd:,L�p���-d�-��Ƀ�Ϻx������^�#k��RB�N��;���3�&�KI�fUn�i@M"6pmV\@r��5�(~c�z��;���=�`��<��]9���h���룰�$s���������8�	��ep�Ҳ��Y��M�3�zQC��JH�����ig�x'-32�AYz8����U�\��UW�4u�� G5~4��������#�d3%n��5���v��+l������{&ݐ���f6�r�sY�^�$(yV�n�v�$LJ̾L�"�$���zy�u]���&�\�\�j_��ҷ��SvE���;"C��h����-�X��V�K��3~�V�{.�-�y2n(���(e��
�KViĠv�=���`*��l�Of|�p����<�k�1`��_v�6�j�K�>��=ԝ�S�ˌ��]F�����!]�(%Zl!BP�&5olvC�ǗCit��#B����+]d�ӻ�{��1�V�!;�WVp+��*�0ۭ\�ٷ$����z���+��AQ���o�\�!w��� V��N�3�}e. a}�����Z(�%:�����k���F��.�Ҕ���I�}���8�an��]/�Z**WQ��ueX���[vl��_t�J�X'�c)^HL�/+�:m �6�m��6hy\��ܷv��%ك��f;h�	쨸���Z-�2X�1�e偖e֓l\�G�U���⺫�t�W

B��3V���v�8�%gM ԗf�RY�:�ge�/9��v�"v�|Cn�]��ү������,;m�03��9[J��}����w��^𸘼�U�}�e�똷�   �
�Ń[���Uq(d���5�M�>�&��$	$���$$ �TL�7��(��M��5�.$�H�E�R��9�dQȆ�5�TL�TE��!���T)Pu.(drH����PX����Pȕ
�j:�dAͶ��\8p�{��9_<=�mx��ݓS�M��s2R�d�򗔓��3i����w��˙:����g�ky�L��=t��:�����uq�=O
T��R�}/t�>
"%^�Z_OlZ0T.Y�j��-��k�S��ۧ=�t��>��TL�����Xa�u���.�V�q2}�%e��FUe�S����ѻֿ���Ab�����N{lS�m��eo rY�}9�K�
;������ٽ�0^�n�!�C���_��B��u-���%�~O�k��Ir��_�rȖ\������dWV�yӑ��;��&��'�����6�����L�n����Wj�;�|����g������k�q.�rn�������PqR��X�`իY��Q�$�r�C�7mqp�l�R�\�"?��PĽ��{�wߥ��75����`�j)q�ɾވ��d��Nt�L���bM4��^�+/y���ݱ=�-��fMY�I�ҷw������ʄ/e/c�uÊ��7qk[��Dq3!�R�t���N�z2����E���_��q��༎�Y��0�1���2|nl]Uk4>��^9��v���e��b�ӱb㍂Y5��2�F���D�Ew�w��;[\ܯ�\�'�I���rn޹X�����&ߺ(�T�{^ɋ�\��١;nu�b�Q�v=]Zd�6̳�����]s���hcn򭗪�8���@�����}��U���$��N^4K�=^� �}�t��C\V��K�V~���c"n+V��SZ��D�b����apоt3k���ܫ����>�[���X�����}Z4�bϿA�2g3P��?MW��>��Ͻ�s_�Mf�(��:d��4{�o�b�+E��p>�U�\�?�K}� s-��*wS��,�y����C�U�^�������{���<ˊ�\)��{΅����'H�^ӓۆ��(Y����-[��V%���~��m b^�o٤e�FT�U�
:�\r�f���:~���qY�Y~��U'����8��VzTwjA]k�"rF0�5֘�J���(<�i�"`�ȇ��VҀ�Y�K�)�+J��l�َ�@�&
eO���r�&5�y{s�g�>�z(���׻^;g�ܞo�E�w�ꞻl��s;�9K��O���:�b�/��Dn^��O ���Y��j��]��#����O�Y��4٫�����o�]�{۲]���L�]����ru`���Rv+q�:X����IN�d=��⫘��SS�k�: ��W%��G\u*�#&��o7T\k�I�}�3�o5� �������б,��.;:,�I��+���@�Se����W���w�of�r.�0�����W6�X�ZNK��ˈ^�lAf�@u��r)��憨�;ٸ�17w<��랮�O���{i�E���٥�y��<�K��{�<�v�Y�P�8�s��z�ѽ�$�4׸HvwHU��������㚚Ԇ����h<4�����3��M��ڶȣ9�K��uו��*g�\�����֗{��^!��Y��Ҳ�o�D�a&ˬ�����xG�kk@�lul�qd�$��{���l��{̮ ��r6<'�k̙�ڋm.\����/I%�t�D�9�gf�T(U!fO��)0DE�0��or6��Sv���0E�ID0� ���oT�})��5E���ko#Da��3�Ayԑ�Bg��H�Sn`�5.Q��@#������3���ckAw���i�>s ����ʰ���zH����8x�����ܵ�
>&K�S��z�FF��oFO.F��gn0�U��5�Z6�z����B5���~�LMu������x��+�SW�v^�Us����K�������$��
 ��=�y�1�I�C�}����NE�aLg��^��?%
#� "3{
pPӼ�s�ƻ�l�夜 L Hṡ���6���ǜ�$<�,}�OHb�Ck4�/�Cps ř9��y!�D�@����(eڈw�8Ԙ��A��lk
3K���Yۨq�eq9�(q��Y��#K&׮�n�C~�Z��rr0�/#$?�����J��\؄ku�*���.�1�P�CZ���!r���t����F��ѽ3�,V.BV��qO������c$c��m*
����}�f�୑n�y.xÌP����\�g%�����%�+�N�T�;�^�CO7*՚N�0!TQ���M��!$+(�rb��mw7��ydT���}*l<�}8Bb�Ei�&�~aΜ�%a�\�q��g/$u����Wf5p�݌��F!x���z·YuX2�']N���0�*`0Zl��䡊��EIP�q�j������r��+��.�0V�4X��������\��b�����2�i!�]gp��ȹq��0��E�ڮ�n��W
��
�Xk��ڥm��J�֪�W���A�l�o4`Q���5�Y[������� `Ei����4 ;��n��R����ƴ�!�m����q���.6r'HZ��8ƨT��Ċ�D˔.�t�@�iN���j8��GF���[����`P&��y�pl�"�_%O�f�L�չ��  `Rb��-��VS�ٻ��J�pj I� G���I"@�@��q.S*�%Ad�E�n2&C5Y$B�5
�F��@�d�G 	�H��)�qj	 \ut�:�Tr�L�D$��� �##S2�ɐ+)]YW*.�BDnj$�	��L���p�b�����mX���	0'�65]�} �}�G�h�Gt>r��,0�M�S�ѻZ�>1ä���b�ψP�8����wۮ"����Ƃ/P���q�B�w�Bz��${�t�cgoCd���Ն:p�hIEY��u��=�}`�Xa�ֆ4M��YZ��x�!դC�$�hš�R���-T:�� ��`�6!3-�6,�H}@�ꆝ�"�!ϺŻ�;�P��)~������)�Q�Cԗ��$�6e�㦋�N�`����^)��h���m�_oj��P����ڈ����m���}�&�K���<_��&8|�>#H�*K�ы��H�r/i�W���*Z݀�^�6��I���"�g��bb0���z��B�,\��gXF��w��|A��2W��VC���W��4�Q�#B0t�q�TfY<Uf��dpن����ϸ�FJ|����/7���-4}��hR}�=rL��������!���,�@hC������zC��B��KO�����2R E�������1�8�����j�,8����Wz�5��&�X�F�Tvi���s��:�H{H9���*�Y9.��$١���2E1�u�$YӸ��E5��h0}�HwA,�
�$͠�ʶ���2w�� ���Qs�:y���ѐ�6ܐ,ٓ�.�iDF�qW
�oJx���Z����d�"���$�L�
�����,1�4/#&��E���!v�Fۜ#�Z}��IhB
"�q��p�����b�ϸ�D�e�� �	V��΍�t���50`X�0�E�-�'RGeZ�Z�-a���/cٍ�.h�/\ �WB�m��Y�,�i~QсVD
�"�]�J�.��ՙ{Ɖo�1]#�\�܍�q[��X���M#:v�!�J��ȩ��~G�������8t��l.h���Ӥ�d� :^E���k�|���`nIձ��+>`h��9��ZEPde������)���=GӉ�)��Ƃ/I��uq�/�����*���ܛ�TkCmi&�ҲKj� 9�6�t�),p�2o�5Ybm0#22,u��IE�L������1B��V�K8p�J,p�!Qr*1�!�*��Ύ����*B�cR�᲻UBi%��*{��'v�f�]�$���������F�����Z����%���Iq����׵݀�`	�A��0��2F��>�z��#�YkCH�XDհfT|���zё�P���6�"M���<p�2k���׻��$6�4\��4�!��d0�C{h������J2J�a"��/��V���P��F1�@AD$*�1������l\�� �k5HzO�� �/�J9�����_�ͅ����aDGȆ5b���WHi�@�x�!e�FC�������?��WGP#�Uh��������pT��L��
�a����={+�hC6h�Z�8�v�SE�ZFZ�D	�ڜ�x�4x#N��+HÔ��i��'�=����{Ju��hMn�\��(cx�]���8��2[CkZ�ƴv����!�I`\�59̤�vl�2F�Ʀ�í���(��i�}��5��N�(ABbڇ�`�M�(�5%X�r����l�~`�/YP�������A`�D�DA�>�ZTYNN�1e�lO���.F%"K>�z۰�c�J�o�H��4��g����}{�pϮ�P�'=4x&7]d��X<<�`��6+����9K��5�(��=t��}НHFޱ���,�R�'��"2'',"a)Ξ#C�,;X5�
$FX�e�}5� a��T�"��Ř8l�C��������f�H��Ȣ��\�����]t�2几����q��
p�K��7TP�ZE��!���Qpx��sc�
�"��L�a��0\�.D\�ڇ���d4�:����(�cz�ע�6b5��D�	nw	2C��� Lﱯ�B��D�7)�n
3dĬa��I�ːmn�H�C�Df�y:V���&1�FCM�X�l�#���K�G��%�yڅ�Zh�������Q>�RB�$�̇04!o���f��^R�x�"ϚԖ��-���'d�t�k8GH�qG�bB��N&��",� ��M�293U����%�^�Ǫ6}���P��x�����l5�7w*9��|DQ&���,{P�^��h8`��u	u���@�a�|1mO��B�W��='���r�m���e>1�����l�a�
#�!,��>�.O?DA�cSX�����E��a��c�x�8��0QYg*��b�fٖ[�L�(qnB)Q��6I�$�A �{e�nP�����F����t�>ؗ�,����Q��Q�Q�)V��J����\�}E�9��M[
,%
榲y�#�d����Q}��,d�OX�����B�&�#��LC#01�o%��L�D]saV�>E��t!�0}N�6��ƣ�Q�7����̙>�0�Lt/�p^�G���kk�\�0F���0�"���$A��T6v�ĊM\j�Z%^��番��k ���!�]]vTΨ���!��x��4p�����u�DA�>t�5��������xk<Cj^��t��I�f��-F�2��s����"������u�]�)��C��ӂ��`�A ���@��i�+"I'��VgP�0�������q!Ir݄���c&U&٘��l�>��xJ��X���j�����\����P��(��<f��kf�����J��<d�#���`�mޜ.Pt4� ���7� ��˙"�����䏎��w�u���G`��Xo'��t٠E�i</b|��˔�օ)������tc�۵��v����΅�B]j1DzR��=B�G����w�̎S�&��b�뵋N<ԕ�\Ȣ����R���:>�mQ�P�}�q��N�leh9��J�n�����"Y��O�#:p�̵���_���&s[B�L9� ����bm�α�m꡷f�^T�{��pU�i�*,�]�
y(�Z���k��*���IK�34%��sf:��1�51�b��I����ޫ	G��1�֚cr�QѢ� ��K8//VX�G|N6��RĺĄV.�u��/>c���|��̦)vV�p�����'Ñ\)�V��;tW�s���h�A�)]�̵����*Br����e�mWA��L�˪���^�	�� ���Kf�Ȝ7
�i=��`�Q6v��,n��HŖheK��   `+v`��V��YS�`kz�Tf��]��rA���Q��K� �
ڇ#��FA&�Z����	$�ȕT��MD��R\j!UL�#p���Ÿ
	���JI �̱�Re5��.Q�R�]Q!!��Ԩfe�C"H�i �\��"��$ŏ�"FeIfSW)#���YtHkXZd�T���!Y�V��&Cr�9C	�8�ӹ��9lɳ�|q��Lt �(��6GRl=����E��������
u����e����r0��D�Ha���B.v�51�Tw�x��.`�-( .�'���e�˓�4l�)>�A��O�����緽�X�9\��m0�ܨͯQ�\���;QqaDq�H�NkV����Jr�l�1QH�Q��4[��0�q�8j�&��X���,F�u1��l�8�$@~��6)����0D:���z�g.�f�/��j�)X�H��B��rZ��=UQX&/Ch<��뙘'u(�T�2�r�j��ψ"��jd�-���PCЂ�`լM�6@r�Ξ�w��cl�b�*��n^�B��l���x�4X�:`�c�^XQ�d�g���l'w���=!fJ�.��ce�!�"[��[�w��Bd���1���4�a�+r5C�n~��ިe���<hپ"����Rw��MN;�b�5���m0�A�i��.}y�t��C9"�C��ȊZ�ar&��TojLk[��c`�@��2p��%�b��L��:��|IlV�CS��g���u)O�BLN3�tS
�NV]s0��Y:�^�Z�e\c�6�I�{U�@h�M���3\WYC�\��ܓ��j:}r��q<�WuT]e��a��ڬ���d�xơ���ɶ���:`��Zu���-Ő.W��o�Q�4 ݮh6�a���<1�,�DIE5[s�����\D:�N4I����yΪo!����PBgN,,}���*[2��(�Aȇ\\�,`��	6�~�����+�t�
�ō��a�����we햵[k�wu���%�%2k�Ƀ���D�3�DV�D��ؕ��1B�c��0Y���vJ�\�wr;k��Y��Q��;�v�"� ��׶�}-����/Vt���rT1,�˳ֽ��;`�a�A�i��s�;KaeR�q�܅���ʋ:�Ð���=�n:�^�y���L�`����Ɏ&��J���s���\C�d�D�d��Aj"��3�q�Ng���l�!	"ƾ#�4�!7���Pb�uG��l�C�g*��@R��8*S�8�&�a`��2W=޹�y�[�*2h�u6�P�
�%|���AeN�P��b��I`G!ȃ����ʲn)�'�OC����2ʢ�h�+w{H�w�V�WL��OA�"U{L��<���e�".���ͶyG!@������}��D:��F0q���5��GC��H.Bءe��:��Dj��/6��f'l���ya���$�D�3j�S>���\���I�vbX���DAh�j���b3d'��)�CL�
�������{}�q�ǎ���3����S�副f�N����}^F��$��c�z%�a�����\��r��H�0�[bz��>�4[�%�Rh��Ogm����:F��ao����a��Q�XE�����o�A-��;+��!�m���S��AuA]3�$9W��7_��d%��u�e'4������q<�Y�}�&�FO��̘�k.EN0��{���B-�625AJ�D�Ys��u_J鍶��YTKY�Cm��l��h���/,��,-�Ko7p�ç�D��C�oOd�6���r��A�m�d^�,A0]���s^���BX�4������ꡡ��[Lh�#�r����!�B��[�_$v�6oW��6���Xђo^��-��t/=-��L/(RE�$�	�VY��	�!�O�b��sS��+`ux H�,����f#��n�L/�b�2>�����ݘ�U]�B|���·#
=������N�#�MFSh���jsd3�)i�B�5��`�4ds�G��0�P��v�5�iqdT0ax�(R�Z�X�DX4V�#(H����pC��yj�N�� �!���\ݩ9�ǟ�l���a��aO��aj�Eiy�x1*=��Z�S�<d�U��/*�qp�Z^�(3�<�)#q9���㵌5��1��A��峖+-��9Cid�0��Z`�&q"E���B�y�>�B9�DΰÆ�$r����L؃`��eP{ǥ9��g�0R���!��N�-����jj���2�3�-�4��rD,C.r��X�ͪ�[��"�l�G�p�u$Qb8�8iл��}��\�b,�z���!R��r��o1�nЯ��ɢwa��#*�_m��jW��4u:{q"5z���0X�j���i���em�!͑`�(6C�܅��D4��a�),����(�2h��)/q�Τ����5�$�f�"����L4�� �&K"gr��u����1����m"b��d�"H���~t�M�l"��e��&�
^�N\�� �m�wL[�I����ewwVhU��Y���!ò���@:~��m�Aw��F�{�݊�/aJ8�cG���,�׫瑤i��*P���,aZ�塆]Y��㌠&n����B!Θ2CńX�k"���M穀�(����9��P{B[�[�ƥrE��D���>E�w^ҍ�*,�����/7c��,��s("2����c�Q��e��"M��P�&��y���A�{(,RaQ�A�!T�4D{m�ׅ��&�]��@����(-(Ll�4�'�a5��Ne�r$�,��`΃��V5L-�q2�&fT�LS\ˮg����Xʸ]>�23�L�dw��v��8�z��.(C\dRX�瘩ZG�g4/K�ӡdIo%�ˬ��Ƹ�/9��M�g��8E��"0(��챭l5����٣�NJ�*|�������0��������	zn1a�E�X�;����D9!��Ơ����p׽/�*�H�c� 9��m,�SNlvQә�:O
%{yQ6�q��s�NEl�{��6������7�a��l���HQ9�0s�F�ٜ(_C6l�\E�>� ����-�K��ب����F�։�yb��⢮����]�7���q����NɌ|��p�S�
�O�G+�;[h��²/I3���@�����6k�c��f�쏟
V��o(�!W>�[���&a{��%�����ti&\G{t�ʑ�ovt���Q�Wl75*4h̫Rav�� �(���\<p#&gc�\v�h--�x�l��y��PYx/O-��B���$���Y/��ɬ��5�`)��������g��w��o�������-�l�/9�٦n[�m�t�"�]��Q �۫b����:�O?��;ה�*@���豞�k��Q�-ɋw$_`���R�)K��W{��d������ָ�7F�8j�T�y�Lzc�+k
�to��TڝR�=�}�DJ�8Vs�C��a��K0L-m��i�hL����B���M�X���:�"���z=��A�ud���5yLlSz�����Μ.�ͰE��<���+�h$0����ƺؽ�(�UJQ3~�ם�ze�vT͒ķ�
����9���Sx�    .�ك/1Y�٫r;�X�*E��N�yuyY{�dc�����`Qv^%Ģ3$��'��Y �ϝ��	 ��)}����0A�`S2�N��ɐ%������Qd22%05�d���(If��|�$;&A�< 	
� j!xT��$��eԗ2�`��$D2 8( �>#6v���v#�"�� �X5�9f�S�����ܹ�����i��ZE�t@��3J*#+�b�Q���b��t)��S�z��ǒ`�-dm!&J�'�e���Jv��=�(��`C{��Ō�byIP��%Fl�9`�4���1��Z���m�l�Ԧ�;6�9�'\C�����
�`�1I[���g�n�!��E�~��iqr��Ɲ��C7.ScyQ�BH���W)!�!/,0�c���Ķ�"�IC�\��ܓ��&�EU_k�je���w�)��=hM[{�Yb	��q��h=�۟����<4آ�]NK3�p�����2v��0RQP��ȕnu�����r�$)~�//��_�K�� �>ڽ���uֈgX!nh ��N��Y��-W��Bi��"T�
�<f��g�Br�^�Xr6k���b��!-:�9M��9�9�8���D<�r��;�Nb+Z�L�'��7��.f���H�ƧU!�3M���Q2t�/)���!��޵�u_.\�:��"g�Q��k2D���v�Q�CK{L�?;�SK�W_��K�����E<�vn�ל�����,�y�23��б4N�4���X��;�N]mXIXYNb�:�V�ݵz���ZF$ĕ�Ԫ��œ]�)�l\8G�dN��z��c||�(��H�~�|�7�^�\2����U�9����8�����+�u�<�"e�wc_c�����c{K�s$�"�XS���s{+7�e0uw7��=�����^t���瞞���ݽBY�)q�ټ�mM޲WVm��)������z�Wn[��T�Ծ�Y[���DUs��y~Ɏx��,O/�3D�
|�S�fVb�+v�J��
 � �N-�/iw+#P�O,�@�ܛ�3�l����+G���^\O�{1=V^�s%�{	gŐ��x^����+���gO����'���2�`�����\�Ia������ݞ�����±N��]�y���U*^~@W�h3�V�̬�/��.%B�o̶dl��@�<$���8�{Uhú�k����o�����s��&_=s1�#w�����x��&-�C�4֣7�J��~���|]�9+Zq�̷��LND|Փ6�`�c�^�y��ѩ���"yv�e�N�� ռw���)٢��s菵V�c�<Q�٫}��]���<z���VW�%
�UӄL�0=�Ē�i�lZ�$d{=\e��ֆ4v�ۉ�W�GgO��'EW՜d�OS�4T����ūq�W�3޶�qR*����xh�/��ɸz��O]�x迋Uj�O�4��]W5>�ⶻ�Ҝ�{��㤌�F��m+��:��]�G��Ȝ���J��n��F�^��k�mϞڵت�ЇO�,��m��Ù�55m�P�W�euE��A�����8Oo�:K|캐{Vy�n��o�zQ�)x��:�9�8,�j��zk��Sl�]��9�j�%S�|���.d}.�T���.h�sc�+.���zfL� ׽���=�<��!\�{���}g��p3r��+S��}CaꞮ�+i���)G��}��d{�;6@��,�m[��k��!��4�SuV���}Ε�|�qЮ��4�\����l;�����̋8�m�q�4���oPק�����٭x�S�^AL:=��dU�/�S��@o�U�&�W�l���):z6�d#�3}�������=���;E��h�UM���0�b���2J9x�b������X4�K�v���
�@b�S�%�{+|q���n�h�v�{����V_c���R�*6-�MٰZu-�0x�C����Ł��dm�S�sz{.����-��(���wxP�9��ﳝ��32�gO����De�4�#�,xWq�����xoE�Χ^v0��S�#�Aթm�zó^s[�K�}��}���u�;~�]�2�����ۤl�b�اl������]%�ޣkA���9꠶>��'�0��D"V0ӹSIb6��҆��]^b�Y卙��]Q4�����#=2�-��JJ^�����w^���^�Dฅx1���wF(�h�~2'lw���"���No��K٠����h�'�a0z��FI��K�sm[=�s�٢%4�t��~�H�i:[�oh���5�����t��܍�%(��wH%���ڑ�8���_���~�Y$;��RI$�I$��A@D�T{?4O��h8 �"r��BM���݄
�Mo�o
rm^gVx�`�17�g5�C[�0!�F]@TZ "��y�� �t������7.���t��p�A������;&�g���W!�-�r�Ifɭ�B�� ^Po��~�m��ݱe��n��û�(Ie�..����!�$O�y}g�q�!>B�w�E@D�����'��	��S��&{G���?���`}���G�������Oi��:����A@D�~����a��B�Kg�o�u� >��o�p�4p_�Z�	_�1*�W��5��{ �;=���t3��װCb��"���ذI�S�L�u}r�ӛ�D(4*���D*
*��&����Qe:V�Yg��p��� �p�{�P9���	���b����q���h�%v���T�Y��u�Oa��q3�i��Q�y�i�ɿ�7~4t�Њ&����2�����W�G�؝_��Q�è۲�8�@�n�z����6�����C؆����:����_5=��A��>��u�@(�I�D�7�|}B�}'=���Y!������#�@tPPD�K��@D��C�}�|��m���(��撅z�v?��D6���$���N�X~f�:I�QA�.�N����xl�>��8�6��n��[Sm�=���pkFo-7XSB(�_q�{��v����0�<T�B C���)�A��ט�C�ǰ�����Ρ�[����('�z!��zD�r<_.R'�> >���ӛ�3��B�P;�cٮ��v
|��O/�zOh
%/�A��&������8�#�/���/7�[:���]��Ȑ����aa6��M] ��{��o x=�wl����7!�����@D���{�[�R���Yҽ8l��{��8N�z�|h�΍�Wn�@b%�:�r^�,E@D�C<�<���]�W�y����w��z�P= w#֑69�'��!�kL�)�C[��i�Ѱ����P'�.h�����"�(H+`�P 