BZh91AY&SYH� "ܨ_�pp���"ߠ����  bB��           ����@mT� 
 
  (Q*�U(PV�B�h4  � 5�-C@(6PgA�k��n;0��P��%Pɣ,�	kZ�6�H*�e5J�%@$��1h4[iZ��m��Rئ��f��   ���QK�2� Wl� �  ��� 
�rGT�\5ـ���@�t�RP �p���b�T�NA݁�ճ��>�	I)o{�w@��XIf�j*Aj��c%QCVش��uQU�k��&B�i��֕
�j��J���Z�=����k@H$�k�@�_Sj��{z��4�u-^���mSUM��mkm����{��6�[�n�����*���'�׽�j�C��{ٽۻv뵁�^��G8����o�Pu@�K�J��M��B�X
�5�Pa���t7cs�hx�ޅ-���gx�����N���wG�5�x��	[(���Zi��7�y�^�iK۠����Jlǻv��o<jZ����J��Wl�.,�
i[�P�� .o�>�ѫ[}�wL�۷�tu�e��e�b�ګ�t�{�J��������z�R���*��+��UgC���;+V.�t�i�in�p��w�n����4�f�F�+%� 5��{eQ�);���w+��kc����f����oq����d��޶�֤�wv�멳Z�W8Uݭ�݇5v֝:j�+����b3n�-�t�Mip]�eU�T��$�F��ꪕݾ}A�UՋ9�Jwm[�=x�t��T�� �6��2�졧p�ֻ�����m�J���s(m�X��:^�R����F�*A��@� h [�}�UP�1���ʽ���� u�6�6�]d�[�ժ4��ƀ8�庭���M�l]�s�s:ե�n�+��
Н��Z����AB�)wrݫ�PH��{�R�7]��{m��=�]P�ot^�.�F��c�	����w�E��W���a�r��ꆙ�ҕV�v��SLpfv�S�S�SCIU�
^3�P��I�GޔU}3\�)E0�ݡ�Uj˜wj�t8Ǯ��=gu�Uje�i*uj����u
̀uM�N:�N̬�#� �*�m���W�T��n�C����A@�U�s���T�	]qn�U c�n]As��.�wM��AZ��wj��M�  Tt  � 50T���z@ `F�@5OR�@      T��U)C� L   O�U@�A�@  � $�J��� @  � EzJ��F��$��ѠzG����l�����y���߼�[hO��\�8�w���ӗ��Y��g�_5�b]=�;�~�� $��6����}��@�OdG�D�$�� I���	�'�����^����m��� ?����U[m�m+o�HH��������?%?���AO�S�0���vjaL,���f��S0�˅0�tS0�eaL,�Q���h�,��,°�
�Y�l�
ac
0����0���X豅�avS
�Q�XaG�¤0�#$�XY$0�L)#
�
I����0�&$adI���$"aHaA�A��TTL)&PaRL,�0�L(�,&A��0�*I���aa0�0�,(�,�
�aRX�
�aA�I0�¢0�0�MY$ ��K$�RRL,*;*F��XD�ȘXY��L,C�ɅD�TPtXTL)&A��a]�!�!�I0�'EI0�&QT��$
�D�Pad�
C��&$�PaL,�K"ad&�A��0�&PaA���0�&!�$a`aRL,�"0��E�(0�&
)&�Da`aI0�&�X����,��H�d�ĘPaA��ad��PaI0�0�0�aa;,0�0�L(:,I��L,&$��;0ԃ
�tPaRL,,�
$��H0�&I0�&$¤�Y$aQ<+
I��M����0��$�PaRO��0�6X� aa0�&!��aRTR�#
$¢0�0�&�$�ĘY$��abL,I�A�I0�&�!�HaI0�¤�TY$��0�����&�*I���A��ab&D�K$�PabT�'EH��0��l�&$�&A���I0�E�0�0�&HaI;*I��aA���ȘY$��#aA�I<,�aRL,�
�a`記X�X�
�I��L,&!��0��L**,���0�0���,*I�D¤�X���0�$��&$��:)0�I��L*I��d�
*&PaQ0�0�0�$��&
(tT0�0��ē"N�L*I4Y#FA��0�I���XZY��Y�af��V�0�.�¦0�ag��Y��]���,��,��0�
ac0����Y�tS0�aXY�aL,�JY�F��)��Y�af��Y�aL+0�Jaf��S0�aa��&�Y��X�Ʌ���)��*aSeac
�Q�OJac��e�)a������X0�aO50�
tX��,��,X½,¦��,afafaXX��,Y��vj0��L*:,��+EVaL,��K0�Eaf0���0�K0��
Y��V��,°�eS0�<,��+0���f�0����0�
aXS�p�E0�
��,��+0�U)��Y��Y�aL+0�,��,��,aL,�YK0��T°�0�,���L+0�,ac0�,��Y�0�,��,��
Y�豅L(����g��,��,��)�;.¦N��Th��,��,��KS0��p�aL,�aZ�}���0��G���)~�(h��x�ƪ��b�ԺD�ghE�lR���� �l1op]���!����Ӎ�Go���TJ�-@�6a���n�Sk7d۲�Q�٭W�^VX��'z�x�Ū�-���Qr姧v�wY㷗��[��Nݫ�b(�i��K���׊�>�D�S�-���i��u�6��M�J�UOmK�b�ѫ�p᜼���Y��5i�J�]K��AT$2U��V�V��ݭ��J��I�ʕR0�����ɢ��۲C!�v.�	eQ�I�r�ݱ5�,���~���v��q�8�tOP��W7�h��t�mlU�5��ö�f�6�j�fL��r�̤kf��\�;{l�%T�bEV�ݴ�M� ��f�w�8��Z��Yq����,^����C�#�hҪ��D�P6� wch�
���YtU�j���i�>���Ϳ��/e�	�]"�2�$�^%�,3 �#�o������o
��U��{��t�z���z��ťG"1�T)�E��
֪6*�f��3h�Z���{R�]n)��Θ��٤髵uS[�n��T���6�q`:�T4�YZ�glm"�ΤN�8W'@λ�t�-��p��1�/]��V6݂��n���:�R�S�hmhi�fHv=�}��T̤
���ܶ��T[��#(ad��:pY6�^�ܘ��G��G6��ct�;v�+/u�qͩ��[�V��d]i�<&c�z���
rG1v9���ͫU����
�Y�dc�2U���e�����3\%��,��.g,�%5���*]g7Nd��xBś���bkV��\8*�Y�<��c�#@�gub':w=|�9�+��:d�n���i��K�I���X�)	�S�(֥�	J���pcbE)�^�%qӗ����
-�.�^d8�h�0%� ��B!��/]�f��o2��4)R�ɬ��J�"�2Faڳ�m���-\�n-�CM]mB�m��Q�T���p�J0zz�`��(:TSnq�Z�Y%�n�����3"R�E_;ʹ}���k�j^���;q�oѷp^4�̘����s,S��X�2�����Ҏ⠺>���ț�Ϭ��)�T��H�\�iо��כn�5ģ�����ܱ�׭-��;/�]}�r,���K-U��N��j�D&�2�nQ+^�"ʋ�v4�[4R��A��Q1�CJ��#pRT�J�nr�4<x����(J:�=�˩�^ Y˖�>���;]��8�u���C^����ڤl��dw�9y��aUm[.��V�<I��K�Bh�fHXYf���dOZ�u��*�hb��-�sR�V��e�6ӧ3s���g��Y�3��ӂB0L��"�7�����Vػ�2���
+l;�x�㏶�b�S�T�US��d^�,���c�OULdڇ�y��U��]��v���%��M�eu��.�͖���D���W��e��Y�=cr�^F��+*�:�#sx=y�����۬ʩwZ�GQ�:�l�v��j:�.�^Խ��af��!�ٳ�H��P;H4m�8�b�y2�2_L�������#����ʮ1�ސ����-\�{(��K٥6�)M�vQ'��#���keK˷��SMe�Seq���^R6��
�i��o`tXܦb����ktM�����X톰�+e5���l�W�����[/�B��
LM�
�1^Ѹ���k.��
�y��fܬ�$�����*��V
7ha;��E���,b����7s-�b��m�n�4n-�횂8��v�*ۮ�B1{��Ѽ���ՌEuj���ˠ��]�ν{�.�G$1l�Cm-�{z�B��e3|,�̳2�r��u�էb�<X3(��䫅�Y�$�+.̶�"���pz��5&�M�n�BӇ*�ݜ)¢�l:�{+fm!�T�i�l�q�VozA��k�	켼�d����	)���d�WPn<�&V�ѱsU���ŘE{Ϋ�cf��V���ʔ���K�W�#��G���*^;�F�̗
u���d��:��
�u,��j�ӵv�Qޜ��:�*�[�!�Up(�EV�M��L,��;}|9)66$�Iʮ�*�l��;x*��<6{�`�/��skF6wwP̻J��E:�L��u���z��VVҘ�elH�Y�0�
�أ�[��[B�TL��Lxe��Y�0]#bt������s1e�R�wZ�;z@uX��8�8i=�Bf@���r�q��b�v�s�Ym#�0�T��j%t�G�kcX�]R�G2L�.�c�Bk(ޥ(��U�J���Ӡ���'B��X�+b�V�F�c;�]�+u�fd�4�d[�^\`(�ɝRU�b�n}�ƻsoe,�na9���Ɯ�RX����ƞݜ��0Ub�^�L]�v����f�м���t�^=�	��{Ub��6��`��ˏF��e<�Ƥ!'��&mM̍��Jj�e5��7Xڬ��n�ɮd�[����a2�s��p��q	I��l�P/=r���0r�r��vĴК��S&b�
l`�w+%J0�vm�61hR��*2J�u��WK!4�5��
5-"o>�A9ݻYFb1J�w�'	$4ov��.�k�=�߯g��i��AxJ�z6��Cm8�Ke�Rd��"�p�p�e+��C��EZy+��E�A��^��/p�E��4ռ��ԩy�UZ,k)`�L�F	�:娨֜�4L��sN b�cɕC7��f�"����kt����$ ��Q�f{Q����I�me��u��-[������Rb�j�ܝR*f��Os)�^j�Y×�5��d��lԤ3�Ʃ��$�i���9���{h!2м���Z���I�"Mnuh�Qw�[��՚�T�&���l�X�pv�̭�\�
8p��`�khL�AJ�E�S�Q1t�Yo6�^]�Ys1�wY�u�e�rT�����R�t����Ԡ�Z-���IJu1��P�m-:(��f=�ͱ}�Ob\�4Yu*޴�޻C	y
{졢��7�[U�d˥�Pn�+B�E��O�3��#%��C��^5�⭺��'��eLc=�C-��nh�U��I� �ɱ�+7-�mDD��ة�zk���Zv1n�qGyz�mre���Bie�*��w+��"0B�ʍ��N:�}��+�kvX9��'+[�FQӕ,D3JɑP��˔������q2>Y\zc':���*�{Z$4VR*n���c:/Z��hf<wl!we����5G����w�����|]!4��Y�*KR�eҶ���p�DM�6�`��5��7wZ�T�ѽ�F�,��U'Mqn�wm]I�v�=V^�[�W�$5N.��fe��$IޑU{���%M�Y�ZF�u�l��*�;����6�6ޖ�Հ�5WK#��*}٘z�zv3s̨q1v�%�^*;z �S�R��j^�A��Q�3vK�Ә�d�( ҬI悝���0��K�5���I��ُ3/s]�r�;�:4��T�$�Ά��&�@ Н�S]n�N�)�w5��u��ObSc�Xp�a�/ar��F�7�Θ7���/0mTZ�[õ�~���7Pi�����<N&��Z�$mɷ�Ɲz�9w�|�@�n'u�\���m�s��u�U%��Nb[{�j����b�y���9.�~���U1�7��d�����0�y�{J�nD���/�2<J��8��J�lB3��c���0�-0Pn�ˋX!���T��r��
T�I��*�{F�5��[l��|K�a8R��]�ӹ�,C7K+Qr�1�I	6&нŻw�ξu�{ڇa�Ƃ`���a+Reh1����eQXҧS#%�b*جq�!�+����闶d�t!�i��F���*���Nm��v��.^T�Y��3!,J^%�)L��fꄢ,u�M��o1��jHݥ!�[�tӔ�̍��GD7[����N�e�$���f�aQ�]���qMٖ��6���T��l�;����WW����6<;fGϴ�ȕ��-'woa�O��1�����,��Q�ո-'���o��R��-�����oc���m��(��![�X�DFɎ�c��Q7x�:پ}SJd٤�r�zr�M͢d$=V���u+��^od�Ʃ�s$*�ݚ�tD̩Y%��e�y��(��n�n�7[o,ջ͊����P�l��řuCp�J�u��u��F�l*"��i�����^ۼyJ��ȧc���x~�3n))�Nm�.�gGز��S�Y(�ya> �-�fR,�����i�O3lm��=&�"�3r!3�=W;��w��MZH��Vɡ���5��n5fY�ɹ�n��Y5�=FR�'�ZkS�p^:ŵ�(JȆEV�;R�M�jR�8V�nژ�n�Y�K-\�Ң)��۩�Y:\/4�!����Pq��Mf=�Yj�V�u[�vO("�c{b/�V��z���pT���n�*�D7rJv�i�,[����nN�MR<wY��m��֯)�.�n4Xb�Ne`x��ӵyD���ه-�6�lV:����4]k�Oy���M�!lmn�ReԀ�a��X�RAٛyo/�f뎑{�1���ۖ-�C$�� ��-�����g&X�w����&�݊6!������NOef���س�f��f=����Ͱ�"�/J�!卬37��[�1pz	�v4�3]L��wP�k/ҖK�Ckl�cԱ��J��Lȯ'�Y��|���%�U�ņU��&>����2��Y�;��/5�Xw-�
�=i����Ý��Q<
U�K�T
XA�����b�F�m���H�ڶÚ���e�f�Ֆ��pv�"AB�*��S
��Y�U5�"J5�T���^�"�*M=v��>RՔ�|#�)��Ѥj���uuB�1�-�y{*;-҇�cF�xs[=i��ޥ¶�Mtwm�x�%Xu��\�+Fn�J7ugF�ǵlʅ�k%��|�����\�]�5pZ�Ir�u��Y5��(*�oU��,��ܖ���R��WWl�'Z����*(�/���^.��zk%���H�ѵ�bP�Z�Ux/V��C�i&��z��֓�6�C�Z}��V۶`t뒬(��)���B����ID��J�c�w���3��/��s
ݗ�\�̂o�fno"�V	U3a����t��9x�9�c8�ɒ����fJҘ)�:�ݩUiE��7EQ��fjХ��ӂ7:���se�SnE�l0�4(�r\�Xc2�!���:6�!k��i�T�,Fb��ܖ�"T�������= �+�ВÑ�R��T�HmJJ��r�&ͳ�(!(&�M�W<c%nˢ-Q�:�4�*ǧ2�켾$��tw8Ô�q�/졑��"���^�5;v��l���g6^ʛ�j�\4[ʹ�R��Iǰ1׻\e�[N��X��R�O�⪫OfKv����uʥ�z�<����\���#�T��NZ��᧐]�W�7�ȣc:�Jw3F)��<W�rh�-��GI�J�%���%wKT��� �	���VP{�]l��d�mk��V���iR$�bVJ�k-��j�Y�4W=�X�G�(͏���n�*݃6ԑH�fݔv��A�Ւ�GR];E,�l�Ydк�OA[�S������D i�'S���6��~\n�3QuA�G0�/�%V!E�-�%>ȕ�p�H"��#��Xs׎[W6�V�P�2��tӶ�s"9e����"�tͰa\�TX��ݹ2�Gۨ�f5�w5sj��{[cl�o2�y��k�R]5��7mJ�1��'-�*㮠�h0��z�wrVH�v��rma�d��Lv��7uc���zo|����$-*�B���X:a�'�p�A���C�@U����1ca�1 ��>E��H(����6@�B~D��l@�,X7A�08�d	PtE�[�&È$��*���-��u�o���.�u�c'���7�(@a�j�[`�z/uXi>��]
��>LE�X@�7��/V`�R`-�(\b6B���ng�,XoC�f`���9`�E�����~�2���sX��]
�U@�|A�1�IX�b4�z(У��ڨMh��a��
�ӂ�C�%![���,<�n��
�#a)��1�=�]�)��h\���=�|������o�2*XǢ ��X��W�e��x�u���u��b��@��r#��`��{(e/b�`��C������:pvУBD}hJ��z|�	�'m�L^������9����'�!�����["VDv!p�PT�ףC� �FN�4&ta!���cfB��>��cS��|�3E憐@�>Z1P���DS�*�T1`[~��h����HMC$��B�F�PăG�b��;�C/�,.���vA-��3���ׂ���;~z+P�"��B.hH}}����へA�-!���@t5p��3S�.�E�8�3C%�S��O��6`v��	�qRÝ���;��c��r5�J�}`F���"�/�,]��p����;8}�_�a��>���X�b�Ķ�X�c��`7�퉔�QQ����i����+�`cd@>�����0j"���U�9↪	0��Z!��b�� ��;X�c��m�� ��.�k$4���zЅ����ՋDZ!��d�
"H<D��dg0-")t;�D�*@>�
 ����1����[�B����bB�(%�*�2�j��8U����M�`��1��ds�j(\�%�q�������쏗��PƂlE���%�@�0U@��Ţ�Lr~4�W�C�c�DHEcs�Ghd`]C�B�D��qbt��1OJ�b��)1��_x�͈�2P�Ńx;(s ����3���cn
�p���x�9�q!i
H+�N�8"lgO��1ż�r�D;�\1�X&(^x\ōt9�G�&|`�	h:�-���¢�AkA
�E@9������6&���g������	A@jB刨[��B/��!ˊ�Hs��o	��?��I~�x~��~������������&��c���䔛m��m��m��O4�Uw{�2�6�m�m��a��m���e�m�޶���۶T�Kn�m�m�p�-6�L6�Nl6�m����ݰ��2�!��Q����[�VvM��cqL�S+�E2�S�m�0�V�&A�V\a�
N&˰ylܼ���*@�Q���k�J�tk�wC�9P��~-�Ԧ�Q��p�K.�\���j<&�jV�]Z�7��u��5"�;�I����7�QZf�Vl[�v�F���S��d����&�6�p�v��vv%]��'u�)�4�Op�Rͽ����r.P��7TN�h�9�oR��XZ�;i��2��m�ս�J���x��8��3^���5r�D�2�2��00���M&��uo]P�u�Φ
�`���^�"N�i�����`�iڵ�����VU�FE�UI�l�^+ڐ��v�ԝ����2�q�/FDklkZ���ؘڇֻ:X��i�ƒ��]�_B�r���uS�e�o���2���Sڛ�ʪ2F���H��0z�j%�G*+�3n�n��B�fB9ftL����Ԏ��m39�6^�[f��Yz'x�����Y4R�~�{��:Op�a�	T�*��C)��mu��.�y���a��p7}��aa���c�ۣZ�v��H:Y��`�	����r��[/̖M��k0'�]^!��v1.�R��p
���t�ᯞ�{r�	Č�I���n+�\�����1������b�J^���Pem�f�>s��$쪤� R"�^nkatY�mC���ЬZ�D�7��;r�q�W}h�f�+��s�y��d���W����u6lx�4��W��"�m�X�����Z�XE
Hl�4��,����ާ[aV�`hפ��U��W:Cv={�x�]��yƍf��}�U���XWXҨ͔��+m�YXVVA� h���r�*��A�_Z�m>�>Old�n�qde7A<�!t���y(�u��P�6^�T雱أ���Ν�RS����������ж�`%3I8�VƇ�N\h-�8�;�q֜����$ۥ��НN0��Ӆ�J�6���}�V����2�H�)V{,,�(j�zL����b�R����5��(��pI���r�����׶��u����մ.��/��#0)*���Os���%�YF�hʻa�Ӳ���Sp_==�F�4��V�7T���B��� P��em�$���b��Y��g��fN�H�˰bl����ը���3�Vsu*5����e]�$[�7�T�d�ר��'8�m�2�vr���W�e������+y���Q��������՛˥L�n�Y��[r��C]J^u�t�*�#�.�V�X�i��.p��F�1��Â���*E�h��b�ssYxIZ4�!���9PVµfJ��:҈uIA�8ynb�K�7%e���*�b\�M��i.���v�	�Z�xl]�%t,��2��̨Q���9�1�v���F�<lPn���T��*�=Au�{K��w�ꠛ���D�m�h#�h����m̢J�	�����ugC�dm�X(��9i���.aӪ��&�;U=4
7:x���j��S�6�G�2�c�(����I"�Zl��1H��,�L�UZ�F���AoIpv�
�y�ۄ�tҍ3�f��e�=2����s[���k�U�AzE[9x��굃U�]�o8��6��U��卛��*��5�]���kZ�PaO*�ǔ:].4�juQݖ�u��Y;ei�a���ˤ���]^�&��A��SV���2�r�m�,Z+*gK`���؛\��DGv���#�e�ĭ��<跨�a��7�.+�D�1�"��O�t��_fۼو��F&�])ܒ��{U8�	Ȝ�e�d8W��!}l�y����Gq��U�4�Qo$[cp�L�D�	�N�MX���A���]�T�ћ��(����̫s#��0�É�F�YB6p��Jqf��1;�極bmtp�ٴ�]�!y�T4�V�oA;�#.u��"tS��S���^9t�7�-Z�Iy�����z��R�Ŀ]��k�Vj)vY����'(Zͫ�m�r�V��s�υΐSξ�w]�S��3p�Ec�ܷznƽ�Q3w�[;���A�nM��B��CUY	��n�F��^F��ȝ�ĳ2��[��S�����W;Q���hU�g�� {��p�<�kF��f(������`!&-_�,H�ZK���t=;}2^�f��T��+L�v!��T4�U�+/��Eyu�M����6�7ap�B�9NF��9����kM�o�9���!;�z�T�};-�t��*�e�1�+ӆ���n���XT��|F�JO]z�d��m�Ia;��E�ލ��Ug6��;�Z�ͭ����FmD'vj�v��<�UW�6��NFK#����m`�κ��M欧ě}k^�q"9&��eִ��h�3j�'3(�I��2��5Y#�H/mH-Kj�3j��܉��C��Ͳ/)"�i�ed]�MɩU]n*�ZW1�q oa@��V�
��
+LMĬ۫V�i��6�h�p�[85����ʢ����Y�:�ʗ��N�ޥ��|��L���*tZ��ۦ��jN9]���,m�HN�gn����M��W1`�t��zꛝ}7�[&������w��e��	K�Uj(�IQ;9v�;�+��(Q�[�W��C�u�O�y�Ү�Ӫ7���Q!f�6k�a�/M��Q��h��RD��&ԙt�����0wN�*��'d��>���0�)x�T8m�ǯpa�qV�&��&�)o\&�^��s�1���w�J����6K��p,g�h���T{/vlG�d������7���%ǜ�@��*͵CwF%ty���id丩��dg5���N�tԴ�d�E�d� p���I��ǒ�bw�\�wP�Ļ!�r)�`����m62�t;BPp�{��	�l��J2"Z�2r�%��Np@Td+�Fu����eј�'��h��_WSf�ͭ��6u1�c�S����M�*�7����76��:P�<D�
᮶��y�.�9[6��v��lz�:���;W+n�*�Ն��Oh�Z�%W��y����2{B�y ��I/W�z3��2aT<�\磲��	��	sqB�I�D�9w���gk���6�F���m����N�2sd���//{j�ČE������Q�2��8͍�O��-�#��ך"��Dsy)kS�l�<u�,�O0+B��ɐ�6�j�E��Z*�n��r�����7���L@���D%����2Df�ڭ��,���2�����ζ�C[泲�eb��=�q�W3[�Pc�1ݕr#t�%
d��@�6)�X����`��i�޴"R��crnf3+yI��$X�Y���}Ea���j�h�9wc�x[%۝I���[hU<Z�W��O[[fuT�w^ѩ4�z�۷J�&�J�.�t�R*���u@�vy��B4��[��/��n�.S��G.�b��ʷ�l��-vD��.����[���fK��P���f�#)s�N�U&���Ɨ��)M+��A�ev�:�;�Z����8��zeV�zؾ.�6�J;[o����	Ӓ�s�&։�(پ�b�܎��h�۽�k���͆]<2�Rh�C]5�ܕ�`�"j�kL��-�,v�L�5�[��U.�>���)EJ;UH��j;[I�W/M���ƨ�0�L�n���p�P[L��3�E�ɉ"]�@�cr�.W��I2�T��#���S;�uk���Y���g��LH��;��i9���h�zi�_R�U�]^o(��<P��<U5�yv���Q��ɲ[�UJ/r��6�)���Y�b�w{V�R�.�T�M]S�Y������TYiu�����WϷtT�f�cZ�t��m���������q�L�-�4FIфU��&�Sx�M�KenZee�N���I��'�B��%3:)�Fko�+o6)�K�ۯ��кbv�[T�)���]�Q�Zn�c��>��'�Fˮ���d����um�D�z<��WK�uEϰ7�MVq��1��w�v].���]�sH�jv�
118�Ë�o!2�l��������}:��';�.��B����H�P��*�hͫLV2k6��xy�3$�9�������p�� �z(6[��S	Y�bA��&�MbH��w-�qo�,ˋ��h;�P�m<��w;�l���Yl��TP�j!V�ìR��������F�{v�<ޖ�D�lǬd���_�mUn�$4R�����.;���W�|�n���
2V2* �ܲY*۬fq�i�HWMr��թ.*��wf�Y��..⍾�BMv�K��H�F혬��2i�0.�2%qt��m�䘅��^��fK�[��0��{�u'�ev4k������1]��]T���՚�Ɋϟt-u?F�;z��[2�N�jHg'�;w~��Ƞ�N�*��i�
��v�8��vj�2��XJ�0q�z�ᓢ���*�b�'�O��CމL}��n����@�d���C	+nٺ;��V�B'K�����.Q4��Z7��������;m1Ƿ�wx�ejD����K)�ᒯL�Il�̇Vt�Z��L(���	����ՄJ}����U�#�L[ָܪ�w]<b��skB:j��HwD�܃sL��I-�.��d��6����~�F�>����}GT͂��*�,rWp/��;Xn-iyt�E)U��m��/YB����J�Wpj�p��~�N�u�ٳ9����vri���:�3����yX�`�5J���,5̺�r�3	�y6�"�MZ�W�Z�l�ceD7�LIvjT�7��/>�����m��䑇f3��tnV:���6@k�����N�U��dFTƛ�1���5���)]o��q�Q��SX���[^��E�x���I���н���X姷�"&6�C�W��a�Y��bwi9�����;�C#R	�� ����7L�ꞛ��-S��.JU�6���L�wkq�	:Od�U�a�)�����i��y��8UK*&ib�0](g#����Y�kV/Y��3j����TL��ø3TH[�/����N�ݲ�X�)]�;pɥ�σ���+��^��퉣c�BR9��&�x
��i���g3kp����%����;g27S�s�ʱ3�6�;��J�/l�M����Z�\�]i�z�p���V��UN�J�U8uC'6US�0)�m�h��a�;T��yj/VXm帻q��J1և.3gX�.3F�+^�4���wn�T����C9�p�d-4��uh��Rr�m]텰b�-����(�ڶ�%gu�>��r�L�U�ùfCY��Uͽ&���v�
<^:�1����w�N��Sx�fe�"�"�2�)W=�\�Ҕ��;�3'û�M��[�v��TɆV���IӃ�����I{ά��d��3��ܙ��]'a��)VV�tr4Ѳ�)�B�#d�S3O6	(��׷X�N�^�aƒ��lq7���5v�1&lu��������������h.�)[���n���u���o(NYH���އv���N��ֱ�$cř[f �(m:lQߒjB+�"Ѡ�S�R�o����U���:J-w�A�,�>#80Hd�L)c�pT�j<��m��f�nj�Ԡ��5AjU���kA�7�����{�Q�GN8,ŵ�X�8��n��q[m8鄁I-75���`EE�-�A�F����V�m��a�v���nU��/(���qC1�IH��m��I-�m��A"	��fg9�s��8NݴmEzӊ4��O^�V��m���ǭ4�o]���ӧ��ڎ�+����;zt��M'j�vt���_���o�m^��Ul�o�z��q��:x���vǬx��4��m�m�i;V�;T�[+�6���v�ۇM=ti�l+��٧O];q�j�ںi](�4�N�+iӦ�(b�t�S�em��m�8�鶚V�b��M���x��iUM�x��U�J��z�Ѵ�֞�6�Ɲ6�j�fݫ��v�M4i�|��i���6�����N��m���b�T�]4��z�M=c�N�c=W���+h�;4SM���t�n;l��'�z�v�ƛvѳ��+j�t����m#Jڴ��<m�֞4�ۧ�Zm]�v۷z�J��O�m۶�UT�=v�:v�ǎ�U�cN��gjc�=t��+�Hںv�8���W��+�Hӷ��t�4�
x��ۦ��GM�WJt��\tۥcO;i�a b+�7dCG���$�E�Hr�"���p$���HZ�!	Q΢�ܵ1x3���.�Q˄|!�U�M{J �ìxj���%��ރD�,�ʓq6�S�!.��$/��
G���H���
/|��IP����*�:`�{��:
��ܶ�,�&ê+��R�e����eCp���uW/�#�(-��� w�D�a- ����-��X��$>RAF�Ĥ��)�fָ�� ^͆�y2l�m]�b��+�QUFȋ�|f��鍓��A~�b�&qH��!
J�h�a��q0�.���Ȅ���RH����~u��z��R@=�����_��>�?>�ߧ�P�����,X�2kB���e� �k��H��\z��P���D�Pm*�658�52�T�Xot�џudk�,�|m�ǣ�
��F��;G���܃Y2��u�n�%��M�)��&*�Zn�a��N붒7��j*��A�%���������/m#[5�3���p�S�mՍ��uE��40q�M�T���2�%X�bT�ƍڭAJP�z���F��4/28j�Е^s�3�#R�oS��)W4n�W
�wC��
���կx�$⍔���F�e*�k.qR(ڭGk���V+<��D-�+.�i-��]�T��s�!����4�`����3�W\�D��W:�����7k�8��u�b��ل�w�Χ��+���r��:��@A�+i��lRG58�學�DLؕ��Y���5;ID����W���=�I�9�T�݅[e�Օ5��i-�:˭�Be������mЮ-�+�ݥCB�M�b$���M��;����q�v���f2�a:�f7j�r����6(�pݼ��}��fS�8a�0gd*Ӹ�l �44zp�Çg8tp�Ç�8p��Ç8vp�ÇG8p��Ç�8p�ã�8vpp�Ç8p��Ç8r=��B�6.�j�#fVm��1�ۢ��r�eU�M�P�R�Y����j..��J�|E��v^(Y�������q�£�J��5��0�<�������vQ�6&E=i���[MP�3�"U��`�������{:�^j�G ��ޕs�p�4:�X^Q�l\e��s3�w�j�"�eZ�v��DW"��޷��J�#�l�J�V�e�6����BS�Ң��Evw|�&	9�x��
mq�Kw-L��{\����|C�ۙ:�#^�u�[�Br]Ϊ۬ʔb�A��V(d
�jv�í�0�(�sr����x:��΂�B��W]P�;Ώ���RjH��v�A��/�y���iY��^<B���FLt4�K�&�n�����s�ֻ4&�o�&f���e�5�U�%��A��2�]�Q̷�i=�7	1٠�Tj����^.W���7nr�9X`$���8Y	QU�/U.�E�`a7A1ݘ��$�7D#��U��a�iN�����"ΣA�U�]`B���6��Q܄[j�j�"�B��@95B\!'e�G�8�y5l�CfX�a��QH��1�G
��F�]8�x��p�"3�����//f�g�ᪧKX��@pѣG8p��Ç�8p�Ç8l�Ç8xp��g8p��Ç8p�ã�8vpp�Ç8p��Ç8j�F!���2��͗��ޭba�lf��\�A�dkP��jfC+jV�yݺ�1���5ۚn7Wp.=�ĜX���:�D�5oP���ʔ���ޡ�*����\�W@٥R]�ee�X�f�ht&�eC��y��y��rݒ2k�O�w�iuA��K�7VQ=��2&�����]c��_�z�����<�A���� �8�2�� e�P2��)��W�6�m�FM�=�7�V)g�ꠏ�Wk)�9��F�C!e�;Y�@�hbH�PH����D��0(���yTQKkkV's�W��B���	C�[�<�X�<\�7pՀm6����DB'!���l��y�#2�Da1�	�	��"�(�B��j��N@�+�?{��X8(�@�Ll(c;(	h<����2��2!A/>G�5 ��5�F$-S���
�<�r�^[�m{-��͠���{�p"	8��؅�?C�Y�����s��9b�[�u�H�;�B�"��A+<���
 Um�!��Xv���^�
77�F��R�=�#o��du�;[�{����|�5[{	��D�1j,; �N*����._�P�X�;���@�s����5��u���Cu��{(�p3�P���n����=�=�=��(��20U��C,1��ym� w��&\���4�Ä4�U03_ibP�@z�����¯��Hz���xp>�O���p6���ۻ�n@.��DWS�1�<�����zm�]�:��,��^DW!q�<H���̈�f�@��GPb~�B�����X�y �U�Q��Y~�v�c��ً�ؓe*��7��Ç�4hÇ8p���G8p�Ç�8p�Ç=8p�Ç8p��Æ�8p�ó�:8p�8p�Æ8S�8c�ۿ|��U��M $f�u��<�~C��8���6�>\��a��B��m�\SXF�`t�!��=pk�hDA������:�p=�X�x��#�c��cI;1�ю�cMl�{cص��F��0gO]�V������1��Wt�1�6��`X��lq�b0k�͹���� �/tH�����u����+�_�nс#c�[��u�.���3�Q��j�A��*�t��J�ݏVu�������29��B��E�4�����b��"��f`�����f�@em��`������Z�A�/��N�7wz�%q+��g{����E�|�Ч���"T��S]R�ł6�����Q@� ��5K.�u1��ip�qD; :�(����N�i_h�<��[H�s8�w�i�U�Wb6�v�ƍg]=a�E�z�F�}:��B9f����X)r�
�^<s�mINƗ�ŧ��e���s�j�-�-�����������-6rP}2{���)ZF�C/]��������^M|Đn1X�����m[�L₈ӴshI�+1�`�2v/�P:��l�ǧ�׫�����.��WX�kE;f�G�e�ɳE��]�̨�u�Q��(�J��چ�_hb��:�+�3m�6
���v��v|j�*v�f֬���UT+�t���V��é��/dUXF�Q/E�]XeI�t��1��eSQu4���8�@a�F�8p�Çp�8p�Ç8S�8p�Æ)Ç8p��Æ�8p�ó�:8p�8p�Æ8p�Ç���FE�jg������{��V�̞-���.^�]f��x���a��tF�Г!9�x������\��j7�Y��jRKRŐ(�������Ai�MH=7t%ߍ:Ty]i���;��X���f�w��uCwϬ#��-:�Y��z�뭽T�s\y(��o�� ʱ�"жT<��$�v���b�qRc�7��V,i�*��N����4#�ۯr�{|�K:���#�3$�Z��!�azA�[T`[��p�ӵI���>ڮ��yU��ݩ�*I6�݉p-��4��6�-A�fJ$�A�}���UU7����Yմ�\c�̽BR��G�+��N�8.ǳ����z���Ave6MrۚW`�	+N�W[.wFN�9�Nm���K{)��m7��0e6���:uXF���`(ۣ��Τ+cyIU��d�ܕ���R�\�n:���(�Ê媺�k���m5]Ȃq�<4�bj��xJZP���˛K4$�a��v�z�fE�<"�c�KoE^1�mT���;A����=H��W�)]�8�{r�1�~c6�����0&q�����kH�xo���i:��N�u�E���0Ɂ��'г6����R�f�؝jN�2>��2�����tzp����F�p�Ç8pp�Ç8p��Ç8p�Ç8p�Ç8S�8p��Ç�8p᳇8p��Æ��8�yk���ØE�,HT'd�y�y�N�(,�[2�4�q���Q�`�О]��ʘo���9�<}�,�Ɲ�k$��5+诶�nպ���H՝CU#�b��r���D��;�����X���ݴ���=�}���wu� -F�s��Pn����l5�
��^��Zhf@���-9R��1=������V�c*q){4C�BUc,a�ݭ���F���P�k�3���kt9�Y0�X�S#�c(n�*�q��7VC�8�Fd�Ĉ��)��0iۻʻ�O/��l^t�U�I،!uo�Q��Hhx]����ɑ�v��5�W.�y�_eV�.���ί��n�lWJ쾩��A��Ҫ�o+ywda�=7m��[��}���`F�`i��ke F��0L�էԘ5�g���^v\8Z��"zΛ�5˄�q�Z��Ѕٙݾs;��o�T��-��7
	WM�g;J�����DmQN��uԕ��������{���8ŞQ��u%����Uz:{p���yݮ���oc����K���NI�,�n��g(M��B{�z����2�㷵]�\\�:���w��7C��j��+���sGr��v�C�HyPd^�:�:�g
a�g
zp٣F8p�Ç8p�Ç8pp�Ç8p��Ç8p�Ç8p��Ç8p�ÇG8p���`0�4�ծ"��bp�)�hI���
6��ǕM�/���xFZr*�@�UF�n���/wRۊ�����Z���8eN�;���b۳��f����T��z�ks/��S[E�u�T/�P�Rt�Ͷ���i;W[���`�q��Ne��^����mB/;p�-�����Xt�ˠ���UY��4-吖�����eVIQ�v��nnс��lY�-1����Z¬ԡ�&��j+]I���y60��f�%�)L���zA��%��[H��L�p埪�k�W}6"�5�8.N���`��m֭���$XH{�0�n<�W��Ûּ1+��;Z��&O)'�Z�3q�iѬu���\{�}�y��U�2�f{Z��_#�;3�8ȔY�ѾMJNX��\a��a4Bޒ��7o��dJ۾e�	���=�Fn�9%	���V��FS�
Qa"�n*��0��o���ذ�Lw������"�����u����{ �;��焺w���*���ӓq�Ǩ_��V�N���IY��T�b�y�J�+���I("id�$k왵�R�/�c�Ԗ�-D*�ZF�5ٝU�f~��n���ۀ��HF�-ʓ�n���F�K��PvS/�\�غ.w[��	��V�|�5߳��w]���<=4zl٣�8p�Ç�Ç8pÇ
p�Ç8aÅ8p�Ç0��Ç8xp��g8p��Ç8p�ã���UlJ(�ƋtY�$v��M��f���U}Ε3���ޝqU��<���+����GN,I�,{-�Ή\�穘����B��R�\�Q��)E�ܛG;*��"d�p�K�z�)���)@����<����u�걢ԖmeZ2 �&�B0�c��q��({��bĈ��(��W�d�!3O]�f�E�x�+���D��Z�Z�����̰�.Dg�K�c�.�S�z��nS-,���7*��"�ךV���S���2j�\��ݭ�o>��]�Y��	��Mk���ш�5�.���wh3i�{%9%�:�$�^!HE��B�nm�3�	`�Z��D�p��t93n��S��Q��������Ux�!�	�+�yX�Z�Gwr&�wXq<�{����YTv��q�M��"z�(fd��;R��9�;���Ս�cX�ry�A=֎w�ܧ�E75��}����.ox'�-�e�ƞ<n�Q5�c|Bŧ#]&���sNl���V3Y�|h��FDΐ�wI�9�lf8niͼӲwQ�Jճ%W+�4����NQ����d��.�V;��2��Y��
<��S�|�ͪ�����$���̩Gb�	^n���e�Cr �oK�ِ]|����X���4h��Ç8p�Ç8p�Ç8p�Ç8xp��G8p��Ӈ8p�Ç8a��8p��Ç�8p�Çg�{���jb1ĩd\Bj�T�MY�m�rДo]���)VE�Nv��ĥ\@C���X��d�y��mY>�9��D��)^e\dB����%.ʖ�5��-v]X��@�5yzR�@���-
(��<�۝��ZM,�v��'H�:�L��)�-��=��.n ��A{�� �T+8�
�b�2�
���	N>}z�Tbf{Jٕ\;�<Ź�<��a��&n�ݢ,S02�e͖���YT8oK#VI����]��óJ�U��M)[��D�7����)U�U�4i���؆$"����r����/uX8��L9f��b�!Ȝ��SH��[PE�Q���B%�0!-�M���3��UP�fh�6�	��j�z�*IctR��\z�����viĦ9�5eo]��Z&���m��~Di�L���L�MC��(o���%ﯻo#�W�ƌ�e��T��[9Q�{
)igd�v=9�)�Re��|�=��cc2����1�ٓlټ���6ҿ*-��nf���ʰt�˩N�Stƴ�
Z�N�Ǧ�I�컚H�b���U��h"]�ғ��T�,�DRr�iW	��GuO(������D�F87��:;��;�2ܾ�����+e<u,���Ի�/����/w��$�❝[�q���rޘ��/1��K�/D��b��9��Tv�+CCp�����̱�\�i�zR��C�����k6��fӴ�S%��Yh�6TXۦa��C�z Y|a)�3m�#Æ�CțtY�v'�U�oӷ �x�����:,O9rΠ�U.�od�z�d���oq'1]�v�vҧ�F��^�� �����p�:1�b�n���n�ܐ�M
F�-�I�>c\������Q�ܕUP�U���ƻ�Q��2A�9�\b��ȉ��9Z����Z�ov]�}Y��cK�Ы'U�l	�EX����	����M��f�Vऑϫq�L�G3b$��Y��yv	d�|��G^Y��T�(aӆ�4�{�T��)��e;����[9��i�N��$$�4��eC��[�����yp��.�l��9�s�;	�gK�1�'Fԑ�R&N?1n/!�5�[M
�B�%]@ɔY[�/�/k�1h�;"�e���٢��)�2dɥ�u���v��1DB�N��*�BD(V7b��t:�]���r�������a�If�חb�?M%P�X�7r���{ױu]��{ݟ���� I'��������l8�����'��~�uz���iz�ۺ��,3�����-@��cL��2JMY���t��!B�/�( %�JVq�����;CU&e)!f��j4��R)ҁj����ͫ���j���Q���n�p"��n�r�^�Q�c��ㅾ�:�t��1U�;{M�-�1e۴�Y�3�KG"�η�u�V�&����k5^�rY�^AZ3����di���+�Ĳ��_�kR�4v��(��vu頽�I�{5�;���7UB��j���̧Y�HdĴ:�gt>+���oD��rV���\c1]z�:ᾲ��V��j�xj��֑Z��(we��A(F�鲮ʈ�q,�6�8������#"-k�6�h�� u�N��9����}��je:-AYX���/�-YK4��:]�:��i�*��Ձm����ڎ�iӳrPa����N�8$�7Y9{���:�I�s���T�[�&o(7�+�t��^Ǆ�Z�Ptɓm���*e�����Q1�&�7{��u}9B���^J�N�uN�)�@Z�ɝi%"g'e�V�fQj���1�%�e4��� �Ifiy�@ȫnf�	�i�Z�8I�FqLc����Ƨ㻗n`;(V'�G1��p���1bc��>{��
�'c2�m`N:�3�r��ಗ#fyT�3���U_;��T��*��{1;MF������S4�����[mҼmD�:�m��H��(
%�l�Lmъ�j��M�t�U]��]�W�:m�O:m[+GN��v�qۧm:i�㦕�M�M6�ۦ�tکZV�t�M��Ӷ�l�OZiڻ+N�:N��n޴�ښUv�m�tҫj��EiѶ�xۧm+Ot���Jm���f+n4ӥz�zǍ;i�M��t�JmN��]��H
@"�0B"���&-Ga���R��Lv�1�ur���$�uwBQd66��'r@����/�=	��R�D)3�Em6��Tn��$����W}Q�Hey(��wMj9�6���EB�$�����GwT[l���j���VN�;==<8a�O*خ��7�k�^������b��jȵ��Ou�8a�g�g8����_4��SU���MRK���\�/K�$I%S���'u�%��r��$�U�K-��,TZeIlX���*����*�(���ڹ=ut�+�h��(�-lY�����[%b-QEh�
�H��EKV����g�8q#ڑj�j,Q-"���X�^:�|U�R\�먢,IfY��t�(�J����RRWwE")�|]$[�uM����WD�7����I2�wIL��(�U�;�KU+Mp᳣�Æ<����-*UjX�e':I�H��&��׾����R�*I�M��v��i��U���+�����Np���jiE]T��m�R��k��^��*k�n��^7M��%xk��E.o-�X�oKf��GG���Hyc�{�|n�������&��������������x�x��ۥ���eS�u��Ç�O�-��Tw{����b�*wcm�w-����t����id���*:,���wGj��wi�Æ=8y'Vyd�X��V4ֻ��%��L�rƄ7��7��J�<���m�-�k�]��Kox���Uޝ�ȶ-�������FA#�Xm�&�-�hB}"��֦�V���+fA�2�64j�S+\��������X�Z�
�y;cp��t���N�Һt��<tڻi�M����6WJt�z֦�iD$,9>2IQ(i�qB��A(/2��  ?��f��χf�{���
Kډs�Sw[��.�����X��4y\|�/���s�[}�����cz�s���2�V�+�ˬ
�f9��:�o����w={�V�ӻm����o9�,���kl�v�(�3% iH���{�+2�I���08��� �5ky
ڋq:ܴe�p8�ip�e�vD���6���r[���#���'m�}�f1�	�k{�_n���6�m`X�9o u\e/7Q[=?>��g-��s�� ����X�@5�����ɛ��nl�����P�r��/rW�_ �Ŋ�Q`P�Wّ��kc�<��� |~��+L�J��U�V3�[��R��Ĺ{ٝu��,������(Q���s/�U�UA�4�kE�fVc|�6�j����#Ϗ�Z�g��K.�Ȍȫہ��4[��^����iw�j[�&�ݦD 1's�߄�۫��@��W`֥5���ս"H�����75n)�_]`u�!*J��U���hur^S�l[�������zvgv{=r�B<��	��G��N=�\m��օ��M�����Io&����z�A��/���fȆ�'y]�n�
;�i'o T�H��Į��=�r�r"�ٌw#dGD��\����]�yG�wq�`LnA]� o+�;00�Ά�H�d���j�m��
�4�s仧�̎[���M���>�޺Ƙ��wl�wd܃�9�H<;���n%8!�D*��뫼U�sX"�h�?Rj��\lwa�*@L��g݀�����T���- �Z�-��R�9��>�7��}�j��&������^� �n��@]f3Ҕ��t'�fD�-�U�^#�>�NF"��[��3��{��{�S�P�=�H�?w �@sJ�uRq�Ɲ���$R���\~�ٗn>�~̸��}�����ݚͣe���bd�*�@�����rѭ�9��=SJ��fT^4����	VU��i��h��z����nص��UP��W�e�uq��C+5Pp��0t�$��­��Z7Js����p��tʽ�ZXq��1[��+l�zx5!��3RwHUB{*[�����ҷ��	�U�Y��7�7�K#���rҮ(C�'C|��W1ĹV�ŵ�-�q��IX+��(:��E��bx�����ŝE�8��������N�W]H8ݮޯ���y�G�7m]w#��m�2'��q��D��Ӭ�V�Cu�0][�7_b�����m��{p=7�B����$	30�����q�lY�P�S0灁���j8�')G!�&��O�d5�CZ�p#��)۰�?mAQXzh�Q�V����d����ϵ��4 �������N�+l1���#7z��ݕ/��[�(�Ȓ#�Gr+$* ��0�ˆ�������H�M
|����^�"�"Q�R{(G���)p%�P��B���o��QS��R`�o��N�볧���������Q��o�i*	\�)��"zF��+uj1[��UB���eJ܋Ԇ<j���dі�r7���y�r��Y?m��OG4XB�^�åM�ӏ�)�W�c7�$����T��#h�ӉJ%d�[�6�]���޷N������w;�I��|A���	�-�Yϋ�Y|�b�O&�F�����0V��V�p����y�x���]j{9����� ��e� � pnA}��i��e.�s;;������=8��:�]٘�S��HL�V�v�e���a�ٮEʥ�����lQdq����O�-��������z�2r�h+��Iܭ�J8[5%>��n~H@D!�wi�K����_u�ǷU��K�����j�QO�]G��	�b�Z� �|�5}2j�LDM���7oi>��D�'�֞�x+�zTA�?9��\��>���٥�@�]E��n��\�+�; >\���o"���,$<o�N�n]�N2]J�D�"$����F�<���(}�������:��F�]�r6���n�[�����S=�u�}�5���� ۫_&�t^��6L�۝��t�ۖ��c{h�Z:���\_^�:Қ�b��n�si�	0A�̭��o�������)���e��k(�7�T*��P|��m�5}V�E������2����e�ڒ�zU�f��ku� ���P��|����-�-��{�X�B	6�2`����H��50ű������42ɋ�v10��G���B0�_H�:c� �5%b���z0�����if�K��w�ev��.�;���=��{��7C�2��D��M�gfO'�!�P�%��tgP����C$䘹�ږ�L�<O"�-�uT�k�̊���i�i�/oA9)ظe�ź��㬋/{��G�������`G�����V�6��"6T��s���^��?a/��8�����WMv,骶��{�ހ��^
*����R�L5���$[�#C^������e�1w�qp6��mweDPo�_����CL�P���* q6�����ɫ�q2Q�x�n�*W}guro���"���c�Jv��6��˙��q�]��u⓶	�KF[�6T��3�Elp������x��%�{��;B{5'�>���C�)�uS/n�>[/�(,B?r|N�}t��}�e��ї��0��%��2i�ܥd%z�qu-T
X���C��j�Gb�*��Ec���ke�;0>zi����@w�:G��<N�;������!��9ӥQ��J3�(��q�0|�9�����+�Wp��ح�u�u�1�/�4]�@�����vťwF��|/������82�y�s˩�d9��۪��M�ᬋ�5<��T���4'U��m���j��<Oz�=q�v����I��N����A�	����}_��?c [��Y�g�J;W<9����3���j�>�ȁC��߮o>�SN��+��9��]s�i�߇H̽;�`�CG�GM{���w��d�
v����|�:;]�E}����z�M��#��r�k��_:K����B%;�.rB	=_v���t�Ҡ��u3 
�j�����8
C.1�wB짃P������r�!
�c���a��X�7��n��t�oUSf*[�Y�����mR/6���̵CũfT�yrۡb����"�V4f�F�sF�t���+Sq���[�cw�=[�HpX�ɢ�!S5�3*�w2v8 K/��&��-�J�O'�*�:.@�ֶO�59��t�u9�e^�@�G=���|���Hl����ol�n#�� �s\�Y*E��ݙG�]�G�|,��4i�o���{�[��Ā�a<�e���_���T؜��yWq�;�k_*��.부NP��x��#�Qu��o܊�Lt�b�0F=�l�î:~|����RM��HW����wsJ>�z-{�}��������C��*�wwԸ[��r�����}Qk�knA��[�t_�F{ �i�6:��fBY�O{�ek�7ݝ����f��~�>�����T����M)�z��&&��D%?=)_^k�gZ�6��`��B��rje^�������?O���p�}g�)a�+s��C���w�]�1w�Gv�"��9��T�f��mM���凱ͷ�=��q�[)HthE��u�\٭�T���Gv��	��(��Fs늢uU	DcdDl�vs1�e�%��V�7�QDPzufڥ��ڛޅΕuY��®�^;�>�O����[?*�����`^?����e]9������LR�w9��}���3�B�FU�&��'E0���⒊L���8��I�#o�P���Dhu�E,��Q��b�d^�A�f�Z�t_�xX��_q�9ds �4hA]��`X	C�*wCs��6��\�t�n���~@�;��v2�+�A���M�x���-c��V�)qP~ź�,������C5�)�|������6�xG8�x���3���k�Y��@oN����:��o&�8J6 )���D5�]o��J�2��{��߂��ke�����Ӄ��T�����������f�k�M�3�����e�O��tiʊ9��������nWۥp���`��������@ѡ��5�z~�1���Dn��oRbj˧�e3�Z�o�݂�t��Y+|���ŉ�4^��݆�wlT5G6�=���T��u)�)*W�� �8�@@؉�e�`kU���Z�S+�����M��kf9�x`�Op�m�9��V�[�{+It{w�g� �&LO�A*"��^���m�A ��@� �P���DB���Gvr�/9�����L�E�UiN&{�E�ɃT{1>=��a�!_m.��!�� S_���hp͔s.����1��u��D�/ u�������}c�-����PI�#�Ix_}ϡ.9����	�������[Ϸ/`{R(@L����hC#�5�r��G;�n�8�De��؀ ]�u���(��i�{�����jw��v!XC]M������-��0�W���36��^k��\��,�@������Eg�au�S�.��\���g/��P���9���b�x����N����w ��Ò�i�ӌyc� �sc�����h���6'���y�꜉�@��_@(&�cy4��%�fL�ݾs�Ҽv��m��eOL� �TO����=5��[Κ̓	]-���~��j�_I�)s�*z,\nƮr�A�;sD��2��*^bKr��Vu�Vwؘ�\����D��Њ�lh�L/�-kx���:�D�����L�T�ث��o5�j.i$U�6�&���Kre���-�ٶ����e֖�H=����,��;�}�4�0`X9�<�oX���'yO��aF2�X`�����g��rT���[��7X)I�#$�ʻ ��;Ѻp�v��!�!'q��3T=\��� ѡ܀��9��r�`�UT���vVoW8}�~�չyD�� �{����P��}�m<�wX#)򾶛�$r�L���.>�x\_�ܙAU��b�;�Vu��,n�ǩ�iI��*���'ܾ&�&��d��(��+�.���TM���3�	��pº���Q�]�9�t���y�U�_��� :9X��\����q�^��l�3=@h�E��+�g̠����޾���'�mZ�7ڱ� �w��]Ƈ1t��bHN,A�q�3{|\��'���Z����������;�\�9�f2y�4�q�<}��D����]93$/W��,g�?K��\��-����(�M���t���Bn%)���F��9��J���^��i=ӑ�f���cگb�zF��_�RAn˭ugfո�U,[��4������G;����gM���˻9��V7��3�L�6%�DZoT�lĪ��2N�y�2c��J��k�f�Mwt�Z[����&U�\����M�p�����nf���la�����ֲ�a����"�A'6倖�4ٚ;SZqU�U<6�s���J�vj$i��n,�u��U�WD`�"������43�Ӆ�c��Ov��wj�^dX�����i�	:����7}���:�c�bYX���-}eS�������u�b�d>l]^�<go*��OV��[M$4�M�P�j��%F�y*�,yZ*�Į�Ғڬ�e3��u'�L*��a?��)ۭz҉H��^�v�YF����n�8�����$9��+^�:�&�=Oq���yH�r�w��ċSmʱ��@�m��my�U�x������,]�6�rݚ̈���Q�wVUeC�a�R�ѓ�h-�����|�dfٜ36r���=�{~M)�c�rAɨi1YXg)��l$id�rS��Gf_Q�IZy�i�ō��l
0�y���?X��
X,A���%�6/(
��g������-�"��!���y�-�0Y@�w��Xb �����F��d`��(SW���C�6ޭ�t�F�{:��J�[�}���y���b#��[�d�Zv���L�����"U��*��7fVsܧW��V��L�(�ɹM���`&X���L���o�_i��Xz���w��;��z�i5�L')D�/��'x��)�^[�sY��]V)lX:eo�:��� �Y��fɸrSv�a23&��$^I)�����e��M]fө
*�{3XvM6iL�8��3��-��;%ӂ���HW�T��tŎzjv*Z�V2�D�i�=�����	�\��Y�Ӻ���PUR�>�bu��P��v�-(u����2���ۗM����-�;�h��U�+y��Q�;{�&�:[Q����aZ���ɥ'�q&�1�V�N�5(K�O�]��q��3̥�k���#8��iu�R��U�q��u>�+nl���P�	F����b���aao�I�)eD�{��.�0�f�
�\ڏ:������e�.���M�Ai0vv�q�ə(����HM1���m�_i���sb�ա��+��SNZ��1�:�^;��d�v���)�M�WRe������:�m�,H�Ea,h#�P�K]��`��?�x}����׶�7*�эQ�ت5�Kֵd[#�M��>8p��V�.Z���2Ƌ�܍�oծQFѱ����k�{�����ǏV#u9YQl�g�^>usnU�,Tk*���ώ;<<>>8y,"�,=Y՝u��<�<�'V:�Tj�\8a���p��9=ձi����5&�:�ÇGg�L8x��v&�yE�=,�RO��wJ�T������=>>=$����7bMX5�{dO�#(�>==<0���;�j���~h1d��M�հ�[!��l���8d<�&�GvY2��=��탔e!i�vd9dn����%�����s����B��G(eEl�3��H��.h�BqYD�����&�+JМB�M�҂�����1���e�4O�� y�=��7h�%ᘿr�|>�Ϡ�ZŔ/
K�]�Ǿ��_�f>�**+��Q �x!�v���ǁ;Vw��>�!��no����F37�}���nAȑ�BBG�k�z�}�s��锳�<]��9��[��@}n �,���]��!�?�� Eŷ|u�>�k��gnÒ=>�������wT��S.|wp���;���
h/ÿ],^��� @ �Z���oG�ӟ�����O���1�w����qf���	�fn}bT/qɋ�p�|������0̈�P�!.�`gE��C�5~�=݊U�y������̛Ãs|;2i�x,�ٖ�?H� �_��4�C��4��3v~�<O�4-d�3,����IY�i��z>��LN��^9c��i�`;
m��1�-(�p�����>����;Ś`�#�������>����6��u�������q���Փl5���3�����3v����hi`�K{�{���6���WHf�Pmj��RO��r{���7�4��L���<4�	�=�z;:G�������0�����������wO�9�vX�u�-�>��cco�q�鴥ֺu�7��i�;�EP�����z#+bL�vbԙ��������T�=K9S�&C�1޷܆g����d�Dbe�T���W����9[&�T��X�>��1��M;�g�#�u8ަH�S\9��lq=2�����n��y����?9��|j��9u��ag����^��g��~A���:dͲ��HJK�!�#�1���j}�������ױ��P_;"?�j��b�O�^�y��
w#I_0�o:o���*�7�K��nO^9��>�]���B%hׄ��
����~�+��֭	�{gx����r�z\|��ǯ�Do�'�=�#uy@������W?����e6-@��+U�EU���1��5K� �zB��B�W��J�Ԁ��NP�3@F��xV���n�6S��~��6!����̌��o�;O��F��7�.���{�^�~.��R��dx�ĩ���>���M4�e|�(��4&4���S��m��\oe<��*u�5�@���ȏ��)���~fj���#����#�s�����b���1�ꀶ(�`寥(p$	%%��4�;�й��z�������N�C<����ו#~wRg���Q߭��Ӆٯӊp��> w���VO�~!P�v�h�<u�AM���â�W��l�ڟ&���W(����&
����p�,�-B��J�O�WX�\�'n_>.�*
�Z(�x�X/m;w � �5g22A�&��눃�h!�`h�3���y��R��r|�5׬���������R]�sH.�a%�rt��;t�M���7��Y��Rw��,!��[���[���M(�5K�H��.s#�i�ջ��8h战P�o3�/���<%(*���1{N|l��l��`+v��)�quF$Z�vg�D����㋕雈`��۸=��^�!�q)͆�ED�5dl�w%�)�K�괔��̉�wt��w�0����e>;6S�l�۲$�֑���N�fI�<�skd���w����=��)�~��/�>Hb�<�C`5��5>8\������x�~)b����r�O�r�O��6���Je~�<�EJ�
���-j��#�q�{Q�%Bo)>Z�k���o6E��q��Z3
��zt��K8t�E���'�J�yK�n#ݏ�]jJf�p- �5Ĉ�)��G�.�y �fuM���?s��T��N���;9X�
����y鈉��b�j`}�y��%����7�T2�Ѧ��he>��O�$���M�-� ��Rb�5'`ܤ<kG�����}m{W�^�&��ZP�3W�'=S�J_Zh���\W��.�F ��C��@���}�oC����;A� �Z���*�S����ɨ�������VD��z�9����vfԣ�n�-c���C��lB!��m���5�1�"?:����<R��<	��	;��v�:�
���iL\���C�bR��Y#S��k�� �������@��{Xm��)��fo������~`��;%��-Y��˿�y�]"$J������E�]�5��3F��`�@��᤾9�ߥ�`�Wʺ5����ew���6�Nq����e�����u��?\�C�ˁ-|Q{�����	�|�nD�f���}��a]���Y�wڒ=���=
�F~�~L��`���ל!4H#��zk�P�r�(w�ۮ9��� �N����U\P�����IY�+6b���4!�?1�X�=�DKH���t��3�˳*v;yV��O�%��oj7�*�k*!�[�jy�o!�x �U]������[��u�lf@"\�����,��I���eQ���&�m,�h�teD
�����jE�63䦸�Rۊ0l蘛�M��<�a���'�;���%��xv�Um��g���oVDa]	�hr�G��t�܎�5gsN/5��.k=�T�q^�^�����Tsu+�K�h}��nj��n+Z��QM�wmgN��xe"��zo����/nc�X�x���]�xO.��˽�s@�%��fiؔ�VF<��Y�VNFN�{J�:m=r��N��n(Q��wJg�n�� p�g��О�M�E�I��o�����va���U���3��DdT�{��<��Ҏ�"��0,+Ս������ ~��R�֚5�4�ut�~=�HS�-�')���~w��,�ä'�aBf|sP�i����@���.˽*���w�$�H6|�������wC�S~���r����,�r�hE���]��;��q��8�c�O<4�Q��Ǿ�5;��]�h!�A��L�2:���4ST�B���XKQ!�A�L]E�	Ճ<�O7��uE�֟�)���`
{o`��{�͓Ǉf8�8=Fe'��\J��w2�y�	z��y�25���O^ʌc�����|����P=�܉� ��0~��f��@����E��� ���Z�@�"�֬J�������yH��C���Z*(b��*�\%�{��E��<��D��
��/� ���_~����X�q�[A���!4�����Y����5��y#�ӗ��vuB��@��. �������� �h���f��Z��
����yqvgނ͎��3��XE�s3CaD>�&�y�V�0p]�	���ܹ,{o؆�}�������}ؑ�;��A_��IЁ��,�Ƈ����0���0�ߍ:4Ax}�OiUbq2y�KwGWo�Zا$�X�V����k^;˝�v��wa���)*��0� �����赖�N]�u9���y�v�]S���"�]N=k3�:�j�[f�6�{V�k[v�Qt��Jմ�/]}����:>�*)f����7d�bj��we�j�T��]��޻�x_{����>j.��[�?�u�Z�.�@�¢��:����}uʓ-6*T�V^�4q���ҁL�B{a����t�[ E��16�j�<�@q=P�!\�#��>�7)�`���H����CV{��?�8�=f�Y!�'6�k�F 1	�&�(�sy�Zow�1u��5n�[fl���51��D��0m�����Օ�`��1vD.�S{�P_}'&+�>z��k�iwz�_9Ȳ\1�>:@A��zʢ�+X�	;�-mU�^n5������zy�/V�|�l7�O��44y�$�]��֒�.�ʱW��Fh��]S���"�L��VޜnNw���z�����	̋&�o�)*�~�G���>Ӧ�p���='�dN� @����`�V�]�G��|�u*��	��s��`��;�tr]�C�!�~������{����
p:�E����!���3c����NlK����t�uA��xP�����?i�GO՗<�e�����~����Dǆ���0v�sT���1���:�Z�M���C\����nO�O�d�N�jk>Φ����Ԝ��)C�R�3A�����U��/��r��ŒU���&�qQ�'h�;�������2n4�ɒ�[���.t1�
�Q�N����T�,5d�E�����M$R�4��[���=�-���ѣ���x�p̀I���>���*�Y�����t�xC��r}�C�RQ�s�h@�e�n�^�O�g.�?I$����wʁcv�Go�>��1FP��X�]�>�rvӋͬ�x�2��[�(i��e���`��x=1ށXNC��q}0��=���9�X�*y��o/ftB#r�F��O���
�i�!�?[�;�9B�T�	mœ�;m���J��5Ӷ ύ��8�c���=��Ċ�2z��#Y�=o%�߲��N��^����e�23��*��mE3�(e�`���q5�\��\�q���EZ�%�|D��b\����~�T�$h.뫘N.!\/}VpS�.E��p̎V2`�z�"�Kr�8�a|��^S�#˟���M#v4�]�g8�yw��O��ԡ��@z�&;�!]RGs�}n�ïm��3��$B�a#�4w��R�ި���R�@��.���V�0��x��{HmӒi�l7�&8�<���5 5��}ԧXH����+^9�0wT̪�.�9m�G���X�.�؜�gK�)콳.��W/Fas6	��Tp�	P=�2;QWF�@�YQ�7u�����lw�!ׂ�2a<\�����	�^KQ4ֺ;m�않�-�s)f�Z���-��ђ����ur��0O�{������މ��E�)dN�#E�ƍDIK�I4X�5d���Wߏ�=�k@^o��2�F8��Fk����6-?*�E��_)�%�kv(�c��|��4�r�m�b�ڌ���32}/bf5=	ye�1Y]�?�P,�+�%�j}�L��kG�5��Q��G(q�t��& 1��	ށ��@6[!��4�=���+5V��6frp?R�\/o�p�O�K�Y����M	������?�R,GF�Ի'�뵳��D�w������Y�d�E3������@G�e+��p���?Ø��|V{�a�8�����Dԇn������(	�3хE<oD��A��f�L<���o:���S;6��/M�َ1�"+��u�O��b�*S��/�2`8�}��O��o
���0�ay^���@:7�o������7S�q ��̘_�w���l��+ߣ�i2k�yʋ���3'����<�W������^r���%f��凜&���Ϯ��?zf��l��g�|O��W���.��fL1�ā|���Y�@7y��b�	�ED7
"> �BΑ�׏w�Dǽ�Ob=K��,LTSaʤ�wVVf�,��#�
oES�;<M��N��ܾ:���J56���A��4�ZV���%�oƔ޹�&s������Q�M�NUcʹ�HJ���=!pxn=����	reΓ,_�?�z�D���TCEBJP5d��e�CVHh������$n��F�I)U&�jI�yg��v-������<c�f9���b�gE6�+�a>J/��uqO�����l=m�vz���l�#�c��a����Y�'ˡv�E�
:�1:����6`ΦndJ89a�V������-~8���@���%�6V�F���Ӟt�`C��p�w�����Iu8V�g*�g��3e8��!��A�ǟ'�3�S�� �█�y<^�ƲXIr]цPa��뒼����	��f�tY�3��="��7�i����1>�"Z��3Ğ�oL(�ꃩj�vja70_ SƙC�3X����:r��q p���TAS��q���bVJ���%�B��3�3N3�$��>�`�c`cC�Hya'�}�v�f��<�K;t^�ϣ`cc��C�}�u{�͓��q4���o�9�"L�D��@;�3���y8�0c9ӦLq�D*2e��Pڲur�>6�DE��3NZPw�&3.�V��6��o�!\����ю͆}�^��#(3�ۡ���4�^�߲�_Dn�s1�Ҡ�_��Ǹ�_LX��T�Р��7�TbY��g<�XQ�Clu�"O'{���	.3����a�`#��T躜�Ζ3ҳ��Q�}�w��Z&,��6F���3�����*�vr����w�<m�Y�j�"I�$~K!�!��
X&�#vDl��F�e�-�6Y$�TIԭ\�h�n��r���l[ƛ[�h���ذi������a���C͸��σ�,�%La&3�'Et�ؚ�=�u�jb��{*%BY����̒��G��!�9�<oTH�=�G��s�	�B�j\��ྥ?R�� n�<���/�ܽ�@Θq~d<����3<OO3k֨�{��;�m��R�Y#������m��-����g�>�����7!fE1��ɴ�K&Vڦ�)����9SQaȏ:�3�:W��7�����?�yP�wR��6
��� x8�ů�}k�ˬ���Ң��)�hb��y�;n�h�+��W�����G�`����[p�2��6��2K�O�L`�T/h�lj�Lz�6�^���Q^�k�bj.��Pg�1z�=�:�h?j`������@bc�&�̤��:����앛��"�	�����4�q�$3k� ��".Q�0�Y3�k�,��-�&bg3T�R��� ���y�7��ѳ�D����>6����d��q����t߶� �)_ v�AP%��'�S�&LNF'�X3^�m�C2Y�F;p�7� {��/�_Q�}����7y��*�]3���S�\}�3Y�奵s��$��y D��N���O!LA�,�V��m�w+=[�Ke�.NӬ����Nmm��a.m��-���5�j[�A���;S�^Y�I��YE���Դ�j�L=[�AU\U�H��b�Ҕ�Ŝ��V��d;�sg��%���V˄��ғ���Z7-��uU9��uU���p=�Vɡ1CR��;j�5��e˻�9p��Y��u%�w{�V�Hv�Zy5p���űe�r��P��%��S7~扯�TS�[V��Ʒ4�2��v����܊��C0�-���Jˈ��n���gu6�TVz��%P9�d�30�=}�1Rʽ��v�,b��/by�k]�MA�h�n��w�`��]���˻��<�T��$;|���}�ʯT�~�����Uc�eiQ��M�b[s{.mKE�꺥��i����Q�(tzT�-gj�mHӌ'9��v�[y�j���M����K\�]29��KIqK��Vڧ%^oU��/��ܴ�U�:Y���"_c�oj�o<r�"�Yz�:����Kb��	��I1@��vC�P����f\D�iF[4�:��]����e�f�K:TllUP�y�:�Ǌ�C�VrQ7�e��%5�-�ņ��QLh��l,��z�T��:��+�%�a�k�X�<�G2v������C�k�%Y��z�� ��&,P%	C��<�2
z�
���%�;�C���n/A�0!�W�������(�B1���$����\Ɯ� ��P�Q��jf��n""���K8sz� �r�I5yZYRY�����V�nF���0�K9z��f�,�L���jtDIs��E4z6�%�6b]
Imb�\J]��M���@�Vq�8ӻ�V+)��ݶ�;kET�rS�W^�B�V8�\��hv�r���^���b�+1�����A�������ʺ4Ҽ���"	������lݽ=�:{(8�哕�'F�!�Z�ur�V��s��YW8X�u�OD�m�aV���O����T$�f�g�gV�f9��SG"����2IT���5E-�B����ް���Vf[�T�`��U��![�:|��K�	#|��8�x�iw�$��j�}ێ�4�iff���X6�i[�'�jwV�]�屖�M2��ejs/��1z[���P2M�fҥ�b��M�M(�&+D$`渼v�X�\�u��M�O�P��b�m�x�l�nZ�)��V�,�vC��:9㆕G�宼�9i-;w�ֳ6F.!�:��ُ�;a_B(�)�]��Q<���Q�F]���=�ܓ�p�|��_j?k�*t��E������q�$]�%���x�}\&���M�g�ؿ@�M�/��F�x�&��
�	
��Z�s+UE���<)E7��*�m>����u�\ݽ��t��a	 �	!�cF:q�
�駎�l��m�t��z�4��o;i��l�ݴ��c�i�׎�+���ǌW���s�63�hdpW1�Œ
����eU���kV�fs��3|��֗�~���vTxm}Z�Z��xU�^[�.o�vMXN�Kge<:>;0Ç���kTy�IT5d�Sʝ�*<�MQ�h�Ҝ:;;8zp�I�6��ڢ*�ۛ����Z�Z�'Qg
p������Ƭ�wR>���*Gv,��V]Yl�������Ǖ�Z:��E�vC� �]+�MQ�t�ޣ�8lᇧ�vޢձ�$�m&�ʒ؛�Tn��i:�ӫ$�M�<=0Ç�=��$<�&��ՑՑ8SG�8{#��'V[#��;����R5c�;�uQ�&�l���ÇFY��k_UsX�|���ky_Z�-Ϟ�6x���m˕c[��}�>�xxxZ~U������ >i��긴�r�y��kkq�Zĥ#N�1]���p��Nq+.��T�vĨsV�v���B�6^ެ����@�+�vi]�ٷm:t��Ɲ�v�@  m&�j�%"MF�X������d=�F�D)P�(��e$�ERȚ����#J��Ēy�w�x�뿹���z�G!B�I;��*_ا�1X��y�PT��Ӡ�s�z^W�>�Һ
���Z��5��=y�zd$Ͼ�`���t?5K���zO"4ȝ<ޖN2��!�G�^!<�r�0�d��^��S�m�xfBn2+̼��S/'f��dC3�b�Ձ@�uo�.<L�T5�L7���6�ڗ�<"�][��}�*�^�Xf�a�y�>�0T�|I��������-�U!�+vkn��7�s*,�4U�y�-���Z�L}��r�Ξ�������#[�_H�
5�3�������"[���ʬv�9{�`3�r�hב{����zb�cy�k��Gl|s�&+"�zǎ�7XӞ��@G�Μ��|>����0�^p@eCF�;O�@�,�GZ��O�Mü�3p�L�㜼xMڋ��i�ˊ�W]EoJ�EP����Q��N��t�΃��q�R%^yn�3J��[��/�?wwW~��m3A�*�K"G��w/@�p���x}�TC���4PK�+k:~o<X��l���L��%? �!��p۩#���2���/��;��q$	��EG'��P\� �$���A��`�%�f�ێ���ej��&#촫t7����v23�������tXa�7� �#pP�U�)��j&a�}6\�z���2�;W���U!�ݷR�v	8��dh�L�o���bl�x{d�������>�?%yRCE�!K)Q!Kn���݄.��4T�n�Z�#Z�j��?�~5��Z��7_w?�Z4��~������
�`̈i[��
?���@�S���Ս�t�i 68fCYz3(�˟p�����63�[��F�dTx�ɭ�`����4�a��[�%�Xf^�����'־P��SY�o>���2��T \�V�TƳ��A�S��2��`�Y�3e��v���q�e����x�dO���⺜)�%�GڪO��=:G��[,fp�*ﯯ��r��R�vt!��3C9�P�f�P2ޓI�
�o4^*^�<h@ay:��şq<�����ڮ�y��	�dn��?�"y��>��5�󯗅H��K�'�-����V�*/�Enp�XJ���T �QR5�yb�`�Ӑޑ�/�G�[�0�����2.�F�e�B}��8jbŗ���q�ZsڧZ�4�'�}BP�s@�5���Cʼ��d��n+�ҥ�0|>��EO@�
�}VI����#I�7Tb(\I{sQ�sZ�3ɨ5�u��x���;(�B�}ЭL\P����£'����êQ��L�F}��?e��qQ�k�y��ن�/ KQ
�Db�9JKÉGҽzo3w^������ �:��cPo"&қ&o�#�q����{�]UEj�h�(��h��@�lU��s�ڹ����f]f����Y��d6�Kr�����U�U����D�B��ը�����]���!��>�Ij$h��&�!��"�7�&�����I�Ă��!��<�RW��|�Ӽ?��� 6�0��=ސ��/�X�"F�傍	s�MF���P��{�]�S76zr��xzj�{��!#�;�3��>6i��0-7�sl�Y�� ���;�8�n��O���d���l^΂$I���~Ye��_T���0��>���ܬS���nj�>���v��@�k�;q�f�ob�;a��)�d�l�X�E��Ρ.A���>UV�/��{���<�����"�m푗��4;�TL�
8.���5d{�.\����b	 �mޝ�\'������.��ֻo;��%����M�9�%x��/@��%�:ĝn!b�:}~
���Nk��
C�N�]>�P0ɨ�4��d9P��f��1i�r~P�΍�ޡ8���@�������\���$ᚉ�?@�<ޑz��ߊ�O�('l�X{H�~4=����(tlD��@ř �H���ͩ���(�%m�O��<�鯷7R��u�q�P��@?-�S��� �f�C@t6An/��	�Rhuk���'C�D=jw}gm1հ_dTi�n����)�Y.p�1�;���Z�E�O!�*�[im	ſT�J���l�*�<7V���U��.�z�#MPbm��ob����Qת*�jQ�8�η����c�!�?~�߂�%*�:�I���7a)bM��R�#v �I��Ձ4RH�I$�{���w�����Ė*:?\o#N��0��7����_!�-�H���b�5�c��Ge?T��P���	T&I����}C�t�탯�g����ݲ��q�gSe��7H�͛£��^���܃lc	�L9P(OF'�Ʊ��썆���2#���.`�����@ceuw:���g`�C��y&�L�d��:҅@�zP�`�9� y�d�l��&�yj��<�ʛ6��{�:�&:�����\]����9
�M�:k1m����h��%kKk��=HX��<B�q3�aM(��`o?�1��:��P��B�k�(��7��!�y��`1��xlaqi�g2Ws����� ��ϖ�"}��s�y+/Q G����!���w�ee��������i1�����і���p���Iu���2D���ᶃ�q�k6�c7Ƈ�F�݈[���@?��~pF�N��g��&�{���91״�]w�H��*`-ol朽>h7�����{g?����Ǵ��F�?ߤ%�\9y�N��rd��&��m��m��3�C:[(���X���*�H�܎.��|�C]R��:i=Or�� �. ��`�ܩu\-D�X'������}cu���!i6���4���l^����E���L��*;V4W�bDˠ�T���n�(�繆N+j\4t������wʹ��̂~K$G�$�*BRȑ�$�A)H9bh�!�4T��Չ'�}ն�I��������@A ������<��1 ! Q�_�Y��\X�����W�"���@�l%�S�F�@xe�:������/��iw��n|#ҽ�7�i����T ��@�c@f�Za�6���Me��gd�;�Z�.p�Bȓ1��a�<���5�,,@�������d'�ϚС�����F�/o��ׇ�����"L�`/`KH��^\&MIY"��X�-���"C�d�5���PV�ʸ��v #/)����@�2=T5O0ʸ��C���=զ�1�%�����W[>���c�8L� �>�:d����z0/K�7a'h����x�ʐ�ɬ��	����wv||>5}�(�[���H%���#�?0�0-����p[1XvӐp�|��0�Mc����t!��8��Sj��P��Ȏ��l;9�=G�F<w�/��l���A�U��ǈ�[|��B*7`@���<�4:���g<� ؔb��!Dy|B`��5��D(���������,��W�S�U�z���S!|���9�~�.ɝ�@`e�t��R��� 
|��L�dׄ��U\������t�wO�B�9�am�0�V8�-ݫ4�ʙ�[YJ���	�:��9pʒ̋љ����ɚ��8vD;�'rq�GoS����L�8Z�!�����J���L����Il��`9wd�Pn������4R
XB�5R�w�g��_{ϴ������}i8��@~�
Q��l�8=�H�XӐ�<f�LC��ڦ-uRq+�rYt;���0�h� C�"# +��*)B#=U����,]��t)���)���3=���闶˖LC�nYt�������(|*��6-{�>��[�t���v*e;�8�u� �R�`V rGu^B粐ȹ���Y�A�,�9.=)�5=� 9�2a��	����-<�a�(�����x[n^�Z̡H�Ƭ�BǑ�?�/�u
�3VF���-���a����u�_6c��& S�~�
�t�7cLŽ�s���{h�ޒ���W�!�l�`x~"3gOLxЂ	�CZQA���a;0d>�T+�T�u+(��Cw�s@�M|v��q��{�o�̅:��;�l���@M����-����xF��zy���H�ƫɒ�s>y-��*o�w�;1���Z�&E�������@J#)=ת=�-�8�ay>�-��O4�*GeoA��\Rf8|"�|,`r'��� x/d_���G��z(,|}�%w��s��B���Yx��2\�ϋe�1�n�]�1*���}:�q;;V'���4�9ʂ��&�7&�)�ܵW���l��q�� �A����U�+�I��y�2(>}!��zI�V�+b�1�B�idE����Ť�,u\��lWv��|,
�H�����=��P�Xj�M5d�5a4R%,��DՑ'��!��R���&�ʎ��m8����ib��|o�A�<��|	aw�u���/���"���iB�mk˦\!��������3?�:xb�`z|�W�'�����9H���k ���!�Yo&���L��������r�K�t�lC9_?T��`X#6̑������I��r*����{g*�ߦ��3�|�� (͑��R@8�=3@�-٭�=w�٢	��4��jAL^Ko0Ow�ߌ1y H :+?�/�%�΋_p�(���̜���C�zܴw���<Ñ螊=+'P�s�2�	YƤe�}��a4�s�'@W�Eh���.�TQLel�c�h�͑�/�J^�����"f@-��>S�� �#>�ڜB�B�J�
���B��q�=Av���θ�%G�-$�Lp�"Zo��ͼ1[�5��U[{0fJq�3�틈dhD"�>b;�_`�W�����Sm��
����;��	Ȅ�/�r��<��i�]c�� `�h�-A�i�DHڔF`��>+$e�����r�F����D��<�0�%B�7uz�W#�l�s�ȹ���qJ}%��!̼Udl�
"}�mX4�ݰ�D�-8�U�d�P/�.���99)WW�39���Q r�S+��,�0��\�\l�Wm��Z�V�Y�Vi,�L�֜4��g.5�abu�dS�9l1�R�#oPG���BS}���h�)Rj���������Nu�}��y��w���o@��B�2��>`~"���1L��d<��s��01�ؼ����Q�I�1[�tnL`~Ң�ב�����yǦ߉�|c~�#Y������.~��~��b�n�}5ͽ���AYG�]�cF��;�����B2��ÀP��vt��I�RXG�{�|BJ�dT�8%����\web�n���.2�(ML
Z'�����L@e�dc�;z|ƃ~_�O�����I`�g?xu-C ��B<�N���U��1���@�W�� ��?�6A���������W �H���T"�C忔��roX�>��`��Yb�$t��2xˮ��nht����vWtW��N��p�3,'��L�/-m�{��6Ű�1����M�F�好 4(�m�by�Z΢A�(y��^S&	���_}PzQ�� u�Q{hY~�f�"�Y�}� ��C�A�1?�Ӌ����/���	���2���	��#��~�cF߯����Z(�j�=�_�D/�+]Pb~�#  �Y��1�O�0�o�9�&#UbFE}�?LɅ�r2|�Dl4�B�^_���,i��I�Ug�B��ICnu�w�LY�dͱkq��^��G�Xbj��
dU�?eXUz[y��4��VnӶ3�p�/��I��	��[s���w�}���<�B��b��|It��_��dJY"��]B�B�&�K�RIJC�Yj�x�s���;���CjƕU�M궺����D<H�5�`��y̟���?*�Bh��-Q�����6C��j^��H������ol��?�,]	_Tb�0���1i'�L�g���GhUS�&&�R���A����lƨ{Pl�N��"�<�m�&h������]x2���6�/�,P�� b3T�9w�R�Un�O�l=�]��'�� �����������
�� ���j7Vʓ��6Ě�;l16饁��q��/n��+duհƯs��v x��"E����'9�b���$DYR�[	Z�c�yc�c$��L�~��}X�>�Њ�����$������xf����oռ<�>�@�0��Hp2`�n�+)�:#���,��L<	������u_���|Zo�v���^vX_�	~e�2D�֜C�z�ޡ�L����b���X�-�Ì��Ӌ&]��؈q*��}=���x���C �L$.�OR���%O��ER��6�?O��
��������ZSk���vn���Ey�:Nh;	qh��� �)<�����T��A��dOr�C���`�ֆ�9�M�i]�2���G{7�k��Ќ��9Y��U+�Ke�Υ��u�D�O}�J���Ca	�@��6?O��ǡ8��!{�&vʹ*�+/q�<곪G�Jή�1I�z��`�R�jÜn��3�C	_� >Ѐ^������5Ԭ��-��Po#j�C�Ը�C�9U��-��!���yt���V���?A_�u[���kڤs.�Χ%
"&��;�i��7��L��O���A�D���G�k�d_<�]QWΔ�ٽ��z�ŝ��
~��D�����{��5���"Ί��.�y��A������;)C�Xk ����,����#�d?52>�J;`>��"�3���4�S����h�i�Gz�(��.v��uq����O��H8����ԉ��#�.x��`����*�"Z�.��1c0���^N<OXL:�p���/��8}A)��GQ�9E�D2#�(Ӎ��:౞�K�C�f5<�F���w��ϑp$~��~XB(nl}#Q_%0r@�ٰ{�A\��~Pf1Рτ�l�	a*J�M=���E��M=��8��}�����_p�F��48��O���*<O��4�mB����c>�3�u�K|� 3{b3[�À�c�w�X�2�����f�`̋��b�]�=3��@
��e(K��� ��I�ِ�� �u�PQ��ݑL��S��R7cl���E�q��x{��=ᛎI�q�=Z��ڗ;m��ۇe�:������T�ETR�n�,-�F`yݙ�lӚ��.I|�t��sz�Sqv�pl7;�7y yȃS7+�}�f۞W{$��&�+������8��N��G�Un�
���^�z�j��f&҇Xo�I-!O.�����]��UWeMe��[��7����V��jM��8��D.�S�����ʙ_J8�N��/�R��!B[��XD]UY�*6���ż�ID�:n�#�olL�PԮlU��(�Cɷ�OM�[G{Hj�K�D\&�^�Dc˳-�wqy�q��ڜ�bM�d�( ��Bv�ꁂ'sӗ��-8j\��-"�V���lenoe���];��kc�lkǓ.ӵ0\���B�������n�[7"�8�^�%���-W��n:�^^]��x�@�W��$[r��k�:�5[Lv�ыΔ�Ze�3M��B��pv�h���d�3�^��b��ʼ�&����[��e�psp�o��u���Աh��T�s\/�l{s[�ݸX���,3�ٕr��1e:�*T�AMd̓�;h���i̹�&Β[{����n�9"̱�r����r�ml�%�e�QS�d\Ӯ�y{
nV�ДOT���Iw���#G?� G}��Xu5;�6�:a��Zö5� �!�vS�(4ŉ��Hb���k��}��~<+����c�JC�H&��H?;���-��iM�Im\%z]��K͛��4�IB�&�'~X�,]�N�b�p��ʎ��8V�Um�K�_oK-��J���{�4���T���뢓v�6d�� �K��6�x�tPN�mU<���W9�\{����o��rd��N�Jt�P.�^i�Wiƭd���3V[bB��1����ǒ-3���vLR8U�A�Ό;�M
�]�t辕�6��7�h��ÖM,��S�g�`�_v�tk��k�7�
7��_[�����r�b�0,�x�^lʺ6�T��c��|��&s��]�$�MlP�/fVe��re(9�O5��T����Ў�NcQ3/V�٦�4{A�Eu�W+{����{L���2��/	�zJ�����\�5#e�Ӱ����;�-�Х1���me4���#�F�d]�/ZW�F�{�ut�T�*��\��n���i_QK%^K.��Jڀ��R����5n��^.7[�fIr�%:�#ٵ�W��∊I��Xp��lF��؃�Z��o7rV��Qr���,b;��wnd�b�*�Q'��fK�i�*ݙ��U��]�v�ՊmS� �+��ۻ����gm'�}�v��!�@B��y��mw�.yۭ;��;�;�}R=���ؖ�f�������Q�l&�Hʓ����:<8p�b{P�>�7{��&*mR{`wP����a�9mO.y�k�U$�H��)���g���*:�Xn�������h��Æ={gu#ꉪ��:��!j{N����Çg�E榨Z�&�{��{Rj���d�;�V�)���Ç=Hręby\���V��e6l��Çd����5"n�j��I��^��o�C��|G�=�EA}����W��b�H�k�#D�yf�ֻ�Y6�Ը�{�^���h�svFm4�ᨭ�"l��緜��9�<6ܷMo�O�H��KJT�e7�u6�R���{[_l����=2n���e�V��0kM&ŷ�\sz�2�iq<ڔ,p׊+�����Z����l��� EsøR@�$�r�#Nlx�D
g��}Y�,Jq �Nβ6�q���Ӵ2oSp���i/�脄�%�XZ�"-Ǚ���.3S�ϝ�û��t��nA�7�S���i���cy�%�_P��J(�����{�=�{E���|ס��"ò%��]�:�FYÂ�0�`��;yy-40�+~ˈQƆ� ���\��q��"�܅�#��7MŚ��i�Wg�ס�z?u#Ƅ�xcH|�\V�j�h.e9xÆ���""�R0����]5]����v�j��ɌHaYc�/���HA�$�Bs i+�H�#��B�[L^�M��j;:�4)A��&<#�Fȉ��@�����ր֡��Xڼ,��z$�"�Cr^�\���x&�Oz��V��ئ����a���$@�Q����J_\��Հd����M��Ź�f��s� ���'U�"w�rH�lh�ԟ�9_����Јq����`��\b�%�t���`�O���[9�����r�M=�9�a»,�!�*����Z��ʮ�Jmߊ����! ì`,��b4Un��Pz�k&�����F�vUx���W	�ԥm�e�3I*g>�;�AU�:Z�������y G�<+�5Φ��]JS��non�7A0�ֽ��"³@�X�2.V Ϯ�C��$f���GB�=� /b�EY zi�Z�K�����>ȉ���J<�ı7Ƶ��U勼[R&fr��G�In�f��B�U�~ú��;'���t�����y����YN�sw,o���l@��J�RQ�MP⮇�:0gQç�<��N�&D�q�i^�<�F���0<��rANy���d�J�7v%V��8�T��K;?c��}��si1Mp踶�K=�	JD�g��mz�����\������	Ü��gwG�U��!�Ҙؠ�3zV?7��`����������1�8��������SX�L��]��y����G�0��k^����;�D�z�g�+@��"#��vEw���l��K����u��"Z��w [�TPG4�ا����X�_e"��ǓQ�|k�'��3��Q��읞��=.n(p#�V(M�대���k��<gZI+� @W���i��ߗ�vj��"��Do��&���������UH�Ri�X
����ڲ�6���Y��|�!غ�cE_��#).���y�\Rܫ�J��q�2�M�~�Z����1Q$�gvLLp�^���j���;��C�ԇ����̝�Wʐ�h���2�WX��	+�ݭ-�sk�S�0� �Ҕ��w1[ܾ'9^�XCDpB4f��ߞ~���֭h����R�R� �� �7�������#BӷM��῏�/��a*L$N�~zB�O:����Բl&8��#�T6`.�S1���ܲw=�������Vb��V
"ch�A,~?0���5����^ʇl42}0P�Ԃj}|Q���C[�	��`!!�qO�.^�XP�A�;�@��3��EK;�!��y�__���b�2	��5��M�4vC�֒m�<��^�C܉ߧ�Q�8?~K��3�w��F�u��5�qL�~>N�:)��=�4�f�I7;@X�]¸��|�*<�� ݹ�ld�Bz�}S��MH���L����R0y��H����)E��H������{,k�n=>�U/1���	Y��ۂ�_D/���>����'ۘ��y.�is-r/a\l��ۛ˜�Y� �*s��U�Cu��4l���Q�����q���A�6}�+�	{�|`/��">&� ��MFۖ�@걝g[Ռ�\(u���{a���_}C����&�1�w��QIm{D���H��3+W)�F;��Rz�U@m0�41��>�2�ޑ��3����x{ЫS8[�Yfr`Cʸ���ۨ������v��u���Re���ڙ�σ�����{%n�W�8���-k��{�txf��%L�n�6_kLRXE�r�`���v��u��X�1��v����s�]._PB�o��� �@> 	�H��� �
�{x��N�4ky���6 f���&D���#�Ĩ tƶ�H�P����1��٘�-$z�DW(C�P^��z@G27�᧞ӈj�^��2j���'�ౢ[$.�Vrbm�|&����9
��͎X �0���� ^��ܤ��}b��͟_�=�T�tC�GU��~gੳ5|��q�~:x���M4hڶЄ6���{@�9Y���)k��3�������*����iX��y	e��\~�),wJ�k�� �0�M��T`�eo�.<�{�ZZۢ�"���j'1��ra]��
}K��� �O&	K���,���.������n�@�K������"Ȁ@1�=�$�{BA���^~/x�!�H*K��t��.��=��/r>H����4��Y�IxUp=�]Y����(��B-�	�Ț�qvL�u`3��v�+!�w �'U������8&>��WB���Ͻ���d9��9gh��"@s�D��e�l4���M��43C��rc¡�@��y�8���S/��Q���(���Ǹ��7�
T)��ۏe\^�����Gl���	Q��=#xܫ�9.�L�ݞ�P��iu��#b�� ��@BC{��r� t��ۧ-�H�S8�qeZ�5V+r��Tc̝�n�Q�/e㺄�f�sT�;Qh���Hse�{���i������K���Ѷ�:�o��[(R�ߤۃ/�ik>�ڙMr��+7���~���~E=�뚴ʢL��݂�:�mg/���r(���CJ���ض�����u�����TO�3�{�e���1�ķjt�8ͯ�L�:F;�{�98� ���j�B7�c-�d@���K��l"n��l��׀�>�M�p44WP�B������|LS.~*=���a� ����-zz-�6�L���6cx��.��%��~u�'-�d�}�0�p0[{����)����i��R\��e�)�텚�31��1�H��1O]Ŷk��Qz���\{�F��vW�2�vb-e����س����H6w�Z���}�}�����@���o�i��o��
�I�{Zź���I���`�,'؅N�"y����%��~U��Y����=9�1n�+�Ҕ:���1��>�� �v�xf�29���b]�i�?�h~2��A�?n�}�|%{;��ğl'�ڠ:G
��и�0$|�G�pЮ��"{���n��tFC�s�ip����]��.?����L�ڒ\ǚ���2�j�:ͦ��
Dk��b�#�P���: )<��	p��nk�W�N�B�UJ�F�ieY/S�A��O�{����),�&o
�U�� �иT�=�]gS����֋j�R�/����\�W�a&��_����z�|���� 3fzE !�0>͊�#~��W~���M���]��g�A�;?= e�>�3�&�z����8=��c ���`�|i���ZWK�̵��.�5��C��и�0�H�6ΨGmDD�:�x�Dz���˸?7Bq��A�et)#ge�6�/�p�ԻcG>��>�v��?+Ô��@ĉ��D�1����5��
�uЁ� \���u�-g��0g��]J�fp̜�����rt�z_-w���.�𢒁fm��{;�Ut7<���B�oiX����)����ٌʷ�I(k�r�*ﮡ�i���h��鎸~�����1�[�cz�[�����m���X�k���vGf���;�����»�n�P�}��#�����H��=�����A���Hɉ:�n1۫#���7fn;u`p�sb�g�N"��w�B<A�.���K��+vC�JW>�t��Q(���"2�X�����z��9��V��\1�Bg���'�/�&~ݲ����7�\"n�C(eT��X^S���//�@W涢����Tv-����SL@�Yi��)�G;2��lb��:0��]��ôZ됷�/d8�M�eӪ�=��'�;BA�M��ӷR��s���_a��Y)v!��w��zq|D,D,P˷���� l@>j�?3)�i&�J�#�@`��kx�t��Η�1�U���sߓ�sI~wo�
�:��ϧg�p�|ګ��>~Mz��L����v9��EG����J`BƙA�n�:i9Cv�SO1�'�|<'f�Ez8�QG	��U�T��|nWf��j�xH�g�H�#�Mk�'^���N�0t&���!����N.9�d�%�V1f-y�^g=��=�v�ae�:�,�� ��:�ޙfM\�ٙ�@m��8�/���!F��|e9xH@�
�lY`b���;�=��Kǉ�ĩ�ɡլ��^�)�9����1���&N�#�s�D>���	����kJp��jo\��b�n@��X�8�	�B�T_*�I,�*�3'��˯�}ٿ��uB6��-=q�d�;D��o&�k���0�=M>&�C�uӗ��ͦ^�O�l4b��X�U��ر~g�ob�����j �oL&�O���fu���N������0�x�NL����LΞh5�\����;�'���?A��U�3j�g�����YG���sG�w]Q������v�:~��h�η��ܺuFT}a�Y�1
:)����U$�9��I[(m�4*L:~U��P���N��K��0!��(0G�C��D�]U�U���>��SáMC�v�n^�[V��8>�:��;JI�㽮Ȭer�2mM�ep����� F���ei%�r+�3���9�wC5��P0;���PEdXm�k�Ǩ������:�zs�ZE�,��%�^�B�R��ϻ&
w1��$O���E���CD&���gg�R���ks�NuM�W�V�#=+^҄���B��V0�F����{g�@ő9ޯ�A6��ޥS=����̟w�3flkk��1I�n�T=�*�������y`s�K�T�_w�Ok��|�L 'ѪjX��ޡJ��[.�T���1����ww����?,��X�<v6FW��P�޹��:�t��Tx��n֞�D�	KW��ӏ�\dS��ƃ�i�ߞ%`�@F����ϒ�'�O�zh]���atۓ�1�y���jjn�'s;�֡O5�j_�'g�2N�Y��/�D=���*����ҭ��}F;����Tk�K�[I��>U�wJ<W�2"	�x�b_��[���8�&�&wp����<%�ENG�(fΑ�OW����^�h���"O�A����M&U��=v�E�{��?��S�z�\�N�g�������9vj^�>2����v�f��W���0t@ @��l�8�0�+*�7m���;3���-�˼S�t�/pb;��	��J��D��!nJ��r�_p�!~�@��ϏE���b��ŏ��ـ;Y�g=5��O^����M��6�\��8����Dpb��B �N��o��V��2`�x{k�C��`T3Q����Y�Ih�i:r�(��~���2��PH��S��l�_��ԩ�=��Gz*��`~	� Y�lb����CUx����s_i�C���=9��C���N��T����,GT#D_�?g)B������;�
��y�2/p��&%T���aMX�a����U���ɶ�c�aR�ߒs>�.ܜ{��[}��!�x�SN?6c�Ȣ����+U��a���K7�� �\Y*�j�
L�����w�e��m@��� ���e���f�l�v����;AdR��(��j��(���#h���.I�լb�=q��9m��CW8fI�>C�~Ίe��/G�Һ�Xː�h�7��߯wut�߯#�>C)@�VP�}u�&�d�����
����)>k�Ώl���d�*kD�{T��V*Hs����@�3������t����{LO�#��+��ɇbN�+�m�J�^���ճ��i��.��{f��p������Y�]{ؘt C���������D!�r�]�պİ�\��[nԣ���u���ֽ���C��Y���}uҞ��}�d����� v��� �Hi�X�q�|5)�K��Ŷ�q:}1��TF�(	�E͊�q���Vv��ꋒ=�W7�rqc6z���X*I��T�^�O1�heqc�	�����܅Y��ya�9�����@_�b���ӊ@�c3��c-ǚo�5�0���tsk��.&g��{��jUyoD������^'H��ٯ��}!Xф7{ӝ�+�� S�*�6��}�f��A9�{�G��.��a¡k���N�!g �|����c4�8�S�[�k����3�f1�@.�&�5ӿ�i��S��3NAO@c�8�]÷�[�|e�w�WR�9�մB�^C ��: ߻���P�֨L�6���J� 8\{-��k�;D^���� 3ڵ<�QnS�cçbb���7β�/��#���~�~,RN�~[�e�CY�9�J��o! '�:1�Gt�3�v:;g8�'��/��uSa�G�%�H���,9�6���[Z-_#CM�̥>,�<�2i�1���6.�V߄ï{߯`���|[��t�Wt�P�j�3�S�MQj�)����U�S��D-7Ŝ3��\��ݳ+s�]ne�Uq@r�Ⱥ�j�i`J�����Ϸ�k�Yd�pܴ�HVe�4��5�"R������U�3��$�+.>Y����p|t^�ZtK^�W"�i��o>W�OU*�7gq�9���g�q���ñbj���K�sy2e�0F�ժ�V��g�q��9/���c��c%avU.�͑��ΫK����L�oN������a�+���<'�y�U�|�zs��uX�D�$Ow<�I\]M��AC��f��Z[yg���n�^��Jm�o`���Ď��
�5Uu/3u֚�Ҷ������j���5%��9�U�ڸu��<�s�q=�R4:^j��.��#����+��4�'�;��}��ڵ3's{���i;�%m-Sy�J��܇��ath.���Go���}����d��R�9ر��n��{�e�u���;�B`S�v�>��R��:wr��ܪڹ��S��f��hϦC���H��P��w��:6�f�S&+���x^�hVLQ�Q�1�f�7�����i���UM>t˾]���OUU���E@�)G�H����f��w{�/�VP=ض��nB�774�*�J�UX�b�cZ�Ǡ�B`!u{�K��-�A�X0��_��Y--|�hX�+=���0�)��0����7�6�bW�����Æ< X!��~ ���XgM�;#�c�f�wp�_q �����LB��"Ċ�p �u�x����2�v��g6�ڢ�ud�w��gX�&�A��J�lА�!���*�u���V,f��u�yU�b"�]4�����iq���8�e��΃h��o�_j����t���.n�KyU�{��^N�C����҅yƻ9ԛ�]��v�^�Drh4fT*F��G�����˕Uŷ�[�jU�kj)��]��g-�s^*��KV��N;����N�Nم*wkJqlIj�c+ZS1��6ؘc�
�6���i�cu�^ʧ5�w/W]L��L�9no�����+!_�R����I>���"���ªJ[4��MeT[�-8���1J�r�q��6l R�m��UliE'�cgY�!6gt�:�j�J�Y/�2�t����ʊ�yu@ON��q�I:�v�V.�wm������{o�Ԓ+>�U:�������i�y�5�4�n�\�!�Ig)���FqIAE������l���/eF�M�<M1y�g��
X��p1�F�̹���.�,Z�-@�6N+F]�u�nfŌxT�tl�W��/M��֢�U.�m�/���ګ���.�-�y�j�L��9�Y���U� �I�Q��ҋ�oT���i��H��1�:z�Ӣ�UmX��׮���v�ӎ�V8���ҼzWj��O��m�Z:V��L�W.�0�c!َ�+�L\��º��f	����Լ����C��^�������U;��'
tv~�{:�=�����xvh���Ӈ"O.��hZ�R,T�4h���0�l��:��u\��-�����8aÇ��uSt=�jC;0��<�9d������S���GƏ���>><�l�a������Z�N���=:4xtzp���˺���Qd�u�6a�a�����[�Z�&��N�Fo��]�B"��#�}��d{��'>�F\2"��IB!0"�ݪ�e�s�u�^U�P�P�je:v��M�f�
�L���tM��
������5j.D�(��{�_j� � !:*�ۤӦ�+f�4ӧ�@CQ1�2�!8ۉI&Oa-��@�@^ " 2 L��e�0I���L"0`A�,0�B0��r����_ԫTJ���r������Ԁu�&�\{h���{b�����Ȫ�d*U�ڊ�G��n�Bw1�T@�5"� &Ɛ/��+
o3a����^�M�uɌ��5 W��o8��>�u}�VH��;90��sE���}Bp��PV�95���;o����Nj�p��ys��(��JV?5��1������Tp���蠻8�h��	 �i%�\�̴{����lB}.��.y���gNt���BXՄu��bz7"A�%����X�DF���c�dKM-�k`���Q��c�X�/�"�6�d��p���u�\���w~�}
=z^T?�
����*�9���e�=�_/��ެ)-�}�l�����4��rC2��֛�)=56�zO>�1�>G'�����mi�-���t�p2^���r��n6O�X2NB"���j0.EF���db����Σ��d��ս��.ؘ-���s�=�3�Z�t�0E���|"I���=r� �{�{ὡ�H�awN�{x��iS�9�o��&�[�ވ��ʐE蘥��W�T�W�ޗ�<�xx`�E��F$V����˞k~����Y�[:d�4������
�eG���8�^wC����	]7+oc�@��� �'� ���䨬�՞��L׿��kd`a��{K��H�}/�)uE��%�$�B��x�ͧ��(�Վwz�Kx!	�X��Ÿ���1�k�Ca���,J��t�{��'�R��^�^G����L��
��K�F�O�/d��cٯ�a·�}Q�;�T5��^*�Wޤ��1�������1-�Q��ߠ�׃�(�H^E��Z��ni�b�N�b��#����I��-i-�U�3���@p�с��E��<�D(�C���cP�>��Tz���+�!�Tui<̋g:���-{ޫ�g�z��0}����� ��PgÃ^r����v��E����T�dŗOJ׿	��T/VM��ғ�u�m.���p.ޗ\H���fh\J~����S���I����d �o�w�9��)>�{� ` ;�ɤ�M�c��#~�m�o�7�Z����ݵ�u<���`^EwO���0���ty��I�SJ5aں��m�*$������1da��~���V�w��b����Z}]�r�i=>�m��63�zd��pL�	�!�v�	�4�����n���*8ag�h���HHb��v�}�|)`��!ꪋ�I")iu��������1=x�}Nc7¥T��=2c:����ۣ<����T��j�m�`�	+��p0�F�7�Kĳ� ��L����H|���Ѽ�/%�/t��{�dUS�0��v-�5��<�ˎ�-T�a���S�"�5� B N��?�d�z<P��6k�Dbn���-��E�#��T�V��k��A�ה'��tQ���8I&��v��!�<�:Ȫ�3ɨ(磱�g��9 F)��#����=b��B~o��N^�mA������n-�kf�#�'� �$p�˵��@��:�,�?@��Z��q���GJ1���iGjuO��Z��}�������;=���B�T���ˠH��^�\���9y+����k�x?^̖���[zׄ� W����3-X6P�pm�����S9;��,���_���Z�W>ާ0�(=u~�ޠ��`=�p�n.P�N���p<�w�_�z��X	V3]�S������E��3ߑ������I��3���?�vVd�=��Ǯ�H��2�����$f�7�/!eK݌e5���W�^m�L��|�1��
�K`�EdR�rz؉�B�e��$�)�:g+5��l\@��Z�n>3ƴْ���D"A�M�Q�
0;�bryIפx�՘�fb�n��,84�qumDN���\�'v�֩x�^�u�<�y�/~I�~O��KKKMh�m �kY��?�o�4�C�k�!�Ik�B.l���N�����X���	�0<�s�6�\X`+���V4�j�J=�5埻&�p=��ʳ�/�#A��A2
���Cf:��1l��SLj���L��t�u�Z�}�`��l �ýSx�|�5�Ĝ8�~���5�0�����9/ٵ] ��Cm7��pP����c�S��oP�Nk�C�Q6�~��hP������f+V����\�,=<�g��0�����;W���!%��P(�/��:����s;i�U��N�y8�r�G	M�X�G��U���vvF	��'H$�{��kާ����z;���Yxhcq�[ӈ�-����S�N�{b����Hϻ������&t�!��{� �G0�Z���zr��	4�!)����zo���6�O�6�9��������y�C�6�:2#����������aY�z�a�!F��p'�Z�k<�<��p�1Tc%�����/�bY���\22"D��aq�>�G`h��z�ғ�}TB�O'��W̥!����$$���==�c�cF�)��l���MS�����Cn��֬�^�=�_YR�+5.�q�,͒��;��W)�e��\na�. 2�S;��{1Y��;LH >�v����Z���?4�Xo�o�S��Q�Y����Xa��)��q3l����	��4"
�`�#��Vg�f!F��7�ܲ(LwzB������k�t�m��<��>�4'aE���\^���0"�sPEeL�VMƛ�תܶ����Ouzyu.5��[�����
��?7�F�-{n�\\�1=�YF��ken���Q܄xL
*�#�N��tצQ�~�;�4{�r��"�,Y���x��·��{�)�TC�k�iiU(hx3�}���A��dE�g���,�Bf�Fꑦ��C.kK�Y�8r-��)�3�B���6t��	9�[S���ug��fQ}a�1�~���3�z�� ���Y�E������"0@�G�Iy�3�wzW�r��ik h~��!�~.�u��eG7
ߛ�[�Ph�j�P0�@��wlhz��4\���8x[:ms��U�7��I��K��*�K ۯ@���-��=T}3|��S�7�
Y�Ϭ�2�>�j5�7��4��J4���fycL�Fr��*T�n^���鹌�E���&��]a�pB{G[ImE=;i����sG5���=׷�]b�2/c� �K�ҏ5�j�>�[�{�e�"�UN٧���]c's^�n2�⨈b�h��1�f�ٙ��*d��?�c�X;%�w��3?�(6���c�>�P�r�k�C�<��Z���b��G�@w����G|��&���kvb�6˸\�`�Ɂ��`=y�rxnl2�����t&4����p����ߝG���^vR�Dl���e�����r��<@�7������nȰ�ӌ�*��n�������L7���T����U�������'���,?��c�3��j��dڌ���"�-�������p,p	����/��Qз%LI��=�"�[Nd�dU]ό���Dşm��~��{�=����#��!5Tt+̷W�̑rT�BDUի�p1�(V�?�S�&'#�i��ʄ��釶G��H�gKP��8��9I�v��ۂA��ndZ!CT\����x竂w�NB.�FtS�=�F�h:\����N��z|�K`/�������:3�����o�6>�1'�W�?�@덪�e4�Y��wP�]Γ��z�Iփ�>�1�I>����3	�
��/�cM|;�.3~����%�d\�e���:�K5�a��vk��N�!W�r�.���ƮY=�Y7LE>�0�d} �V�Jz�Z��,L�+Fi��,�m����};Gc9o��c����+���_�@Y�y�k�CB�L�>`;���7�V%W͋���o���GQ�װTx&&�н��l5��{s��L#),>�Smu���/5Pͨ\k4WHf��w {��<(`"���T=̅��H�9"ں)�։���J	���9Fu
!邞��e�Wt !�gT��Z���0EB3�c\�����(�l�w1��� C�`�A��sϢ]42D�ȵZ��}��w
æA�֣+h�M�q�ǽ~`����k?��G��^��X	Y~[ɗ����Ը��2+�t<�P�P;�o<����5�*f�_�y���3k�B'_�O�$j��1���.5�c�����k�-6R�)@x_�n�H;�V2-��]jՑ�8`L0�M#���a
�gw�>.�ɷ����n�hͼ*����j���z�Y��g�:���"y �	�
%v�g������e⠾��=& �OP�СkА錋�k.k�q�)�7�w@!�bK,�lщ�@�s�~_��ZZ_o�� @ӀSߨ9?N"y� ���z��P��-�	�>$���i���vN���h^����uRB�rA�`�7F+t$��D&c^i��Ncn!Ҽƻ-1����sS-�vR����uW/3+"�:*>�9a���\���:��
�}��s1n��L#~�7��m�$D��K�,�kz�1���}kX�B:��W����gp`0���S=�Sc,fΩ��ͻ���j�\���|��dWӓ~�4@d"�nFP}P|&�)��-sQ�;.�m���%��NC�S�L\r���A��o��*1G�֯�Ւ7�p��Ͱf��)A��%�"DG[�D�Q|��ܶ����Sl%�bɈ�����,�}U����Tq\����#�ȷ^��t�C"�c������zdi�� (��2��P��.x~V�7�5�ҝ��Ų�x	����ދmj����|��(ߖؽz�(/���,��
�M|9|�����s��h�E�C��5s�b���َOD�2��ɥ��Iq��=���ά��`��&�2lG��. �UG���xhe�e�G�c�Z��0�^Ð�/�u�s��\َ��7a�m*�0��۵1X�Ϙ�P���5W�p�Z�~0�}��s�s]��\%Fq�x�O1X5��`Z"�`��V�o�$�hY,g�Q6Ag�l`��q��ϩ����G�ު�qM���댱�K	�*u�$	�� �>7>U��K�cwJs&��ي��O�Z���1_Պ�eb����F1�_`�����$����K]ho\�dj�Z�v��ab@��t�:��{쨾�8������s��ȸ�:���PÓz4L���C�o7����:UNd`�!��,�]�a 1�0 0��}��aJ75���Ђp# ����z�>0�A?��� E
����/-�<ޟ%P��ӑB̰a���<h?.��}�D������r����d`8NXd�𾫚d��N8Z�^������tK�I��c��]��!�BB9���"�䊁��y���2)�g_���\�	�����}緓���.P4�M�M!�K;�ǆ{sB#��H�Q��NAOX�Mp�:�@�T��n�֨4���̹��ٛZ�g)���^za���,?0�%@�I]sO)���@Ǆ)��1���4h��Aup������"{��
�`�T�v�?	��Z��M���!�_�Yt}���� �M����gW&�>�3��V��Uu+*��?]���q�����]	�@��0)!#+űDKH�@��,��-������]/�lN���-�{��¦��?}�jf(8&��|B,��z�p5�Ӏfz;R�6`�g��^�mv
�#a%�/-�8�@5�Q�2dF1)?Bw�ؐØ�c�nc?w���OuM�w7~$F,2V��{��S@��β8Y��t,�R�}Z]�I�ݘ;��k��C�{��ڢ�CA2Q�  AtX�J�r�s&+�A�]�/i��E�AH��X�l(s�tvp7δ�鉫�J�ʗ�ss����RK w����w� � fԭ$Mj���O%�� O]&'T�t��hCMc\9aM$���i�S�H|p�16���f����E2)H}�oI�9E��1I���EJ��P�8��4x���GǦ��B�.���\>
�m1u/�Ʒ�YF�r�$1�Qx��E�5x�;��m>�N�󨖭�زtp�4�+f|�b"�#z��ުk�a�-K��ێ*(��尡�D�12;4=�M)��\�E����쐂X�@' ��_F
����x��,^ώ8Þ�nO���+z�sWG�����it����T��;����YBOR��^��<��#��fs�B�Q����c[��U7���`�W"nw@_!���:	���!�#�}F��fԞ.��Ϡf_h�ٳ���Q��ͱlzw)�d0[Ćv���ɨ�B=BX������kk�.�״�d%ǯ~��;`�s+�`�8�24W���B5Tt$6Q;���d����.�ϖ��+7��z��O��۳=�!s�ǝ�Kq6�>�P|>�)=G���0�$��E��/���Ri&���f`��+-�nZgT���K*j�ȳ4WX�*���U�nvm+���F��+#X��{v��=��1h�]8��(j�n��*`�l�N�,��%�V��x鑢[��%(����Z�ewU��oT�v��c+b�W�S%-R�eFf�0�P��u}8� �z,8u�8�o:�Y�Cz�d%��S/�������[��Ll^*v��#,1�v��V����íh�=���-U�.�%�+�V^I�ɪ�U5���	%o�gz^S�q����3���a�$�v���%�*I��ef�o�;&r����V��p��՝�R��!]<4��ϒ,.+��7mM讄Y��v]K��3��n���S���U�yhJ��:\y5�̷��ڛ�[�CtP�/(���&�hh�t�3F(�HݜN�j��S����ȏi��\Al�0f�S�.�� �p�]�:a	o���Z�ؽ�%ʍR�R˙�"������)�}�����ǖ��:��hl������M%T����/5�t�����Pꝛ��&�1ݬf;���!E!VFp�ɚ�ZwU����ד�����v�;��U�~���"���h>��^
N'Dc��Ն���%Nñ�-���ځ�B�D!��`�C"�PY��cM8Q���AoA�'�9�&*m�h����BD@�(p�+D<bcl�U��P�-�#DCB�+�Ƅ��Z��������'ӫ��W��n��L{�+�K���'k�u�e�N�q 櫽/Bju�z�^WY�J��Or��e�r�+tj6�w�q�)�����Skj��T���X�6x^�K}�1v��g�S�{��)*؍���6"݋�u�My������İۏ�8�����K�@����[@���-�tʻ�mj����᳛�r�J�â*���%iɘ�i��YkB&��_'� �2�^V��m����V�`E�LӲfkS���56ʃ���Zz��!9#��m��_��D���w�JӤY��VSԺ�����0��mE6r�	��E��!Mڠj�\F5��d��m)Q:8�L8���M�79i��I�SZ=0�`�O�wT����2�Lq���'�A�<�F����^��PZJy�9�(�u�bN\ͺqh�3zwiٕ�q�i�*�Uc�uՕ�Wsor�Z��$��;�yG��+_m)�"䡋���w_6^�:�����J�$�^�۷B���fvkD�Ir�b��ì��י��`�;����o�����<Nܰ��'H��(���+T��WTp��jޤ�o!��F=q�߫{���/��(��9]X-�f�\�O���Æ���>0�5S����T�Ku�S��[m��WV=ޣ�F��0�^������^Z�/C��:�]�wr��Շ�F�>0�����m�;�m2wj������׿s_����Zܰ٣Fzp��֫%���ݱQAi-����>>>>=><_m�ʱ˫F6�-^WJߕ���'0�ڵ+�jݞ�7�����l���M4|x|||a�^�@��-\1}�c���8p��Lޓ|�ke�;��n���_���4������ǂ��xt�C24hK���/ί?|<t�)��I]��W4�R�S,��^�-7�b�����M�d�V�QuP������6�������3�д��hD@h~�߾�iKϛ_���D���M1q�z�z�oM��	O�;��2�68ͳ$�H�����;�7KMz�KJ=�rB��f�C�/���
 �:�L�/��]R{bf�nx^�b# Dpve��L���-��P��G��嵅��w��n(�~��&��ѥ�T$ �2�3	Hjg�y�˞�G�P >�����JX	z�LP�SdW���62�]{wu��w-pW}�\��dt*�W=��
z*r�-�z�i���9[~��y�i��`�ݴ�f�l9>��3�������QU�a�#�>"�kf�j�p�!�%H�"���y!�d��N:�`Tx��~�Pi;T+����
n�$c.�`�T�I���h����b)?Z�g��*�r�~=��o��_�!�����h�2�ۖ]��y[�X��Q��CR���s>V�-��5�������y\�3���K�mgnP�̆M���w�1y�Mm�1�;��+>;�|���6~b">S��:f�6��5���͙�Ǘz,�C�9E�e��i�F��ͦ2I�;��UϨUf���Z���vqY������`�Z�E��1\T�a�W�k��5��S���Z&u���u��s.R��Wٔr"WJ"�(�{A"ݛ�O��p�f 3��=Q��9��`��/E�����e�ȶ����&��wJ<WA�i�W~1s[x�s�'�Q�Ch)�! x���Ns��e�Ѭx̖З��k�<!��Co]�bG�y���;> ��3s�|�^��YHC%��\��쮑����@!�ʴ۹ٔ�_V9%��N����]��&7Ņ�@��0�?C�|>��//U4eFl��v���u��I�˖M{��� 4PFp��<�#�[�\�
���&�2�nF�"��%�>�!#
Lvdo��O��0d/up:�Ȓ�{i�<��|sQ�b�S����gV�0c�
{r���-�[�E���-�e�{yЧ�<��U��f(V�&˞7e�A`�X�q��ݾż�A�KUt"�X� k����~ה�fH�
� ���ڋ򩓭lǽ�J��I������e�����)Y�c�1�/�����FWP�v��B�Z�+7[�����6jpl���F�vbh	�"&�v��(:�6c��zư-i�pA�p%Z��'��ʜaK2�.1�������G�o#F�i�ˇ#���i~|.��WZLS��a���m^�.��%q�qR��Xɓ���A5If�i�xo�7�V���i؝�x���ò����L�9H�&�;�zS��CA#H1H@�����"�T�5K�y�R���7���{��;��o����41=Q�5�� [�~IW��خ�C�ot΂�y��li���\�lL�Y)���L��~��%0X���?� ��)-��[�S����1��d=��Qp�
�Ie��;�ǐ�r�D��.+�N��zds��ψ����^�u4���a4w&�ܚ���34b�)ev�����_�DȜQ���AN���,�����{3�K�՚!Vdz��)�V�&��_g�&EL�̱���^Y`��oX�o&T3�coE댍�C����+�m�1a�52N���(i�^�r|D���5>�+Z���V��j���3n����yt��u"Ƽ��$��]ٵ�:Z(*����A�Y��;賾��a��{3���~*C g9?H�:� T]��|sB#�@����� �k���l�1?����o���G�b|�5·ƍ|O�HBSxP� !+&��S�e~UѭQ&pZ�����k��uw��5B�p����U��`=6A�kxH���C��t�/f<���!1B4�}N$#e�e��3vŋ^{�Y&��v�g	Z�1�(=�$Dnڲ��g�%�!�=O)A��jP&n�Cz���n�0��n+"�مe���%^��P����l����n��w?.}�-�Ҩ�ѥ-,k�z��s��+�,k�}k��[6��4]E14���.�h&T{(V?$��Cz�L�=�\����~�a��&���ϝ�4�겦����3^�G�ؿ�8���7��۴4���s���[z�F������{<�HCF�[���?d�Mzs�C�j��C��K���D�2N��6��(%Q��Thw4ԋ�D����ή�c+�����]0��SwbUm�5mkqyj��0 k�D[@I��i��[�X��W9d>c<�r
h�b������]��}m
�n�T�r��P(y=sQ�
��b�ej����7!��-��J!��:<��xtҞo_. О*y=:�9ܗ���T[H�tV�O~���1����|���l���"��ށS-�jG��lsSTP��Qkm�w'��Ut�o�@;�L�0r��l?Ͼ_��|��ȡ�t�X�6:gʘ���u7/k�:4�ʠ��5B[|�8qh������Z�� �G��P�,�E�{0!de}q��?*���͌���32ӼX��<4��W]y��"!9���uƺ�cC��60u;㶹"�0�+���w��,_����iP�:OC��%q<J��劝�oU+%<��/��!��U�]��3K����s8P����W���'�ꌥ��h�������ָq���'�r�F�ի��Q4tو��]�O�g��!�<���0���6`d ���������� נ�o��
h3�(���hT��DB�7Ni�5+�K&�K���E��C�o�ٳҮ|m�b��b?oL{��#UGG"5���(��T��c ���b��7B��^Z�Ș��y>�w�dȟ.��f���_/q�v�x{/ຠO��H:+i����e�K��/p%�ߓ��z�n<3]Qu>W2ӝ�L0.x�[+�~�qg�����쌈;�m�ʒ��5e�l7��c�K�L盨H��bpH���J#�xsP׆,I���	m
���?��%f����tB��>Z?�O7b�2�r1��U��:厽,�
�.�b�[m�S�v3�w/"�>�i��O�R[;����og;�){a�u��S��9"���л@�%�{l����e��pY4�)��q<�)�PͲB �_@f��F��`���Ҩs7�8,�㟯�=��/�o�n�q���;U��)ĥ7���{HҪ]��n���bu
ѝeS���!yK�K����<لZ�j�' q��w�V�K)+�ܣ[;IXjt��^K��Π��8V�g:�g���`���"j/�4j
����P��� �!����C���5���(4aT$��7����L&y�i��w[�y�zk!0�y���������e<.t*<w�Э�~�H�#\�G�yS�ĵl0���ug���5�V��b�}<���� �kĂ8	7@ }���UK��۴��0u]d�Y\�-G OdkChЗ�C�����!��.L��LC�@`	�vH��3ʶvV��M���̑ϫ�o�N��S� P:Ճ�خ�x�D���c���������o-�x���C=K�K��"��P���3���#�O\�f�Ϻ�����C>daS�(�E�噼;��c��CDd_=	r�ݚۦ��K�d�~.�7��ZyF-��V���'�шXi/zDE3��vEC���	L�)�tE�8���~C�RE�uy�Xa+x�P\{�2�&��#��0	ܽE/���w���[��P�M~L�qL�Ո����;O��A���c�9}��fk��LiA�KhKꉯ�
���I�3]ґ��pXGC���j!�����mM#V�w�,TA�!9á!��AkG5����۷�H���t�)�q�"��"Y�$5yC��&Bڎ�����)����P��qS�;	�H�z�ԩ9QH�{nt�F+8u���S&>�}�D�,P����� $�!��.�`���+^��!�C@���UQ��vCۆh��Δ|<C��AYB�T�	m:��S/G@��wu՝���"�ӣ;�)��:��"��}�k��@U�c��P��N���<i�z�g�U��J��������A˳,�@�q�+�x��*p髝�W3�|�r�x���ꥵ.ȹh�D2nR��C޺���k��tY�aS;NF��;$�\�Y�1�m���{��u�)�~§�H�3q9��xw�����6�:���RU�����@�#n1�Ɏm��HI�{J�caB��1 rf�;�A!��1��U��7qEIX����d���m��^E�H��\t��ƏW1L��c�cs�H���0����/�⎫��-iDk���No����B�^��qq�״��w8 ��T�4sn]�
�c�\�y;D��2g���]zf4���E2}�o[�y%c3��1a�.m��}e��T\�֎�2�2�L�Ƣ�y1��_�)���^���J?
8k��Jp��[�A{�i��)|v��桁�TB�Uf�ZzvHg��v��4Iʫv|��������$#��A����.���+�J�c\����J~����-i5`���[��u/��Ƀ��;��pS1{�p#*�]�3��:Q����8��wt 	�/CxKh��9̸&D�����ö�:R'Ѵ\๏I��6=�u4z㎑v7ޅ��.d�-�P7�%@,�(����2�<�jC���g�ZL�.�F��[Ʈ�n�w�~"ƨ�� �-,���p�O�-���<[��5�,��ʄw޲�4'ʓ�J�zm�KC���ų�H>c�G��`�L��2�zz�c��}�g"��"tt��G0b���d4��v6l���c��ծ�IS5&h+Ő=�P耻z�og�R�X�l���G�"]]�b�?7<9�,�NlE���H��:���	�z���8�u[oq<պ�4H��j�nNI5j��{@k���5!�e�q�\��b�>Z���|Z� ������)+u�p1w���5p��|���[L��(�����������wB�sJGX��l�X�wQO�o�Qfd��Ԟ[�7Cm\;5�6c�$�S�x�Ru����q�����L�HW|\vM�O!��IF�2rŷi-��w.���"��CZU��.id� ��ACm3�ɤ�Q��oڋ�]j�ݖ��w���D�|��:ֺ���+���Ӯ��E��T�^�m9�<�%���Ʉ1��ȼr�>n� ��7
����L+�=�j�v�+��A� 5�M����&6�E7&���<��ˆ�����tS󩚼�^�Q��}����o&.����_���a8m�S�3T�+4�?l��U��;��� ����� {÷�\*䔡}+ы{��� U����������PM�#P���[�#���9�S�� -P^�2�-dμ��{�L���n��v$=���E���YQ{���0����U��$�F̀k3���~W��b���#*���Z�Nj7�_b��
�	�.�^v���4������?d�M#vt�>�ي�9��&�FvN� ����R'���Ko�.6�5�����b3�d���v�q� hj/�P�E?�OS��rkCeu[�>J2�SR�b����3�W�5�̫sě �z!`.ۉ��'B�o)^�Ŵx�McY�c�B�P�"���A�Ҵ��;W�H�F���1��d(�-Qff�'sJf^#��툞l���v֫�gx��|s�~u*� ��-�S�)HW�Ry�	��T祝XƤ��|�I�:^"�7�Y6Ap�X�w	us����.�8�5�B5���*��LV��&�̌�?�#̒;��hMM�n� �l��3*��Dd��x��[A�NsKZ �<�$�C`U»Cr[�x�+vM�H|Un�h��9K�9��W�z�=w^S^u:�U��k�������F�[D>]�r�\�Өܘև�r�װ�d8�2=��t��L<6",v��-�Z�(T� ��ߔ,j���~����9+������g=?	�tt���v^84�X�Kpw:� ��OȈ�<�'�ɾ�t� ��^�y�^�̞�ు�S����\���Ó@�A.�N�u���t��u�`T�{M���i=����=���\c#Nz�3Z4UN:��.�ҵnn�^�˥`�K�3z�1iclB:��Wp��|ss��+�j�z5���,;{@�͜qκ�еm�)Ƨg#i���s/U�$�U�yw9|x
$;/�n�o.�-Y�7�T�:"\�P�ϵP']��c[�)�ٰ^���$f�"U�XR��T��C'
���K�.��m��bSuU!c�z"�fŅq�R���RM{u%ݑ���yI���v�g�b�H\<Z��h�Y�n�֦Sc��\2�`�z��[2BH=�n{qY�K���iŲ��T����Jŕ��QJMH����0p��;�r�,�ނTNJ��nn���_i�!���Op�QPكv_e�����B�۲�p�;�Cڑm��Q,O�xk������c�/;#��wX��otN9�WRS�vYې��	7��N��ZN덠��:/]b�i�&Y�;O"���m�mTW�w$GJB�ͪ��/��O2��c�!:F�c�2QsF�0i�tm_-�+hS�{P�ZVg��G9/R=�{�*�s8Mon+�3��yw*�˕ۃ`���ۨU�U�2�8*�������w�.�K�P��[]����g�&L�z��5H��*��c�֌��r�Ӣ���(�R� T��A����[5����p��{*��3�;Ef ���2�h�j���e��Ű�oA�X�|����<|���y�wX�X&�k�b�U�N��J���:��84��読���>�UE�A�������m��&	pP7�kȄ�jX(��@��˴Xb��Рl(B���t����Y�����|���E�hZUD����٠�9��m�8����k죛WgļP4��J�:Ome;AGxX\4e�:�Tz�rUEĜ�����^��U[5�.
���0� M�=��q:y]��ܫ6H�̩u�dt�*��U7Fm��FK�i�`��Y[ϔVƺV�k|�G��<:���\�}R=6�k���bZmok�t�7M㑾+J��
�zY.��n�^÷-Ӽ��Cyg#�J�,=HRf�M�Y���BùY.v�)��/)�r���iE��"M/���V���G��x�����;��*[31e���Uö�>�Z��ժB����4�z�q���W��ݦ�����Y'4���jw�G�4"N�Y�G˪�V=�Gt;]NtY��<+Y6�a���-C���K�nP���cm%�`��Ri5Tuک�c.�ٽ��@�C;V��W�C�l�1�}�Ճ�\�ޮo��%1��S��	36��j�Š{[��"T��^S����P���V���w�ܳߺ�|T�iR=r\p�3�n�dj4z�J�s��:qN��X���'�UO(�ۙ���m��@B,H(P�ԧM��1����OZv����m��N��c��8�1^���P�����F���԰�j��E�X�6��fr��"*}��k	Oqw����hn��On�ٕ�[*��ԾчG������ϫ����~���Z�Ye�~�<6h��������Y�^����&���WWL(��nIO��3�v�F���8a�Y�Uj��b�1�)��J�����Wf�ta�x{��_�v�:��`ґI��jjU�նZ���8p�ÆW�Єs_<v(}n�7��2$y\���WW��^��}�����M#��DƐ�d��x� �.��4l��0��ut�Z�oV��x��x�W��(ޗ$bYk+G��j�o
h������~��E����n���W��t�����x��H�!�]�M$_;�<I��>"����(�C��,�Ip5JdP|�k�*�=s�	Z�Vt���Z�yIYy�)��UTO���unUԱ��gs'b�sDczC{&��$@0�6�Ҵһi��V�S��6S�`��5pY.Sf7Q(���Me| � �e!�|��c�y�5K����@ɖ	��G�'��e���3������M��|�'�D@:a�S�T6[��	��bDM�83��F�ii�1�	6��hۥz���:�SX��ϝ��U��ѽ�d��j`��Čo$�:����THމ�x����ω�����>1g\�/79�'W����qgI9W�[�<j�`�]Y�[�7��7�wV��Z
���^���a��c��!R�����1[̟���;8ٸ�^l�
��1w��'���dnc�� ~�k����d�+D_�5�J�S���E��9Oi֕�3��kݫ(-N����ۊk��]}��
͉0�7�w�Y>��O�((H1����&���E#{Fn�@�q.[%��~���#���k����@GsʡoKt�C�mW��4�>��.%���^r�G���𿼺^�XəR���EP�}*�)�В�K<���Ӕ�'���ެWk���+�6W<�Ѫ�4[�A���mY5G�`�ť����(�Sb����4Iu�Λ;��ZY�b��xQ�X^�ꦨuWwd��/�+���=����;  j��U�Z��*F��L���=�[��{��#�#Ԫ����ix��8�/P {F%3��}VQ;��|��ԣe�%δ�髈�G<�*v�����CL>�u#�[�Eev�]]Adi|����תX ��S����@��%�����ؑ��k�$��[�`$a:딿�̋��P=ɵS��9���8Ja|S�N�x��oq^��"��9��n�D�G��lf�. 8"`d�]��F�T�Ev�WWyo�XBD�bh�#�xA�6Z�i��CZ��@j�����z���7�8��*�.�E�Qk��w��@\a�p("��Tf��;f��5�eS���1�d�`��2Ly��M�����m���7w�f>?�6�o��+L�:⃍��[#��V'n�7�3]M�|X~���pK烣6�z�Ӿ��K)��M�/q�0Y��}��
;헷�O��,��q��V��CBe��ˤ���:� 4A1�8i���?II��MP�O2������C��U:��;��W|s�Ps!�\.���]z{g�ſ�j����WQG�O��ۖ|���{ޯ�,ư5�t�[�Ze�w�*�L��������7�xH����5a�\�+jZJ���K0�5�eEړ#�%ӽ�\�
0�Bs��+[�7�;�[���V����|��mk�V�^i�uƥ\�][�|��Ǝ��n����R����bm$PY�]�k��g*��'��B�#KZ�p1���=+�o�y��c���}(���	�]�}�#"����`��]ep�]��jSw&�wK��Y�ړ�u��+�V^ëh�����V����θu���/�>ZQsDۮ�E�~��q�p�w�jEB����Ԩ\��c�hn�C���˶����X��f���<46 _����ҫ�}�Y;��t��0q�2d(!��[qԛ݀*��-�Ό��L�OA���:	S$h�����C�\��fI�����.���q��1�MUf��'gbh�zpWΎ���5˱r��K�SW3���l�[H\7����VK�t=pN��]ho\M�9��2�]ɺ�IK$P�" H��� 6 � D�e��x��o3;M~@6�c <B��E���-�G� �쾑G���s��I�Md��;E1���h���e��T<_*;�������E���/m�g�nh
c O�a��V�a��y���Q�2��h�E�|!��i�:�3�+�!`��]��ސ.�R,3�X�O+i�6�z���`���WU��;㘽��E��7ˈ̩���p���d�h
��9>�iKz�8��DEp���_"�j����рu����v�����o�5d��Y�)[Pi���k{�~���n�H*�|��W�V��͌��O�&1YYMuO]�h�8�����K֮>V���O�
k�F=hq8Yc;�l����Y�R��59�;� �8�f��o�� D�b(��b��찴�~��أ.��A���G�vBF���C�O`�����]5�c�;����f�m]e�f��	�����R��>=Bv��Wwgԅ�i} ��{��YQ1)�y�2މ��s���_|I��\��v�$��;�*�m^�m�8IA=&�0,�j�Z�F弽�H��	���y����0`c���������")�ͻ�d�P��� ����D�p���c�
�R*R�N�7��d ���3�#��.떎�U칤;7��np�l���<�t�1ڕ�	��B����H7:��e�9�|��aC"��"�
M�v�cY� ���X$�T�*7Cv^�=E�r���3���l@p�
��έ׆	�����nA�%�wh�Z��Ct�24Ya�����T*���&��4�_���[ع؉(���! ���*ޫa�K��5�ǡ���|��Yt�8�غ�F�鰰��W#�n��G���6���+#�_I�j��P7��o|^��9����?���`^���՛��m���v���\T�3����fn��_/�`x�̺�:��B�g`�oP�b&3��8ܝ	�\En
8��9!�s��d�^]���'-�<�w�~�4	�8�?M���ud��F��^g��n՚�"���Tɜ:j �F���}�fQ�N����J̪#V�]�a�E\�MHhqF�ϫ�P��-S�9;X�.�g۹���*��ť���zX��G�y�c|�MN@�U��+6�5gXMbZȁ�l~w^�`��sT�3�v�<SIF_�f^��7U�_m����s�zzO흹�����rH�[���}؀�͎���tO�c�M񫐲%f��oa;����5��'�n߸��H�ї�F�ro��[@��^�E�'�O�� ��b{@�����|�C�x��tz�!-|0�އ7Q��=G��ܾ�<�Jڎ#��GN�Š�U�=Ҷ���滔e�7��o"�����V5�����Jg�|f��;��cD��Zb2�'���}�音�҅���&�-2��R"<�mya�b��D�<^4�ċ�A�R8�=��>c�D����,o,�=�0�,��Q���%�T��}�jF�Z�|d���q�Sc�6�QS�Nvյ	v^'�}��K��s�'I,wu�B�G
�.=�Je��󕿶YK�m�aSHvk���+NnS��u�բyVe����wV\i:(�̣4e#���:"^V��8枙��o3�,�@�����YH<�#C3��L������V0d%�l��	Ƣ.^觓.a74��C�sw��+Q�	 �LM�}��S|��W�_�k��_d7���d�3�+g̜;'����������	���^�Pڙ�e���Dٺ��v�.�e���*[�ͨ��.P�#>x�dG�2�#��1�'t��	�J���^��R�&A��8nk�n=S�������"'(�-��T"@eW���4�=�T>�Z}�/��܂9-��=�Ә|fk�W��.��� g^%'�ɚ�����8� ��|X�	��%^��7j�����S-~���nT3>И-GM�?tE� ����{#��4���`y@�P @ �A|���_gv*����  7F�N�Ol���� bAFV���˰
�Ҡ9�Cb��.-�#���J�n���� �h����k1/�K7�S�Z�k�M���u�x(�BGU�L�U�Ր�`W�����Ο�b�Ll
�����r��M}�,D�F��^�LGph��ͭ9���c[�mB����
�S%t��u���l��a��Ǉ��N��ӳ���2j$�̌%Fn��OQ�SnӢ
v(��a�nӈ�s���Z:���սr=��uYK��ʪu��`=��*����S�g�qT�Ja����du��NˎDjJo�ktS�"�֋�R��x���W����M��C�e�,���LG
�^k�2ޒ�Z~gB�1l��ݔ�/�@܁�o�W.�n÷�ܯ�r�p���߶���~6�m>l`-O�0���,�foa��}M.��ϧ�Uв��o���?E�uC��߫�9X,3��j�����s���a�����@FFuH
�ܔ���G���
��\��x]��X8䲨��*��x?�9��op�ɪ��۴{q�����u�;�J�����F������^��o����� �t7�D��_z̓髞uh��C�!�N��r{��,�'T���[�Ɓ�'9=VS�z���+�f���ԕ��K��ϲQ�^`>w5d�+�[޽�n�ԛ���64&�S��Bge���c"��Ʃ�pVZ:ʞ����ݗ�z�p]YS;Qs*�-؝[���B^^����-��@��8��>�b}:N;���ӯ�K��q妯o+��'0�7:�豩�~N�{uܻke�*q+�|^J�ە�nuэ!,!cC����5),ʟ� Q ��U/`�z��f(��bo�
!'J=\'�]4� ��X�oರP��;�����h�n�oT�9��Yû=������kp0��9Z,��F�y�����w,a���Ә�$gZK���p�j~��|6�q>gE���X�L�
o]��VSU���oNމH��ԍa�h�����d��0��gKosc\����7�;�!(=�n��n<��$@� X�,;-Dkhj�s��1��wH�o�xa��V^r�N3.;�Ȝ%S��̕i�E���$���I�ʺ?0�{)�����Į� ��0�e&���+Ȋ-�""���_(�5��®��db�m78æ�U:��h�������4 6��_�ה�d7H�f<�.�}�
���x�w4�'���X��bp:�m��c�	�OS��l`��MA;��L��;�&
J�Qҗg(��Ϝ��'KH٠�&�Fٸk��䙫���tܸ�Z]�~R�u�W}�Z:�H��s��P�n"�U�i��׫5��bƝS�s���r�u�[#7-���]���
q���^l=��<�����bu�H�I��1;��#�u�3��!�G����l��&\½�<d��^g�S�uMg�1g�:�x�9�Mv��4�E�S5o���������/r-S�L���`.sGD��2$�o��VA�[�����X:�3��6Y`�.�[����v3�糽�9�t0�{�t�o��7�|�������>�)�g�[����~��h�D�:��5t�Y�O�E"ܓ�l���
]Br���Vƅ�+�;����=��z	bu��!�pP���� �:�����v���;'��k��-�wQn�̰>Ue��dֺ��P���f�g%;'z��*Ż<��

y��0nh��#\��5W;͐��s|�A"сW�vV*�=�[��ҍ�QJ��mr�Y��k�>�wK�I ģge�P���[O>�h���_7٠i�q,�ܫ:zwN�8�w�y)}��Vˬ��rr���]���7�H�o)&~�k4�zq�V�F(g^�!2�ro����ۋ��Z����
N�>����m��ӻ�0�.ش�F��ء��c��o�-�R��y�6l:�!7&t��&���������S��Ǔy;ջ��{��aj=�U8K���S�򊇢N99X6���u�#s���)nJ?��O�]�zv�kιW����ӹ�KY�.��^6kM��^�%h���v�����Ł�K�G�Y�T�u�Q���rsNC��&F|���6����]m�`��]bPM	t)�ˍ3�Q��<xl�М��L�L�F&����,ܬU��S�5.�w(��}��4@��卩��AY����5��3��P�WE�ݴ�e6P�SKS`��Kd챘L�I6�i{B'^Č[.�u�h%w��dٙm<�ܶ��{�۳������������3M\�jM��qڼ�"�;�'3St�
���ђhi\STqS��nim�6��ેx[[���ݢvm��+��Ao�_;�ʒ������GL��6�:���,��Y���v��B�!�`�3x�[s� D
�ް߃�	w�PA��OK�ϠC,E�#�)�]X���{����5���B �����G DL�h!ס|8 8�+�r�!"���
�F�C�(�����[�E	a�����L$nX&l|LR+��M�n��QU���S���嶾����e����ÃjΘ{pc*��y�����L�P�k�*/�6oeDc���]a��)%���(�B!��_u�5�yr�:��^�n���Y���V�y��0�huȅ�W��\��
���YCl*"�']�ņ�q6[�J�
�-#k.�#Y֭N.d�-�!�2����)Sz����C��T�Ƨ�7�Y��m���̺nDw$f�[8�quRU`\��i6g��L@��戵v�	uR���yB�c�n�*V��izs�Шӊ��m�/*�K�����
��wW�YѬs���g���tjOnB�ݝ�<s�޶e��u׀�SyF�-^�/hDR��fePL'x��Iv��9E�T*ŭ&��c1�&쪀�E=0���m��3e!�۱+������TG���.�����;���j�W��e�7R��xڡ{�|�\�NL7��Y*J��y�gq��C��lh����W���U��8���p���F����5Wjڜ�d3J��Ԓ�/�-��eH��(���Q͢���Bn�Oҷ�Orҥ2�,Eb�}�n1<4&ިq�ܼ�.m��j�\�͓)�V�I˸��ܫpᳰL[Y����)��S��hX��CX��X�@�C�m�.��{pR�6�f�M=ޥYsMRږ��jU�v?{�ŃR5�ه�+��{���_���_)�����/��~wy����; �o}ux��x�}�{��jw�[��;>0����Ŕ�3R>����w6�<:��Ѳ��x�u~W�~W�}���|h�A^6���X���W"M#i�t�M;8pÇ���7m��ծk�	|�׋���ݣb5���ֵm���X�Ύό0��_~�К���\����^3�5�ӂ+��{sSҚ>;8p���{V��U�X�}�Ƨ޸l^ڽx��h�2Y(ީ]^k�}�za�Ֆ}��aUT�,��մ*ڵ-���X�4h�Ç�|�������W}u�k��MŨ������� ����I�g2Fؤ�6-��Y"�$_jۭ��ǚBH�!��v�v�2�+:Z�1��l��R9m���s
�!HA.'9�F�W^�eu� A�n�~��K���b�J[s>���U� ����U$X��O0ZnDθ
4��W�t�`C̰	u�]�'wd��74D��@���^�}��-Ť~�1�㜆�
��Q�[/�=����칸k�U�c�LH\�k�e�
�XX�o,��x�v\�ڧ ���6/cֲ*�ͽ]��!���]������Ͷ�E�2��| ����KΦj����h��\k)w`{9�� \����΀��v)��GdB+��y`;}9�#�&;��8�,쳋br��0����E2�lX� &�Y��wT�m�2�N��cU�]�N���4�/qz��G�c��ofcf�\J��ԯ(dN���u��ׯ�{��!�
�Zp� U�V,w�(-��P�VЂ�귗��|�n���!��T�ݰ)<G��tv}�J�3��IE�g�<)�VTK�B�������o��d�r�mlb��ݓ�[�u}.uq�#��.a�\z�{1^�3���Zu͗�.�z�ޞ��r��8p���G^�t�Nթ|��VtbnZ�:�%�̽�yW8[iҽμ4�S��Z�ӳ�iA�d�̓͜����\���O�-2�����}�ߜ��~9�,�~��r#��%+9%Rҋ ljܥB9�{�e��{�0~:�}w<7֨��s��n�JK�������dFȉt>xo����ԁ��5��E��K�C��Ƅ���r�y�E�$����^xc���}iw��q2P��U�}�[�&5gU���S ΢��fI/\0�9SH����EC�m�m��a�!�U�kv�koEk�[�:F6�2P],3W7��e^-��I�$T{��3qRÒ�q��}s)U>���bV�}XV�l�Q/�7;K6]��"��.؎�X�'�pC�k�����!y��;R��Q���#�+�
�7� 5�ׅ��*Qx;F���!��,d��5�]ߣ��`Q�W%6E��U|=�sX���*�l��ĻY��|� ��r��b���.�z�i�W���S�U��z�&��v��������1��"���0��U���%O]�"��e�bZ{z�\�������u�A�wXj�)��/줦���窳i$.��J�ف��B.��|�-�1����cV�0�Y���]�f1����c�g1 ���ŋ��ִ�����ҹ.���T�ޠ������{Ʉ4��i��T��2����&YI��4	{0)w<��4�R�v C*1��$��/ 
��@���;xv�S�:��N�}Q`,�<yn�3��žx�q�c����F��e�:<�dGoY3�����8{	�Xы�3Fl��bnMW�5�哯�fEx�p��Y}�ib�r��_�{�_-��6���g̟f���@L+�D�dn14��J�~�ؕ�������u�[� F1�v���$Z�oO���u�k��@�������[�T����M'����
�A��Kp]������^�"$��nͿdѩ.ջ>Hܘ23Ձ�����t@/��~�7��t��rV���v�o`��)���o����խl�CvKv�N���T��wW�h�m����H���ܖ��)�qS�P�zeq��Z��/U^�?�Z�uX$�/u���Ucki�!�7Y:1Q���tg����`��ʉ���y�521�"T dK>J����S���Pċ�W3Ö�o3/��]-J�1�`�xΘ0��3�:9�s��솟:YX0@���  |� ; !���M=�o3@�F�G���� ��Z��-u�m�͉�e�T��n'[ �r�N���{d�s�q�s�.��z^ܵ&�w[���W�s֊\ ���p-��L(oo��i�&�Sv���ƀ�|�MC80`�z�#��nT��g2�h����k��v�5���j�EҮ�ݷgH���� ��O�w�=��@��O���/��VD�멥����@x��_m�ي��r��X�\7��_n�Q�		#�����	w˝	��J8�;��[�Ӓ���ާ�k��ok����S�q�ri�i��X6��v&�ŊޘF��v�"������,�]\��)��6�l.��*�;���HBzī=)�n����i� ���9�.>Y8�Մn�Ĉ�oA��涂�)�qДq,x0�d��N�vhӂ+Sb-,�,����_Uv�|���1�U�s�];c��ސM��v�7��Av��*B��{�9�俹k�����jdum��Mͻ�.���JT��y��8��n)C~�E�el���8���뮵��ȴ��ZZ����S�g��	��V���$���JOۦ��ٷY�Ǘ[r"����=�c��:����qw�D��=��)P+vyXf��[�����Mn�m����/3-��%)l+D�H�L�z;w{��
7�&�@� ��E��>�w+hOm���ǎ!R��@g�u�kc���E���hFp���s	��O�ހ���w��^�zn�K�CnDF����5 �66��<��ͱ�<ˁ� ��j�Y�v�p��	�׋O�������c6��=�����<��ҫ�Z��	��UwҊ�������*�n(�,~�����}�,����k���d�psHujD��/��Y9>c�4T���x��8*i^�z7� E{�����a�[`b��ľ�}	^�I��{H��ҭ3��ٙUa�1�����SW��'�n���0�<w�6셪�-ie|�ͳ�G������O'�ᅵ��p�.1ҵ��kԡM���gR�v�R���:�uz���t�E�ii��j��������y�
�I5�j��m���|46=�8`ʥ�k��2��;)f�l��4���D�nV{@��E�(��+�!v�U^x�����z���H�i~2l� 7�����ᘖl��7D��	޳�U�ڹ�
@�!��4S�y6m��1����o^\�wky5�|��Uꝕ�f�X��_/L^#�󐖫�!W�O�X������p��젖�{7����������3��w'>z~�{#��kW���K�fvc�sgA,��}��A@��]Jkcs�@yC�Y+y��s25Uή]l�;e����� 
zì�+S.�z���֎��W}ZwͼGT@�ΐ)#����'um����0?��Ik�z��5k���~ԅt����|z>��w�)dZ��[^vc���+��k%�u\�jۣ4��7V��UěX���f6��J��u*/�j��6�N�f5���<^�1I
Ȍ/ ��s�R�wf�Υy��`7�Z�i�H�wqކ"b��%R�'w�Xb�e���LᕺWr �{뭿斋ƍR�������u���߱n�AO
p$�/%�y�~ϯ�`g��v����nPXe�9P��<�gi>��Ĵe�}޸c��-^ e�S���q'лb��$qܾ2���ێV�o�3 g}Gj�T��a�+�K�z7 {� Ӆ}J�R���]gKǝ���˴�gg�7W�a��_<AP+��a�jhy�{M����iBg{oj��	�5'���l���~Q,t�{�/<���3}�݄F*������j<A��;o�g�n'���M�墭ZOӝˀ� P.N�s����U�I�c��`��e�݉�RFh��,��m6Ľ<��bc˔W���t/j�&�H��7ў�s��\�I�|���"Dy��;�\q��i^T���/g$�ew\es����0�T�bz���VH�JB7oٓ���E�|��A��-Dcr=����t�Kb��n�ܧq; ���[U0��
�J�D��X&�����,n�yα	�v��Q���8q]N8��xh�n�׍>�bu�&G������*����f�5f3ER�]�{E�r�3eM�X�����A ����lEUjĆ��F����\�	&iY��(���t����а�U�O=æm���O=0Ĝ��+9��6p�\�n.�r���ǎġ�D̉I��s/'�e�[��=n`WoLk �3���򹾒�����`�L��>�����᪇3�.��ȞZ�U�wlt[s�̘�Og�q�w/��X!J"cO���8S$��-��:=h���E���度���T5�+I����4�3�j>���w��3�T�Aʝ�VJ\���,;��s��}��ؽ�F��2�Yaa��=�)K39��I��~	gm�+>(�Y	�Z j���\�N9yP{��y�u� 8�ţ>�����;�(b��Pdq��`n����4V՞z��M��3����J���M���N�|���Mij�1o�蓴�N?ӻZA��M�v�\��z)��6+7�.��d�!6��1/BWT�P��dAa���@��'���R}M�m����[7��K^G�YJ��KhU�n0��0E]���>����Sii�6����m?���D�	LV�X@�xvΖ�!�e��n���@��D��kGK}G�7i"����,�`d�/7��l�;�30C򿦯�h��ۨ`�$=�=#I�!������>�hX��C�@M ��\�|ǶJD	�λ�n�X�uβ�y�S��ݡ� ��x��R�� ^%x�5X�m��@�0���2�1�o&$E@
�u�X��}^쑓����#�t=����R����S�5�j�y��hB����OU��W�qw
��䟥�d�x�^oB�i��F������ydD,�'10���S)z��9��=�<��!8�=cz1���ER}�ޮ����0� ��ܣS��ҳ�M=t��/3Us��iP[�����#'�1�g�O�i����1;�6$�;u�N᳛I��1\�{9����}qA3A��C�BאB���W�5�Q����o�I�˙�3B�tj���J�<XL7����>�ge�H�������<��$Ak��vp�it���u[�f�evam�ܐ�b�.r�����J���d4��z4m���m����ΗB�x�$	O��x;_K:��X 3n��!/@U�C�Ca#c���̙�;�jr1��	w���t�T��C����h�!j">=�!{9Q��jm\�X&,�#� @��5�6�D� J��%M�^����@�9,S�"�k�"�ּt`�~/!��1;Q�I�@v)���wg�{"	d�G[d?4
a��so#�<DѨ���T�m�X�N�:
�`w���F�wH(&W��7�b�[��U�8�G�Z������r��F�Y����ά��VށD���)eP�j��'�h��jf�WOMK0C,�2ʕ�^����	��TV=�*��V��g�F��c��T��D�--���h�|�pN8{dF��%e"z�D
�A�pk���yZY�x�2$����=����7�9@����|��ù�wLe����T�j���r�i�8�UJ2�ۮ��h�V����N�U*
���)�tv��kh�JY��6�l��1�m���Wj��.����Lo��뀕2�E�ž=�j����|�2�k	qI��7�ǹ��)�.m���;�)��
��l��;3�����\�c5�+�T
�K.����b�YX�,b�MWI�Ӟul�A��$ڛ�N�Z�ee�mVl��=V"��c�^���m�56�8GuP�H�v����T3���=OL��[�+��Q�{6�^��.*�}��ɱ�C���!��fAfw[ɌyO%�*Y�w�Ɍ����d��u�ލ۝�*��
Y��<!ٽ���H��ʻ��X���>�45-�oz�
�^�U�t�����E�л[q�LK[�T���㊫���&F��.%��fV$�Rq�+]b8]��N�#oJ��+�r�be����_F�����S�Z���Ἢ���4^pU���������fN�ms{d6ԡ|����G��J�2�՚��;6��������d�KV	D�;[��]ո��1.sz�`}%'v�M^�)W�	z:c�*�-O�r]�za���Z�d�qJ�)��"���E�5L�ow6�1G0X"!2X�S*�W�L'7z��Q�v.�"�olMJ\�#��;.�]ܘK�R�Y�g	w��6�W�]0@t�;�a<a�V��$�[�P��b�!PY!`0C2$8��0 �� B�p��2����h��^Ch-�E!`�;�!Lw	�`�%�� �4L�T#ԡ����ݶ�W<EO$����iզ���v�\R��uY1�Y�N�ۈW"jNBceޫn�Q-S��9F�굯��5�n��-Ls�v�k���s�����)�Ye�u���S��1VF�IE��iZ�2��TE$n�>���+)8�$������'�7d+�+]U�������=�ɨS}S�S!�s�Oy�����#T�xL4_nh��z��r��S-Z%m��0Ҏj�٩O�>��r�D�f�Mk:&UgpcuH�e��`�V���R�י���iZ�N��OQ����;�.N��}A3XWCyZ�h�.ѥ���&wh-;o#�9��pZ�6췓��K���ߐ�{p�¾�>�X���o\�w�)�^����b'���V�VV��w&kS�gS�Y�t\Jܫ�T���ompF:��E�G*�4�����ɹt.c����j[ko����i�&�T�$]7J�17{�g����W��z�(�^�A�N�k1Jyq�nݘ��H�%�r�t��a/w
�Q��(���Kw�滏i�9���]�>l�U��\M�Dr^d�^�Z�n0sp�"kԬ�=m�J��M�c�շgM�z�<z�N�:6x�֔��֞;i�m��j��O붕ӊ�oWn8���1�J�o%ME:kS���l$Vd�:�,ބ�a�<�{uW?���	O=��K��d�Z-j�N6a�Ǧ<��-Z��#ysQQ_��4���lk��j����F�<=_k׼mC�\�d����h��\�F$��y����W��_kݽ�B��k����h�b�0e}Z�������Çyc�j��W���k|xƦPbʖ�8|l�������yR�Z�[�(}��*��|v5�6�mKm�-�>4l�����ʽ�F���?F����ۑ��}�C��Q^�������采���ڕbՖԨ��ʋ~�F��!�~.��wW~oryZ���ѳ���T-�T�Z-�T�ڽ��sI���ccTc�z�WKd�r��פj�w��2��FC�H�v�"�I$S��<��vW]*�ͨW#�چT��ڏ_L�V��͖\�ʕӵ@�뗫�|��X�n�L#8�ˡ��J�u|�}��i�Sm��m��V�S��VͫJiM;)��m]�a�AB��:�U��-($�h��R1#>�� 2 d O�h1Yi�����@B eHa�;;0p��3��pϗ�`�[�_�T|<dA���8=>�>�ioi.j���h���˗>���qY`Pt��:'� n��v4�1:��瀚��NWF��:��n=W����ۥZ�
�.ux5��P�֯	㐧t��C����N�gL�J��{��U�*�-��u��\��CU��&�Ѐa
��n�o)wmz"}ۈ���uH~�p@�s�������f�$0�^7WxLb��_Q9��=�h/wt��3��Y)�G�+�qD�D�V�,2C&w^�K�6(�v��F��u��ﵥG�({8Wڤ��d,M�_��;�`������J�vy�1���\_Oꨑ����<���\���@��u	�S^��e����%�*��3���I�~Clt.u��1�F����f�^2�5�mK�no�+���F8.��<r���_	}J�A���V�7��:���X�
"00P����ȷ��nu`�w��;��*�Κ�fu5���k�糽}[��K�f�ލ�)�������
h( H ��g[�GS�Z͙���*�_���wՐǛ@v@wN� ���^�9�Ն��g�y����P��Hs��.Qv� m��m �o:Ԏ�EI�{i�
|Al+$wT,��u����1-���n\�'�T檨�W��w�]�I�(�m�ҭ�d��ueHo���_f.zM�ꥴ��(:��8|(Y)g���� ��#Y[����ɦT[s�vU9�#4CΪ�����>E]���!b�]�s�^v�b=R�{|T����y@`��!�}SbWD�*J�v��$����'��d���T{Y��#q�����1i�+9=�N�Kդ�<�f �g��P�l���@� !���
9H���lY�T��;�|u\�p���`= w��א��y�p����Fo�/�Jk�2.��\�:f�O��w^�û����b���j|�B��˴�]Sirz�v��y���'��o���fؿH�g+1Wi����^�j9Q�ە���ǩF9�O(d�#$j���P��s�J��!���3��7�Y{{2n�`�,&S�������v��0�$�>�,��S�)"�:�����7�@�c�c��}s�`��W9��z��BBP(VǩnU��Ѥ#�K�jSt��e����+7_�r�ه��d	�X�c	�0(7�M�0mp�r��ȳݬ�7��"I�j7�O�l/ �" ������ƾ��9����X�	���h���l?���e��wKk�&�v�Q�D�@K"���E	A;N���c_yXhG\�a���5�oH��w� �&X\F�s�&B���NP�7�N�ѤC�\�\#��U~	����)|'�N=���������⍔y	�/fG�ʺ��rv�´@���L�H�H�em(�l|E_�b��5�>:�ͧ(�K���|L��� y���:�FA�}^�^C��>���mL�BL �O�z�h�`4�0� K������k.�;���DY.��D�#.���^5�7��z��q��V��Uͮ�����g>Sr�U�Lѵ�n,��v��$ˠ�E�lN�цMV%]����d�w��օ��w����G�Rj��ӫ��P�J�s�������  �gVɤ��'�)|d?l�v���O�&���Ⱦ;3�����}Z��쵝h�D��Jkgݬ���5��`P��j�F��k�֧�v�/鉍����)��/���1R����e�i���t�9�LV��$���R�;�/�@E�8V����/��W1�;3�O������"L6C�^ ���ex#_�5g��_;�lU)EF�4�t�OH02:M��X`�f��B�l�������S:�br�8�d�L�rn'8��].�k��+���z�G[{$	�b�l�wʱ���,<�8�.�;m.P5�'����;��o�����^nb��ƣ���S��>�*<�;wHf����Z�C��Oͽ��1�OkWq j��������'(iƼ5`UL� ��1w�)=�Vޱ��I&2��qAu8�����әF�ggKݡ�Mec+0��es�����@t{�R�3j�fCp&�Fp @��jHb`K�B�]��뾳g�G��)Q)�z�ʒ��o�q�����q�E�[��b]�Y�f����ݠ�x�4@�����S�F��r�γ���g��Y�����A��i����R��N��U��χd�{ynj	���T��{1��M���=ނG�e�ޛ�@�;,�o�Uzק6�3ﶵ�zI.Y�n�c@��؜f��z�b�<K�6]1Ezd��g|�ۄ��˳��g��ߴ�����cl��BO��>��&����}��AGZ@��Q�<4y��wV˻�`�81nՑgw7��.h8�#;<5gh��-��(܂5�.V��n�6,uTwL.i�˰�:и4^�f�,	�� �Qi�g���⹠4�h5h��q���n垝��ĪZ�9����6tZ��y���v����A1P$ށ���w�ytA��Lܨ|<$nº��i�7Q�i십P�^Lb�`#�����\b�"��&�w�����sM�:�b�������\4f�Rnh����
���kNU��m��
W��=4_}�`�іA
?0���>��v�4��g4г_�q���6��g/oU72.�S�];%���H�^3�A�V�42ӫR `��J@� L|<� `m�4�ߞ���������������
�v)w�>V�CS�ۻ��1���#�\�������v ��uؓ"5�w���Td�:�$��1WMv��d_�� @������x�_��Dj��0f{0�{t�7U��biZ�13�o��d�A�$	5��~�\SH�4��X���p��& xsP�����̇�S���p=�� 3I��)��J��[�<��1+��=Qg��UG����\����1�I��C�eY�\��'��(n����
̪+9��R�ޟ�����D6�=�z���8��C Ϊ��Ǽ�d�Q�"�9�[��W�|!��\Hӑ�>�[�Tǁ X�7�|��[�%?�_V�4����x�e�����V{�S�d�n�Ӏp*��0$Q-X�9�y.�d$o[+�SN�5KN̙6�j�/�o Jb�b�rw��x5�ɍxhm50o��!�h[.P&���h2�F=�PC�I rY�2/T�u`2�x��r��t��T��A�Z���dN�vͲ�u�q*S4�5��	���p���n��ńv��������]�e-E���	ϙ8׭u��\�����JA;���nn��j�%r�J���!�;N���~���>Y��mEMY��U�W'��C�"�p,�V gt^���	�(�v)
��
'��[�;d�b��z�s�?��7��S�}�=�A�@h� n��� w9@�X#��vO��7��5w��X��,@g�3;����m�`f T��5��U���\GQ��D���`ܲ�?_VJ����u'���9����U�m��3K�oD��xB��� �ؔ[��5�Q�_>�vE	��{�a�GG��}	Ĝw1�Z!����;-�v"G�]ߢ�~>�=锵��4���`GS���Ơ(+<���>�6�������%�!�ua�|��U��`Z0�c8��i�/���᭻]5|�W��Š�G����N��f����[��*F*.-��$䋊v�ȵSBc�e���|���0��6{���\�F٫O�M��`"�QɎ�t��Y��Ÿ�X��vEǻs�*��mn��2^',�̏/��ۨF���΋s������� � !�0������w��d��*�=o�bx��M=����P\*��"��\�+�{��[א�b��Bqcmtn�"�6=���nʯjիY�e=��������@��{�׾&���H&����ڽ{2�r�نR���;Z�f�11�t��Wb��X4�.,��8�Q������޲OYZ� ��[-�� L7��c�%�� �dC�d0����n�4�
�>'4��S�@��8!Xz�"#}����5���[��b�Y�i�%P�j�N4g��˙���y�j��T��Uٱ2y�[rtb��/��u�f���(h�)J#(�n��ʲ�-٠*��p��|��m�e�w���xٚWbx���5 ��P� 0��^�H���Vg���7�o�W�s�_�۫��WuK�5C/�l���A	=KwKXr�k�or�7���w�ee�C�P��WU:Ft�SD�u����z+�/��^S!H�z0+#[�]�|��N�Lf��ͭ�D�ám�/�u�[&wj�C`�uK"
�	DS�jA���޼+WX��( D@���S���5�?�$�  υ2c�Dy?����s��a1�NK�o�Ga@s!�����!�����*n�@91RPDK���f�lr��{�����U s��u��:N�ܹ�P+|���ʺ��˝T����k^��Cð��<E%.�;�����2 e6rP�tЂ�kv�����P�T�|�>�6}�7���H���.��]5��h�Xr�Ic�.����.��m:9��:UCTF��ߺ�YF�w�{�k�����JO7�9���r@�%T�L��W�ٓ�J����uRK�����5�7T(`�V6���c��w�$u쾦�8�y��o��0�p���8�VR*0׃<J܃�cf�[�����g)���!^�����_T�{�g͎4I��Dʧg�1xU����޷y�oUY-
�QH~���;���d��w�ml�M]BPD4�X��yd�yK1��.�l�o�9.;Q�"r{�ƎC���#
�,��g�[v��F����T����±N�����+j7Y�9	�V�td֝6��f� ��P��ldA͘-��l@����xS� 0��Ͻ�_6����O��f��A1�\!cN>S�X�5p&n77V:eV4	��*�Vm�%���鮧s��-�q�̸��T�H	�a��Ͼd���Z��ʚ���N�{U����gd�~�_��|�]�@��T1�wG�=�s��m��7C�h<�r�{�C��;�.��_�?���	�z��"�H��h��}�kO�@z���g�,q��UcM���ܟ���s���	~���EB�H�[�����U3�]�p'v�O$�ֶ�xP�T�O�+5{4}#0�ש��{U<��Qo<W����(Ή��>~󔒫c}p0�����ǩ�%�ڻlC,�c��E:�N��@=���( �VMƘ)D���F&�5�\`���Y��ų�[��R���Wx(��{ځFk��ũ��}ORb]d�uݵʍ"݃�:�[JB��HfNnr����xe��YSJt�N�f[��sKu2S4ۆ��.nv�:�Wv��A���TB���Υ�1�+8�Ǳ�Hw]��X�SD�uK��niUU!R����U�t�;�0mM��ps+abΛ�w;8i]�U�1�Y�g7���!щQęؕ�9�=xyp�幃D�nR����mN�_t�̴�:4	��q�*Kw�V���N�#�>"7p�	�����mj�D:1Q�*�hn%��U��YBGY�ۋ��}˃t���ܢC}i��F�eS���	#l��A3MI�ٕ].�Pz�4v�:��{��3C�×Uf��С�V����d���C%_+>����v��q���*+++����e�z�5j ��@���[�k	��b���6֊炧M�#-
��֯3��ud�)E;������Z��Eֻ�獹��y��w������Z��2��ǉ�gV�ڍ�|Sg��u�yԸN����V��m�)T�O�����������KVͳ�r,��r^��v�7.�������Kx�[f�+y���QJ� A�j\)�f�܍�Ć�(\��@�4��_��4`��c7�0��`�7��P
g�>�����"�h�}�a�	���b�!�Bi��mR�}ClU!�w���DU�'��Pi8j�p�H���CX(0���¶}�]�g��|�T1��0�(5� ���}��6�x�2�V�멝+$�s���:.�_���T��5�9(�Xсd������7X[Q� �����Y�^$�p w-��}F�AXv^�}���=�=��*�1I�c�[��vF�^�n�c���e"��� �W�Ҋ���m��!�;�
�1	�Bɶ�ou�Y��r �U���R�ɽ�yGAztj�`�[F�T�a�%5
w6�Y�ӛ%�^��Af�`�;�&/*5��u��ʆ�ɴC;x/2���V���f��mE;T9��V��M���5נ�Z귳!ES�ҡq��퉼�Lmet�a���"ŕ^�q�L�4+͏[�<�3�3�Q��wu{WH3&��kT������;����0��U�S�%�C�~쎔�{�ڮJЂ��5���B��u�9h;Eb�x��S �Q&���OT����Ib$�f�K2�H�3��HMU�ZҨ	C��"�P4toq�mŜ�O�v���{5���[:�/mՆr��۸1�3kN	�����uh,+/\�os�^kଢ1}��e�@���ŭV�H�n�S��j+ �����`Aͱ/��iX������������ZHб�� ō4�,(AB�⣴ڹ���RB�w�|o��2mo�sW��1���ոxhنzp�&w��M�W�7��m�Ž6�h�Il-�Դ�����8a�����Z|�r�i�^��\���r�4��_��vx||x��E���-���5��VM�Ւ-H�O)�p�g<8a�wI�򲆖KP�Ѫ��(�ԵHՇ�xpᇓ�"yd���^�Q��b(��Ƣ��~W<8p�#v*--��j����#��Suh�RwÆΎ�8aϲH�dՍ[dt�j�[$��������
�mܫ�k^U�b�o4��ꅥ��	�uHρ>�96���+X����];4-E����s�JYXe�ٹ�ѧ#d�0Z�t�:�P/%�]�Ys��=���;��1c� �o��	���/��ܯ����[��[+��[⫨�y�׳[���	�q�'�������1��"<�@����G�	��
�+&�)F��	�R�MY[�:�E��Z���5~��mD��io&�_%%��l]YC���f��6�̬�W1�Ԁ�΍��i]w6r���4�ڷU�~��*�{�I7�8%F�>��c��f����_?`�JT`�=�5�o��:��z\T���z�ᰌL���@w�L��-�u��:���2ᾢq/,�@P'f��Ed�����b�U��1?<tG|�\�+3�_ï���uTݗ�L�{X��;�,�(S�?���A+ǭ9��=���B}e�$|JAL����-���ys����*s8��t�`�LB6 *�HFdR7��	��T����ؾ�0��5�
9ݣ7��R��ꍕ��km�|�a���F���t�ryƂ�-�ڋQ[�p�k'Y�N��+�	
@�P�슗�)�X���s��o���w�L��<�xUIQ�یȝ�Ḿ{��U�N�MQ����� a� "�o��s/��e���K�+>"��O�]W�V�
G2�d%mn��S�h�h��X�@+��2Z���B������Q��x1�:��/�� g���r����S�M�w�X���]�D�5�/Y���8v5 [+��+�i���k@��U�pa�kLMb�����M�z��@gM��� o>�ָ�w��m#��rNb�g�im�k>��5M�.�{Նq�ۼHԋ ��d�*�֒:+#{a���MV�Pw�2\X�e(3F��ևz#���	&����Eg6�֜���X���W����Eqp�|*S��@�,�:#`lP��tuF���1����H܅^К �Mh�-���N`�UgUA��KYy��D�V������}��Q�Y�FnD����rg�e�Z|�l5
ĸ̧����Bh��۵���Db���bv�\��j;�I�n\e��
F,�R�i�WZ-m�m
f�R�7e
��Ndtt������Y��	�X��"��d��Gh��m��ڭ��Ӧ�k��  ��#Tk��� 	$���P��J���=�X�b  �#D2\�H��M��뿕��|T��@�Qa�����pm�
gX�]npv: ���9X��)oKuOg 5�@�Ҫ���Ɯ��l8�%i���o����C��� �V�eʇW�#C`�wjO7�m�d��M�j���v�(5�@(�a�L���Nr�f����,<\,{~�K9�ԥ�"�r�t��F�l&�W� +D�ڥ��á%�3XB��bY�iw��9�.^3 ��w��V� y��/X�4x��4ٞ����	�X�z�<*�Ug�9�̱"!�OXOv��!@u/���� � ��=����G��j��.��ޜ�ɸ���^���8p���2\�̖���Uf��y�=�_g�{�g��-lK�����*�=��MJ��d��� (�e�ހ%y��;=�`��yCZn��F����WQ0��B�2���77n��>o���ݞ��\rGq�3T\-���KrpmD�,H��:E0�`�{*�z��������Y��^u��G��Z�[����^`�1�Vq�]\z��O<����\��}ޖfZ����뿒������{MY�e�q
��k�wI�����oB7��jb_˷��j�����#����ʆ��z���\Yżs�/�V�P�okm�
�ұY[ �Du��n@0��*�e_q�˯���G�����c�ށ#�s�Y�r�]��Uɀ�z���{���9pM���֘A�wɅ�ձω��z�	ٳ�[��(�'d�>�T]V#q��o�������e����|��|;"�U��ΌV��e{37Q�`6�{�{�(Dy{��R� {� �(2Jc��Zo`�Ok+6�TT�TZJs$�U'?]=����k��"��2�p��ܛ��KğQ�jW�oq�#�1��E� d2i��,÷�w��q�W�_��V�r�f��p�Z�j=`Vb��־��s1pb��{����s7E	����5SNbz�`t�P툷s]�:Y��;hR癐��hd_l�����.�#��nG�jL�:\T��z*����>�wP+kB�k���mk7�l��
�݂���\*�)&n��b�B����a��$x׾�,
�|��V[����K|��� ���Ec\"|�ol�)��o�o�1����*����Kd]9��vc��{/�'1Q���M��/�9.�Em��q���t%!�$+�vK�5�\bܗ'��� p��N];�c~j�ƛ�ew�-��c��v���{r���0X��!%?;���r3�%\�ٕ�MM��/D��T��i��Fm����6�p�io:Tyk�8��3)i�~��]���n3��/��dũr����������
�:�ŝYu��,�N*�A�;�.gS�k�LC��!���T+KV�N�����C�:Y���s��pf��B�-8�l�Yl����j��[g�VZB�n���l_B�j��t���6m������������{	��W�Rj[���ye�^�Z[Y�u�X�j�˞����qׅn��V��L��&�1�KW��H� �8�	sǤ����� �6�R��%���6�bUft7���l�'�LYTY�wmE���Ϋd������δ���U�3@�?ޔݥߧ��O_�o�&��vo��(�5��dw�[�xjj�x����S�?�Gs�aB����}lp?��5��;=�=�\���5ywh��DF]�43���["�Ha>����p�n�8΂d`o�9b�1(�hk����M0����������I���<��ϒ�%���<�C������0iwXh	F��Ȱ(bg^''���u���6ۄ<��0P������d5r��tݞꙎ^̊f9K%�9�U�dW���x�
�]n�No>�l2���Z�k�ո�����s۵Ο,�%fW���緮n�Z�V�-@d��ϝ&skWw�1�>�ă�R;&):x�p9w�m?��7d���ۨ��>(�{z�B��u�,�o6alPA��PSz5 b�G9�o��"��N&�!�����m����g���
۱U��7�ֲP�S2��4�.��U���N�A~���>�uo����'�ηzWb�P~`1��*�r`�s?!�<��F��G(ɯ���sVo
��4��ظ�t�sx4k!J�w���i�¯�Ój���l���� ��(RI�?�
ؾ\�90B �a&B԰������-AVʤ3bW!��r	<��~J�0�Q� z'"~��
+��t��ٿ���� 1Ŭ���;�N7�Є�kz�������V	���gÑ�JDʺ;%�__�A����3N�\��{�}������jA:���N�a�`60 5�Cyސ��^�_>�y��wӐ�]���QS�ua[�=l�g
����x���4ԡ�n�b�M���Uo��ӗt�f��^��:�}Ѽе�`>;.h�`&6�����|�����wѨ[r��__Kٵ;�/�Cq?�Υ�� .� ѻ�W/8o�ծ�Cm-:sbF	�<����{�� ��0Y��~���ï�	Qo�7%tUL��=�u{�!���� e�|��4ђ9�n{a�����:��Llz�e)�d�$���Xkn��C�P;b�L��`�kk=�B��AV���v.ޥ�c�Y�+
۹B�%GC��Z���W���LmI�6BL�9��֠����L�cfN�*���L�	�Z����˪�������ޞ����@l�+�^�⩜R����m���n�$�х�N(��#�s�Ky�\��7���f�v��>���u��vj�@S�'�d��M绞��r�R�*��M�Jc�"����w�p߹v��][�r��+���a�|�zUC�6���o`c��:�en_ry���,�p�g]5��<ĂX�*�h����te1�Êay%GUh�G���U�urW�u`d��O<dU������F2,z΃L췰�Ud��;`Pȍ2���Gk�u�Ǻ�ϖ[T�6�Fv�SF�y�
�<�z�"��Y	������
l���o%��!�%v�|c缂��h���{=q��J-?h��A;�9�Ȼ�ʋɼ����	iR6�3݌���J����P��B>�I��:&����pB�#Tl�p���T�굠֦K��.J���ǫ�.��p����Rm6�1xH�"ӌ�w�7�m�ۈqM���)�r��N�יv�rԽ�}b�(���d���1[����u��;]ÁP���U�6aR�:C���K}�w�Ep��ܡ���xoj1`J����ꞷ�	ow�����R� ӗB��v�R l�7'Ζ����gv�>֊��E�=�|\Ŝ��>�`r��L8�7| P� ��A��=�L��X�jV�FWf�f)Y��6����=-�Ā�w��pQ���<�B�&t�  �C��p��C�#��%^'�+u}�јv�sI�w�l���y�t5��蝀֣�xf&��	��5��9�op�^�	a3g{r�i*���u\q}-fC�3x�����i��^�0�/+�lZ��˞�	��F�3�7�VYY21[�w6�UCr���\��L���Kqzyצׅ��/z�ܥGH����C�[�Ef�p��׷<���BTW��}<�.��<��!��H���iJ'1׼�OSBS�EĂ)ӏ@���Y'T����RZ"�S�Y4�Z��g�Md|���j���Y�t��99�Q���"M��ѹ�@@�K�/X�1��蘾�k��$�"���Jfv�^bC��	{���e��dUd����=�Xa�l�UzOQ�C��
��������F�n�A��E�[w�"w�i�M��5�E�Z�N���Ru�[ ���.0u?y-�[��^���B�M��I��q���?B�>��}o��v�0�Mj�����Z�}��	���K*Ϋ�>��t�^�K��Q���r�@x�d
�P���j]n�s�Hq�@�^#E,�x��+��k5�q8Bo�Q[ ��
�l�݄G���=�n=��@H�01%}�Z:���L����)']�{;����[{Hk��=��d�nHl� Q����=����SB���!v�N��dv���'|�*1�}�G4'"&�F���K��.6k@�VCj��v��0o7g�'z�b,틱T���Hhܨ�j�Ca�s50iWխ�i� �؎�0�0��sw����������ψ ?| �M���?�z�D��b	 ����ܤ"F����MJ�Q]�N��:$�A4Y�H�@��PY(,BHl���)"B��PT�#[�tP�EI(,C�$HhH�E����BD(*I:����ȐPX$�Ȉ�,I(,�!
�d��A��Ă��
$�PT�((!APB��AAA
�� ��$��,�$��� ��%�%�Q&��6$�����R%��KE����PX�AbE-$�"�č�D��ZJ���*B��)-%��(*H�ZZ*$�Z�����-��<V��PT�Ii$�$�6��i���E��+D��D�$���	�B5B�REI?��S�v;�Ƨ��~��H���Ii$�$��c�9 ���?����{���_��?���.����?�������G�����~����g�g����?���$�����_�x�H�����IeG�~��ܨݍ'?M$�'��?�����?�$��~�����_�=�J5�G�?ڞ���:F�C�O������sHD	)	)PK,$�V��L�I��5S5�k&�e[I�d�̵���V+d�cV-l�[�k�ՍY-�-lkd�ɫ&�M��k)�Ƶ�[�5��ٖ٦���ɫٖٕ�k3V̶Ŭ�ٕ�k)m�ٖٚ�5f�l�٦���f��Ye�S[&���im�����Klʲ��R�-5f����k+fͶjjʚ�R�*[fʳS[4��Ml٫-5���6UJ��jj�kf�Y��mMl���ke�Yf�5�٩��j�6��VS[*j�5���Ml��͚��lԭ���MY5�S[,��[,��-��l��k5d�fU�kd�ɪ�m�Պٲ��*ɭ���[&�KlVɭ����Ƭ�l���lV���k[�[cU���5jƭ�ɶ�m���DKa:J���$�I"+kIkX�QZ�mm���[R[ZKU���k4��m��cmm�2�cUF�ƫ3m����j�m%�"�i���R����� DBZ�@�h-E���&#_�����~b���������#��l�o����I��Q���g}���:MO����=�;,��L�ӟ��u�G�'����u�ӕ I� I�r?|�~��w�t���:�c�7�H�TY?w����ޤ�n.�ǩ�|k��$Ӫp�6��� �K��#�_�� I'�KQ���_������o#�G�Q�����(�\~�j I'�����$��?O#_���d��1�Sݾ��E�_�q?����?���	:�&dvu����$�G��m�����Si9*�r�u��a����~2�	t����&����'����Ώ������������(+$�k.���th��B �������=����
    �P   �  �  (�      (    (
v��%%$JJ�
U%QUE�(���$ R����U	D�R�*��I"P�2P`�┠��J������%�I ��D�%)RT�B�(
� $BE$���.�(�   nj���4ei���]r�UT�������P	�h�I(�j��U@)*��@�Ԙ �{c�[����*��:�:��=p׵A����i���s���f��N��U��nمk��UP����f���ӛ4Y6]�t�4H�A��U*T���5Hלn���kC�Zm��u�M2mt���sWU5����d���#��gr�͙�f�P*�z��*B�I
�n�{�͢g3kL�9�l+[P�6[��P�-;��5��¤]�ª�[l-[4�J
������j�(I�U�AR���@,��e)\��u6�-����R�	kVm�G\�D���,U]ջAm���Z�Z����-��9H�%UP!x�t�Z��]�i��Nk��6�]��Y�aD�U���k�j��h���Ԩ��w@ܸ�Ut�7pT��{�*�R���P� u(,zgN���p�U�W:��'WV�U$T��Ήl6;�ID��]�U).����+�Y�A=ޒ�T"�ET��  ���UU-^�UD��r��T)U;�Q�*UWp��UEEs��P*����UU�;�AUQ��:�T*��uT��$n�"H�J�� �A^  ��I�T�y;�PJm�Jn���e"	+]ln(%�����]бֵ*ٕ�nQ�@�4Z���û��Eԣ�PR�"٪o 燴ĭcn���W..�*@3L5*���D��ˍ*TK:n%Ii�ܻ�T�nG8�B��S8IR��    )@�@�  �S�	�T�I    4i�E? �))*��@��C 2M i����*4b`C@h�тhd�5O� %)R!��` �  � )�S�5=��z��z����6�A� 42JDA4#=&�2#&�220��F�~�_]w�W���Wz֤JDx�5���h�YU�y���ny�V�{�ߘ� ���|޿��� �����QD?`�������B3�_�8q�{�����'����d� A{ `��P��@ ~@�H^��S��r��$H( �9SG�R��Ϸ�� @
���yh��O�?Cx/���s�w�����D�D�x* 3�" ��"��l��X^6W��`%����RM��Dd���Y�[8�i�A�IA�m��$Pi�Q�Z_%�E�15���-���$����|�ưX@���~#�ćŒ>�H�(�i��?Bă��k	L�I�� �Qg�M��?�E'����� C�� �.	�W���ym�@�un"���1K#s�tgv�c'ٰ r��8�N<���I(��1�8��	�EӡO4�7 ���R��nvT&<8�Ŝ3�ೱ��f���}ƌZ�.{HǊw<~�^�G��T_������`6pS7�~c@�5��?&�֥�R�zi�Vld����3�l�9
SY����2��AOٗ?f�}�9�4?�����!���+�cߩ��sQ�^�G���ߦ��n�°�Ç�[�8s��Ű�']-��M[�I�A����kgT��D�F5�犦:��.���Ku,�;�53`�����oD�K�@iX3F1�n��0�*릾(��K�b��V#���
RZ~|�F���z�������t����lj�Z�n2��4���d"��C� V�q�B�ڡ���au�jN1��W�]���g����%�Sc|q���TZ�Fhs��A�&�3�1�3�������3ALِ�v2�>��f��JI��.U�Y��+	t�" ܇��ķQJV��.	� ����T�n
Q����}�( �֚�/k�C#|���i����n/�h�6�hfW$�u;�n��ƾ��;���E<���p��3F���S��/9.�g�g�t���zf�+�h�1�T]�1��T�/4�ΘZ�M*��ʞD�/S�N:��C�l������t�5u��n-{�/U7�c��# $ ���ؔ�y��� '�V�w���u��� ]Qۣ�0�Xojx��M'�wlf��t��#MNZv*&>@|Ԟ"�6"��ۛP���s��0a�9 �{t�ZŻ�X�)��EǑc�K�:�Q㇫ͲX�[��O=��C�Qb|���1��1a�̺<n�&J8mQX������󝙴�4�}��:�qv���(-b1��_�׫v淠H�P؜�D�-��x�bv]�5Մ�{61��J�T�c-9��݈�%.x���K2�U��z���-�,^���{X���=��Yp�؇�<;��~��4��95�2�+�7C��2{����f���od&�]��gw5��b��bAt���ZH���
�I�n������,
3J�V*�tu=j�DG��ܕ�;�L�`*tӝ[���.MC�6�����I�<ʔ�C0�G��h3�Q���4�t����wI:]����r��uצ`�@��;sE@�K�c�H�}��[��]*�e����9]��qf�b�)�n�8�yӊapph��e��f6eɺ!]gqxt�Y�JA�J����g�����9�':�_sԘ@��E���v��vۯ�i�*P��y�d��:���x2��*;]���*��v	L��
�+��<�іI�Wg-��ft�v�x{z
q� \��H[���#�J�e)���#N��6n2�Sٲ�����9-�r��7%�j�z��M���;%��'����=��0������2\c/=��&myA�N�HK��:��>�ۏ�	�K}Bt�+�7�Ȯi-��e? ��?��Lw��?$�{c��2�EKtK\y�E�����X�=�we ,�Y/�����M�H��W���ج�TCt����ߋy�v�����LD˫G��
r���%̄�Qc�iv���4ꣷxDU���:�BqRfs�pi5�?M�q���FzГ�1�������lع��;Kp�r*���K]v�5�t;%g)�/u�X��g�G),��Iv��w\��o͎,k�|��J�s�� �d��T��;�C���f����h��P�
K)�	�+<W4�-d�ݴ�.���Ž&Y�ͨ��ǵ�:P-�F�1�[oT8�u��!�1
��CK��MN
(��/"��NuR�=�^���؃y������x��3t�ze��A�[���i|s����MѸz�!���.��3�\�E��T�(���y��l�O8��j�SC��ꚤ�x�;����]5-��p;�����XiA{D�sI�4R�t���˶�NG��, ���G:i��Y�E�D��NҜ+��R6��@��t��FһS�Y�5bO��r�'�oq�E�(V7�a��]�6˗:زIx.}��=u_	J'(�;:�7�:c�-T�j�����껸.>E�(`�����$6�}��5]L�{5�	�z�[����I/1*yK��aڼ��j��èctk�5˕7v�n��(�G�fj:냻Sx\���&�Ĝ=Ⱦ�$���ܬ�������I���[�qR��^.����U�qS �@[ױ�Lת����>�8��	XvS5m�i�s�1�h�q ̕M��u*��L׺+�Ԯ�R��Y���s�ݗ �l�ûG>�w7OQh$wL�/b,v�9�[o]�Ӵ$�͹�K^A�p�lB�$��Pt��0mh�z��1��wr͛t���^kaic38�$ٓ�����v�������O�݂H^��Ȱ��F���݆�40��f�W�n�8��l��j�Xɗ^d.t�r8
f���,s�����X&��ܚ�"�nj��<��)p�׋�v��.#Z�vdv�[�o3�"f^j^��y>�q��к\q͸f��	.�\No[����-u��Q�>U�~��N��F���W���|SF�zj	S�/|"�ړ�7��4����#u�w�i澥C��ؘ=���tV�,�C-w�f4��^o:u�w�Ga罐�	i�a7��ǅ��,`Zj�7X�;}��_�;�vbA�Zw�G!nyG,x�wX�-�!GuZ:Ew�Ƕ`}��6�F�[5�p���ǖ�3G&�t�)�w�Ss�	Nn����5��o�ɱT��ţ�p���of�έ�f�a<�����X���v�xV<K�='bz>�Ǜ���p�$�)���&�]P�7��$�hg||p(��=Xσu-	Ş:�üW7{�7uPO�1[�4K�!a м�\q���2�隸ns�ބ��:[� ��³��8��#�����on�{�Y���o�a�$� �Y���	�w6�&�p$�:��[͋����q-0�p��(uǛ̹5Ie3F͸K�zK�s{���N���}yYd6�]{�q��;�b�N�!�0�v��Fq�r�콾4��7����H�C
�<����gu�� �鹽t�:r��2��37�we�F�f.K��l��*16���0&�{֟��%��r6iB����]�MY���\CRz/H2���O�V.���ա�nP0����m�p�Q�x�z�8D:��	ɩ�����m�%�+z��c�v�c�m��ˋ4+���n�,8�v���m�/.�HJ�8W,��/I_�����v}�'�r�[���^*;T��T�+*�m�E˰��ЦA�)�"�&��z��h�!�a�FJ�D�b�y�:�1t�;L�k�9�u4]�9��򂝜��d�SIx	I�c�20Λ��㛇E0Ӑ]�i9ӊ�1^Ԅ��rڰgY��E��z��osx��N����]���-�PP�ک��.�%�-�V#t��1�qYe�uS����hٚ#��{c�w5�V6s
-�N�f0C�;k���n���b�ѽt,;����� ��PZ5�K6i�BН��V9����󩆨�䖙��D��{� �=�����v�����8��{0j��x@h����̘Y^��F�0L8��xGo]D��l+~�na�v�3F��8��)��.4;�� ;��5��Ǝ���Ҽ�G#3,x.�q�{��qO�˘w(����	ws�PQ�0o)��뽊�pv�~�����>���M�I^���i¨�,�i|�]�f��Ih���B#���-�׻��s�G���nڦ��e�[hV��Z�k�vڭ`��p�1=��Czx{BC4��7�����l ՈC��n����o��QN�Bnƽ�H���k��'G�x݌`�Ka	�.�Q��@����Wgv.:x��6!��ˠ&������ ��c���"R�\�*P�ݙ0��"��l�۳����n�fr3�Y���/�N-�1��ZB�xY�Z�<�ђq�v������d{��=�'ڪ:��ݶK6�˽d��MK�y�s�F7�a�]d��1TP���h��3d3C�6�6��AM�*����Â��׺�ự��WD�N-yÓ�#�'F������ōg���%����R��t�F��r��g0��w�����D�7;y��elCu%3�f�ø�@���R|v�kN)�e�*��?��1S���9���[����p�[&�Y���=��3pZȎ��k���{��O*(�5�z5^��m4G�q	�����T��Lݥ`��8+
�x�v��%���gp��,Z��Ҫ�k�P�@ZtT%D�8�vo��g^��)qs����:q`�)޽fILzU��e���Y�����#�x�M!������p�wSS�р���%�N#��Z�V\��o՝��qѧ7�M��S�#�w�\�sg],���U�����\T�0%��eL�j��L�5�'�Ŝ�]�z�)�LZ���N &��fL1��8Xs����t�d�^�[+�"a�o��6r�F�Qe"i�H��r��=�L4p#���b�:�b�j*�'P�!wx}6;:6۽�e�j�x�Xcp����:䇳Uܻ���R�t�D`�=8V�J\�i��f���Հ<�ˣ��Z�������)CGk�An�˭30 
4��XGrb\�;3o�m�U��z(F���@�*Vñ�/Mc�(ǷT�G&�����t.9�[��/LLK�L�^;ܪ�DC
���ow�Z$�wڬh�/(u��3���9�dk61�_Cf�y������6Z#�.Rɬu(��u�&n-�ۓC����+w�pڤò$9�%��gP�-s���^u�z�\b��io�*�T{��f+�{�9�#�1�i5t|���;	�������Qy�d#g�Ч=�A�l<��86�8���n9�p6Vn�v&�X)�rb�
ޙK�(`.S����Oçm��u��+�%m�87]�ĪLjD����ޡ����{�}�V���:�d{���,Z�2J��v����M��7_��rk��9%�M|N��0�Q�ug-qi����5���吙��8ɀa�S��kX�x�>�p
����o��u�F��pǸ~���opIX��k7v�V=���^)����B).6��&��M�m�V�6�j�}D޽���\]k�`Mfnwc޴�a���z�{�������eB�:�0�z���9�\-JeW��1��.��%Ahv�}K��XH1uZu�/�S ������\7��n�)�V���8��b'KHai]}�j���9��&��g3�@|�[��;0ݽs�6���q4*�7�L��^wSvv�>c�զA)�Rg\鎆�i5��&�)�}��C�������b@� �>��GiB  e�+�QP����ᦓ,/����'��?21Q��-b,�H��$Q�A��L/�3���m!��� �k�@ �?!�x1�m�c	L��`��`( @��Xc�q�� ��A Đ���_
x��'L��&�%�`e,)����%'�aD����D�E|��1���<d�0<,�Y�_�����������������W�ޣ����zu��T@�=ֺQD��"ֹ�Ay^c�M#�u�ݥ9�����v��Kp1��+.AorU��ZN\���ǫf,����i򘸮]!�|���e\��7�oR�-�Z���f=n���[w��ŏo�b���5�[�nU�6z�{���i^^�{��U������R�T3q������W�^���3��{�����+�y'f�/1��;̠�9I�Y�q� �c�ų�RtF�;me��)��9�k����Rʟzut��wB&���S;�T��s��Vp)�y`(�[�[�Z��慎�ɝk �56 �]�N��|V�]oa��Īm��4��ʗ�A�c͏����{�� &�F�4��Q5%t������VV�7e���Z�ô�!3�Qç-�F���sq��])m���L�F�O*T��c�M�R�g��6��硌S�`��JÚ���CZ�՘�%x���9�+�G1\9����zů�ݫس�}΀�¼��^��
��{[뚇�,�7\=C����u��)*m��!j�"XcAtەiHG9]K��z���p��á��6z�󂤙�pE���<|�z���>�ˉ>wf-���]u���j��y�D�*���g�P�6ķ�>][�Ed�C+�~ʕ��C�L����2vU��|�����c��vx�+�BxK��R�F�j�0��%�ˊn�'Ӗ.��5;�nWm�wMMֵR�1�w4�M������wPD-��>AwSs����s� �M��a	WP�Y�]��F�0�]��Ȭ�yx�=A�{8�6�������iS;`lO����l��-�]��,��WoFjP�m�^p�#���Q�R�ZW)���.�Q7�RP��+�dǵ�qy��(ZR�8�t�s]�g=}�`i!��Fj}�j�gs���'ZSJy�ח7�U#�j���4�xJ�v�b����<��Lfܫ鏳�U�j��͎y�y���|;vd���zo���<�8�[�Vg_:\�
�ݓfm�6GD�J�`Iݗ#�o>�}����ǵ�� �4vI�vn���ې�5+8c�D�;i��q�X�Wb�gT4��-3�����8S_��7ßes�r�5ۖ{72�S���h'n�	Jwd
@�W�zQj=�����f���'���W=�y{�!���Pҫ�B���pg8���y�8�f9�t��ں�P70���Y;�4��J�Cٶ4	�P�d�cyii�{2no�i]�5h~�c�C�#}���nS��d�7�+���]b�mc�qj�Ξti�+9�Ļ+ռOU�'	4��-��4�AL^���V��򲎹��mK�	B��f>�Y�
��2��x��ճKe[U��ɦ���E�c�kw\����7{x�æ�8�N�N�Ca�&��w���z���`�i���R�3�턽˭�HY�i2���Z�Ю�7R'���ܩ�_$J�r���z�R7��nq�<�3���ld�A\��̲tuؒ�k2�ɹ{�h�۸�*kʲ�'�s&���8ۤ���2��7�:��̵ۖ���~8�oqx�W��m�2�V���Q�u!2�뮝�v�������9ָ�I!�gv�Ys�(V��[���5����>ƧZ6&�gN��T� ŕ��޿{úsk�w���o]�{-D���o8ʝWD�%Ma�˂�.��{���=��UY�B�Zʵuz*�
�j��v���
�`��3�}�ʮ��z~ȁH3v�����p�
w5V�vR�*U�]�W�Y��m��sYI7]�6F�BҋT���Ov׳�H��ԃx͐g���;��}x'<�WW���WܭmV�"nY���ngEP��Y7�5����*%5%�*wi���Z��eݩ�y4�괇ϼ�n�>�4��cX\l���)d��p\�#�-=��\T��,&x�7֒�)�ᔰ��!�1�=(�L���Z��j.:ݾ�+�V�ܩٴ^�y�'�Uv�qKm����Bމ=�T�ʼ��^�TA����xm[æu��G��}EKQp�9��q�����
f3�e^��rOP�� [�Y��.�,Ċ1Ǉ*�����=K���x�]٩�-,ݮq�0�h�9i�p�Y�SzK�����;5Md�.�&j�g���-�գM+���ʹdb-JܻGQ����2�ǦJ��GhAvpr1Fx�f\���҇�R_ot��:�'b���}٠d���ɏ��0�i�=^�"Ӻ�"P�*��̾;�E�vXݙOH��Q箷"I夷8�J��[�]���x��t�j�N׸�>	XE�݀���[�����s3���^6hzܷ���g0E��O���<�3����HvE�V{V�Gy�w�۞�-�%k	��9�s��`�}�. 8�<����ދif����;;.��Vf;��Ҥl��3�(����C�[�7d�T돰a:�N�L	�Q��j��E�}�sц�QՂ�f�ؤ�l��osRU�o=F�D)���y�]۠3��/f����k��W9�6uP0|1��+]��.��\���_/2-�E��,9���!�:J�t-���J��(�yÌ�� m�aɄupZ�-�Ο[e�g%=1lY���L�'yݧ�__Dxq+L7{Џ<��1W��[EyU�6�^s�p�����qG8�-KK�53����nh�:�����W:^_�-�1uM���k7�%/���|_L�=�u��Wv^l�jL�Э6�B����W.=xsJȏ}�u��oւ$Ou�׋���i����z����jˠ.��iM��#�N�g��#ślq���L�Kd7�2�T>�	��q�[�A"���	닷�w�b��S����k���|(�s��I(�lWC�W6�z��w]tJ�W=��5_	Y��l���M��1wwc;xƆ�d��g�Qla��J桔�õ2C|]`�l�0���qw)�Ž�_%$c�-c8�5����Z7|h�Z�W[�|<ew�罝|����w�o���dq�Z�ݘ��f�'=��U��f����r�/�>����1ޭ/x��Q�<cc����EQ��i[��P9Z�;pͶ�:�ɼnf�f@ζ7\�ˎ���"���y�>ͬ ���]ҧ5�oʯ*bg��T����%�ǻ8̽KN������<δ��k��!Ix�х������X���l�Q��F5�r��"�{�Q�|����5r^�9�l�|�켵��e�|��%rZE��$$v�WF�V�Ȅ��o�̺���цs�ymN��;���{}N��x�~^Ͳ�^(�5�6��.������Н������|�sn!�}��F�h�8������DO|A�z��WC)J��9+T�h�����Nk�ީ*֞M�7�U�G�;�7��TޫM*��l�'��\&��^�.�6��4ɛ�A�)��с`������~�����ޑީ���͜[���5���b�I���*�B��aoh$h�g�-Ey��&�D�bd�u,T�xR���b�ϔ�{ ��m��-l�^�ʖ���g�s��s�"��̆`����SW-a���ģ3�R[�.�wm�Pd�x�`4��\�8*8�o���5�sNr��u�]~7.nӤN�[8���^��:��|W@�=�UcF�Z.�7�lWi��d󘟥�v�$=Џ��F��[�7}�{�)wH�IP�nz����W�Z�C/z�����LoT�]�:f��d��m	ܯsu���3��^ o��e�ֵ��;+m����Dր�]Zx��mەd�X-aygw�z��L�wL%�<�@2�O�Nq��0���s�g5O{p�y�����G�s����Ö5n��m��<�NŬ�h;YS}:��L͹�Lxx��������������z���U"�{-k��l�ݳ�ę^�y�����ݽ�'�ĈHg�ܓm��W�X�e*tы�M_�T^�t���wn���&�-?F��I {��,�d�K��x��@������BF$���կ7TS5W �)����c�� �Y�k�J�9�5ALj�nt�0o�����v��i~�E��8�^�u8��_[��Yɔ��m�7��K�7�2��O����E��n�Z������o��C8$�8����V�9�/�c��$�a�+��6L���VڵyH��\Y��B�V��q��4t��ݜ�Ó��+�\n`���]�Dr��ܷ���4�f��w�����#j9^x�������7��cg�+�;z�
�ϥ+������*����[�(��Lf|�U����t;)e��м�$<�S=`�ɚ7� Z�yNfL��+-x�.�.M�t�����{�͟y�|�UA�ϧeٴ�5Xr
�s{��}�H{+��b�F������ߵe��oCE��x}��_�˾2j�Q�3�nk�����$�CxG��9ͪu8��
U�r���/����n"Fۢ1��/�ǈI��tZ��1��R�Y����:Y����� 6J�ܦʸjV!P���ae�7�9��ׂ�m�2����Lp�k�mm����n�Hژ���W_�Ż�{u�ud�SR\�7�>�Ί{6ʟ���r(^�#�{Fjor�ڹJ��l��OC�Sc1�iL�����<�`�o B�4�w��s������˰�����o<ۜ����o���8z����j
<���]��Y�'3H�]�k�}�C�[�I�fi�7V��m��|�BR=����ɒ�l;C���rAJ���� �E���k�:�b��|���I�y4�������Lg޼9��;"ʗ�����?/�,�"'�N��s�Ŕ�s�E+ծt{ה�=�/����ύ*��1!������~��f;��3�Q�uao�>��|-<�,�7���ɾ	����d�eP���UH�cS��_�|F�AX���r�����4��n��F{���_J�9CK�c:�'�;��>:��̀��J��u���'��uX�O7���X�U�:Iה�A���|�n,)}�9��zy�끎b�W�0�p�N�
땔3���Z���P �'gs��Ϝ����{��R�;��p�i���q��*��q*�p=Y�y�A?��@\�U���j3#B�"�6�6�L��[�V��#k����@5Ζ�*�0O�_
�r�*�ךIS��wV@+��ke��rw/l4Y��'�Q̍X��p�k@�k��	T
��!�&����}jܼ.oX�N���2��U�	� �F�0( ���G�JXSGK'
[����5��񩢽���7�J7^=�����Y=�d�3�� �:j<��xyT1���u���b|�h�yx;P����N�Px�a���y99$�I$�I$�I$�I$�I$�6&�g��7���I$�I$�9ofv���w%,����&'�8���\{nb]ٿ8x3��4ܮ��.�b	�ގ^u�Z���%�PU�&��NV�mJ�r�6��a�^Y�fp�lr"��f@2�5�峚`ח�5�,!(�t�8L�ݛ��Gz��: d2T}�6��;�d}�4��c�=���Q������)���w���]8�6�$����O$��2�>�& �󙻜�.|���v�"�Ɋs9���)�G����l�\��x�����X���c��%99����	:�.��Z�aè��fԏ>�랏��ϟ����� ����� ��_���v��I .����F��ԶDZoƓ������#ݿ�7�k"�@ό̈́�z�5��E�3|5�[�]h��-ޯ]�B�f�p3wE�L���L�\y���5����C�M|�@oK���x�VR��7������H�^�:6�ȯ+ac)|r��7=�Ư���o���2yS})��t�Q��;��	9{Ӟ��G�{b�yX�[}����8���Um�%z���e :`ףvA�ws��)������'Q��D�I���OUO�[�+��#����P���-+o)�*hUz�N"�n�y��),�,/����>R��UGK�Ѧ=u�=#�v]׿=�qg�9�kC��`%{��o<.xY�b��1�xQ`�5��HMȳ��������A�%�Η��"�	$����ۭ�j�7��
��y`��u�=4��U��W&��$x�3�VZ���=����--��oW�NAV��;��o����i�ܚڲ�:!�s�M��\�+kcŔ+w���R�\򼏺�u�Qʲ��8oo�z�w�C�Һ;��gXU� �mƴXR��,���K<��;iwc��(�p����u�TS�m�u�X2t
޾�ro=[R�A��ZU^n���`���sE�&/zֆ�F�H�o�g.�j��m��L�������޺.���˩��������h��'ڢ�2u#<�z"K<P�w=d8^;��|���Gi���J���Mk=��L�nh�܎���<;����!�kmyVv�{�0���ǽ�v�ܺ���O��croZ�Ҝ4�%��`�����c+�s��8�L�!����uMG{4BӦR�@�����^d�A�5>=Ƿ�0P�T��t��.���WT���5f�����N��p��9ꇷ"c �7&_^���Vg�o/q,y�Ѻ0AtWfD4�>X��\�[��6Q�0�8	ź�t��Ő�e��i���\���Ը�2���Y��Aׂ��>y)jXZ��l��=&�?u�陮p����N@*]��};!ۻa>f4��GV��^�O�H�u��֪4+��+2WJ�ۄ��y��<��
�|B��$$#PӚ7�SS�I��X���%g:19�87��CnyD�법+�����νe�1�;q���Ί{�On�!}�a[T�b�S��,�f�^��˺�qX�&Ѷ���x����켟w"VZ�4�-(���v��%˵ï#J�:vs����6T8l1�Rn�:9��4�����ۛJ����]�j����ʰo��Ǎ�3�/3����ovG��v_wF��`Z�� &Ú�痞����Pb��]O��C��Z|vz��"�zb����%��=uɃ���#��"�5��Z0��c�E�m+��@Գ�T�Qf_�J�p���&���W׍^%��(��\)�R�~���d5���@�&��oL���X�x�6�����I���P�Lw���>�B�gX��:�
����Ii���b�t�ж�CT�nq�$ڔ��.��`��g�Yt�*��g��r�fZ�j��nG�H��r��j�ky�~�6bA�G�
���נ�3^���[35���e#�p�����{�G�B����n��i �3L҉�e��>W��>���p{H{�'|&�yOq5Px���*���q�7E��
��IR��p�w{��}�n XF?b"�=1؞{!@P]��-�Ǽ^{�����Î2k�Ѭ��:� �@a<��f�:��s8����p���&�q���b���Q�>�J� ����s�A �A��<���G�*ң[��,��E3,����=3��mC\��5�eK�}�B(Ay|��^仸��TB���0��n/J�;��r��D�{�i�:�suV�BLɢ"I�
,�Y�)����u�wM)��C2��b�Ģ�ǻƻsd^^��K�Xn�j/�=3W�u3sV��]j��-	p�p߮�t�)ͩ/pS�=�_t{ٴ��f� ��ŝpsC��b5�*䕩l�v���1/S���y��2<��Mo���<J�{�t��<x:���#��j�/�#]���{y�S��<e�$+�;��I�6T௎���G����>������Ϙ�5tۊ/��\H� ���cq�����j�����FT#z��1D�� ���V8�&%t�h���DԹ�q���N+",wO�{��2,�Uyl.��;�G�X�䅇����E{k���mo�nv.`���YF�1��e�E��E�-�<�bf�V�y��}��7g������(f1�>=gr���[Բ�a���Q�}SF�]�@[3e�4�om<aWf���]���1䚽|�t�\>;�a��������O(q�_>�vJ(���x5z��a��S#ضO>�e�Q}���4�f�(�項�0Y����77>Un^Os���m2��_%��fB����u���'�2
H,��U$����v5�-�[�P�dD�s.�tਙ��PV����%]��/.����ͥ�VSM��n�W����-�5Dbd��/#�z8���nB^U2�l$Iӳ+↿��$c��]T�1��5�a�����?%y^W�*i���8ﺝ��z�g<L���`�L�0��㺞:3a\hKQ�0q6�A��!�xLy �cd�������,�/�Ĳ�S*��ͤ�`���eY�E�|"����\7�����z�;ᇟ��)���N@��r��s}�g^�Qzh�<��YђO�F�k��h�j���h80�8@x�A�p��`5m:pɇ�ٱ%$���[���1��:^��F|&F�L�8���g��6^�ƺ��8��)��8ҍ�x5�֦&�c%pfO�0�X]�XA��)����5��Zy������W�:�1����g'j�ݓ&����%ʶy�ۙx��(��;�a���Y�����<w"w�[�H߳�h�rU�>��Wn����?R	܈t���t&�]*�	�v/V��n�S�/���·8M ��L� 42��ȧ���I�܄�^��z�{��Q�̌uv�e���r��&l�BD�������4�{yq��5ݼ��ֳ�Ɩ����>P�n}��w�
�=���&��&JMc�^��k^}�Zt+˦Bp��
ޠ�E�z�b�F]�k�L��Q�P)L��B����n�2u��~�Qg����U��.�l,.2Mc1�$����Y�����Ց���w�sS��CNC�h���P�,rU��7.j�^|8Mђ�`��S�oS7�xϷ-�w���ޝh�t�:��Sl2!�.����&�U@R<��Do��/E��}�����l���C�%�C���瘰�y!���xŻ�^=�N�}����]�q�II���0}���]�ig�
����{�J���Y��@��top&{pRN�6"���T��(�k���[�2;�Ɇ.�0Fb�GbYk���]���@���?��7̋�9�F��6�^���AVK�j��ɛK~�.k�U� *mc*���߻{��Eo�v�޹����ҭ�ˑ��KU$��p�(�Ç��9d���k���!ՙ��5����Y�X\�̑�0���V��������bϻ�R��ٷU����ct	U�:�Ȝ���e�\�x�|@�\���8=tE[9Tm�k4����+�8n�1b��#����X��L�����C������&����fa^�<.��=������W�}1KsO�Q����,�R+x��7���V�`o%W��j}����橘�Tj�>�W��I�E�u,W��g{s3��6��s��삆i���������fU�y2rɾ��2O�z�N�
���X`d��L'ٽ�!H]
y|Q�+��Ņ���XsB��W*�,�l[�vM��c��o�Ŋb�O��O�vykC\�$0Hȼ���
T�ֺ�G�1��_��q��3��Q��{�f��u�=fp\���)b��Dp����+�S���̵��l������}�~>�2�l��
�0m��|�<����{��Nb	r�a�2�a�"��Z�:Z�h��6�1첬���FC2�k��r��y*��}�?h��=s �1F��O�d�ݜz�Y�[sp�2�:^��<��SX�+*u���C츦��(�o������*
6iW�fA�'y�w�s�g!�Ʈ���
FcX�\��J3�-Q�h���]���"�c�.2��[�O@���	�q,��+2̧�D��;�bE�>".G�%U$FER>]�}_e�G� 1���[���& Qk� �0��O*��5?.�'�՜�ˋ9�_���f��~��Y�HՁ8�k�פv���nW��!ध�	����X��ċEfy�1�z[)�gi�nx=��m�%��^��I��K>�Z�j����y[F� Ί�ZR�N�K�g�wl�Ɠ�s���v;�.�`���1�@
�<-��YN�6
���/6����y4��H���0��p��/R�,9�پ6��T���{��z�P�{�ါ��8��鷺�u�Ci#ozX��V\>g+� <�$��IT(p_ �i����qK9�Pb{7h�i�3Ly�f�mÊhǌvu-�8na�`5�W`@�c��y��	�kP���r�C�5u�ז���'�@�s��1�T��/�_e��x�]��Wy;��R�w�$1��<{"�J0Mj���;P���J�l��3ؠy|��B��ݼ̭ovM���8�X�5,m="vC��q��ŗA�L�Y-����6��e���Z�`�U�_J�=.���C�7:���
�x8.���n��t	�$Q�k:Ou7 Ά�<R%���bת�^�c1�)(�ե��ɴ0Y���bU�"�9��+]= �����&�_�ڏ�����Jց����8g�q0 �>�����]!8׈�m�4�h��і���N%2w7����u����ڤ�O��뱼#C& ���(ɻ6��GX"��]�م^�kt�U=�l���1������d����|�s�W��,/�_U|�c��Z=�ɸ�_=�l�������gt�͞k����n���W]Ы�x=߁YI�هYr7�PL<�*�BNw5Fh7��zK���+A������H�^8�uIs���]�,�������;����>ֈ�D���v/�d(��|cW�;��L���×:�-co�8 	�6=�Fg��D�Z�}l[����th�XD�:�#��O<�{!�v��Wg$�ᕲ�C�˛+:�JaN'��ڎ���>���ɉ:���x,�Τ2�zo�Ur���ɇꦖ��RYaڱxZCGi[�m��6�r�-�A˭a.l�>6l��<b�'��m��٪��b�F�YF!W6{�����9gA��$D�0��׮�a67l����K�ri�Eu�z��u���!�d���/�|4�`ȜYm��[۝�(r�㿍o���n����7�z{�<��{� �IU{����Αk<a�%��W����Sy�uw�"�\D$��e^|�6�BY�L�Ȼ ~g�Py<7�B�̀
μ�bZ��!�a�\Z�*�Y�9�3���wA��֖Q;A�[��5R��|�=i�����>�U�@�)���H�� ����2���EB*"Fl	�(q�� �(�E���L��h���p��,%�m��E���e�+��D�q�N&16p'�����"U�<�D�Q?��d�9o2�2#��y)�~`:�8���C,�1�VQ����B�K��t~�PAuaY.�m���ɯ~�7����.���a�ݼ��Y�&i9S"ڰmok�H/+'���pg؏��W�[�~㺹i^fu+��;P�����LzL761],�Ǥ簿�v�6]��F�W��:�m�f��TV*�)ܻ�rְ��V�e}_�e�Y�G�PZZ/*�K2e��db���VPJ�]nQ�u���an�L֤�u��uZ&��Е�o�r������0�e�u2�8�S"���>{2`��弜�]�3�0�L歁'S�B��p�kw��YG����[�=s�r�e][D��ʦ;x�I���˥w35$2��]�v�$1�Kg`9��d�ck~��[[R��>5���{�EM|'}�v`�V�:H�i�,mӭW���Gv���х�ǹ7V�6`�^�2�u\ �f~�ջ��e�a���^��w�즔{�$=��׍�Ͼ���ߞ_o��(x�������h�hR$(�(R��^�)F�)ZB�i��&�F��)�)��h4��r��!�%�fH�!�&���j�1�T�qI!�DDDA0,C�SDIAFeĴ�CA�	HD��(��&(&���b(��C�
(g4��D�K13@R�)&�!�
R!��6�4��E4%&�	�&
�j4�I1!ED�A2ČJēQ�-$RA6��USQ�����
���IDEQRL�3�L�S4̳�@@TIILZT�b0P��CO������A1$4T2U:ր��4TN�LDTS���Q�5�(���d�P���PQ���(i���*��B� �
)
i<ZT�i�BT4�,DB�=�^�oo��U�[s��1�[���mx.�żq��as�LS����Mv^p�[yڸVc�.�#�z(��_r\�]o�?���k��U-������E3��0��x ўg*ƴ�����*f^WT�wl�s���;9"lB#�0y}ƺ	U�
��HFn@� �+�R�@�=�K��#;���5�x���F(���t�����B�w�ů��ޘ��;LX/븞Փ[(�>\]D���Y{����HGb���e_M�(��z"'�g
���oݕ-d�<kQ@!����#����g��(���o�U)N�-�&�3��gWu�/"�8��K ��z�����=�>f/q�[š~���S�I*4�#O�=L���*��G 7���])`_�^��>F�T�=Wodԝs��K�֠��'�6wa�����˄A��,
�2rY��R�oڵ�j�m����G��#�)�U����G�l�����ڧ7�<?O�73��1b��Xb�T�	�goo]#S�i�n�bVP�P��F����Kt�/%�m�@���XxE���gc������y7]=��\��4vթw�P<���t����˷��3�`���m��!�v��Q���ٹ�ѐ_jK}�҇��v'���K������A�� ���Ф~��)D��^��kjq�n��h*���*�$��b�0�gE�q��3��/���38�bˬ{0D��!�)E�hϣ�'���e��[.��z�m0�x���s�(�f�j�[p�un]jNK��!Q���37�/�����i�W�Pr�0�n/7�i�����Ψ�1b�#�׋l$�Έ��QE70�VV�<0a*�l1����:_�>��E��O\A����\����$ ��O\`�Y�DP!��0�H�`�i���3[͝Q"(�0�a�G��p��蒑�$�U��� S��@�I鷺��g*��&
6d���QEq�:U���+菺� O����9LM\e�����wo�RF1+���I��ç��Q��tG>H�"�F\�s}=[8�#�f�:A��'�Q{~A�]��C���n i$?��H�"M���%����z�$=�Nv����1�4Ӻ�xn����8uǬk�����VS[��71'н���.n�$�OL�ӑ[�:�̫�	�̃z�L
�o4��o8��;�?p��j,[�ē����}\Q7`��|ix�����7ꎰ���:�<�XQ'w�
�n$��b�+T�>��X/���E�nn�zU�F"C�U�r�m}�e�p�w�d}��d�z ��gD�Z���}uQ�h3�ɠ!����5�z{�B��3�=I]Ċ���Ĉ�.���î4�+�A�z���t�[��W�:�3��ɽ�uh�Z�6����i�U�p?u,�3�Ŋ�T,p�W�c�w/b��ލ<;�[��Þ�w�r�=��P)�J��E;�ZGٖ+ W�9;�W�ĻD��m4��� �ծ����,�ZN���}%��A��%��~�3�	H}�=k�G���*�][W�\����J�H0sb��͐�jdTK羱u׻]���Nv=��𛞚��G,���IY�z4�G������\#�K�8N��MO�ǅS��Y:�eQw�*���S>�p���*�f����x�dǂ�F�TC��$�����h^n���^�hܴ������s����*��0�h��P�������V�5��e�A��%�S�����(,�Fk��u(�	\s�1WZu4�)l�Fy�╀�"��61"� ���w�L���(�JvԀ�tz��X�Wݮ���9�5����n�A4�}~$c0V�,;�����
,H���-�e?{�lM��c��f�����{�a�5�$�ɹ��<��DH��z$9��WKػ�nt8㤑����P��ω���\�ƒa�d
�8�<n�D	�d����Ǜ�Xj��[���l�,�@�*�D�]� !fnA]��k[��:��/7��xP�.�R8%kqu
y9oz'����dVA,��$\�;�������C2��<9������]{�<��;��[Xt&|$:*�k�q=9m����P֊R�`3��4��Ej$c��R/��k�z�~�7�yS�M��qb�fM���w	=hv����E��X����E���c�My}��1��T_Z������d�x�gsU�z2�Q@]:��(W6����{�:�̕{�o��u���I�*�q9��)��Pu*�Z���`���ƻ�GfL�*Np����yyv����W���p��2���МPz[X���ޮ淭�_�˃<����eO�9�}�=0x��!Ŧ6%T�U�Ƙ���pU�x�w�
�Z6�S@��W{��0&��Le�Qg0�̂�*�b����1��Z��6�օ��*c����][f`W2�k�޽Ӊy.~h6��Mj��UV�6�b�7��9�+rmVBᩀjH$ތ�U�5��{XBh�����:LC(؈타MC�v~�px��8�#��A�Fwu�~�6�|�Uz%�=d%Gl@���K�"�~+J�=��'l�\�Z���m'$G@�M����DȄF�g��jF�U�9�&�/ᵼ��:��|�z����0U{}�5�\��p�Vw:Q:�t|��g#���tFo<��X��#�,���>W �i|��xt��`���DDq��Eg���6M���Uv���|R~Y��껡ls�����r�f���!��W�7fr`�<O{tAxD�g i+�S������O��Bb;��n��G�)���˥�_ȗK�jm�a�"�EՅ)]��u�X�S(��)�2G}�;:EY�I�t�#�W��d�FCby������%^�s�=ٜ����Pu��ެ�n��]�撟]�'A2jH7h}M����qbἎ@5#7F9��$�1OI!^"r�OCUu��Ò[�Y��۹Q��|�]���ud���~{>p��X��t�x�3-�䦙��7Y�v�ᘅ�`r��$��ʧ;�F�mtȪ�cw���R�l�����4U��y�ス��8U�j�v����}�0Qk2��Pt�ǿ�fMs��}�=�]�G��&h��A���8��t��]�#�n�<��+8o`ݢ^�3n� �\�⇼i�������|7NK��5yq]u�z8�<W�Z�q�_p��/ �s�y2p�4M}8��cLme8J<:��B��:�ye�����h�o�Q�f��T��^
��'.3)}�9C*o��\��ySu�p�Xc$���m��yF�NA讃f�f�M���Y+�.��5�OM��m�]�F��3��r�8�=s`������L�w!�,��W_�֤4CW0�4�;!q s�nV�ݥ�w9!�#ҧo\Z�,ik�ߞl��P2��RZ����Xrzv����]��l|��WM����ק�o�����@�<��,�ꨩ^8^F��ѳ�jH!���7j���WN�d�4��؃ �wȘ����0(�D�^g��k�����(�Ԟy^��*���N *Ӭ>�v�y�yiܓ�r�^�\��.\4��q����uފ�{>p�(i��C:^%ltG�@xGnѾ޼S�A5py���	�C�,m[�j���z!��H���td��<�
��xl���=Y���Ob�펈]��b��M��_:�c�ґ�t=�x���\W���I�ˡ�z���"¼ք/���0h��dH�e�1:��R�cϻ}v���~��e&�]FG��'1{ ��oD��5���j�����1�����ؗBz����g�l����[�fk���}�[~�h��q��E�It����̀��xL	؆��9[kK�t��0?:YR*�V�w�+Y��Ъ6�a�u����ɓC�����%�5S��.��Zgz��B�5\�߃<�����o��^\gX���d�/$3:�V�gw8;m�o#Z,`Y&��R�D�_��9�j	��mcro�o�G$w`|��ǻY�+f��e>�gbPu�eH��ީ�ڇ���֧��u��mӮ�Ӻu��u0�[���`ލ��s��~�~�C|Gtm�s6����U�p##�B5�.3�0���/D�η�~�^����v����W�\��X&�9�&��!¯�b��~R��P�.����R_4�6Wr¾r�0���(�,�ƉkKԳcI�jU�V�Vx�z���r?/.�y�\��G��*@q��>v8������!�Zl�w{���7)�w���`lG�x_r�Q%���\d�tnH�]�b6B�6{#U!�8R�W;�׹r��"�`+..:5����"�0�핅������ٸ��w^�դ��LZ�$���<k�H)I�7Hd���6z1�5�Ec��������Q���)1ĩ�F
lW���*x�}&o��Aј��^����Qݖ��������2�q%	c_�&H��rf�L�	��܃�"��p2�=k�8�}�p^S��WC!i0�\t����5�8��v�%�Fb�>Pc���_��X��)Dk{�0��{� ��
�����`���v��f��V3��YAc��wq�U�ݵ�h{ ,�ySǲ=1�v�ܧPtM���l��]�Uw�m�!�F��vP�$_��KB���5�3szɾ�c�Ww!�?3Uk�Y|eY{�h����U��p9�U!����� 閔�ڮ0M<7�?i���8���9�H��5��!F�����!QyAqyM����)�ƒt��.7�B���T6����u�<n���O���h�U�BY�IA�&�Sc���sS��-_EF�&�p��1V����M	��ŗP�&�!��V�'mcۻMd9������٭�W��T�\kFx�MT�d쬌�n�#j^�Ucq��Q�Iʛ5)d�b{�ђ�p.?4j��P�ɔ+�]+���Ex���j��E	�2�g �G����T��u��#����REM����϶dڭ�}�;t|2;`
�@�3�y)�0��{�"4��I��%�t�f�rTs����JD��:=���t2d�;b�=.kg�{9T=|�:Żt�V�p���]
���M��_��v��|�����GN�;Q�z��\��Ƹ{f�=<9m�a��Z�f�Xv��6e�L�U
n
�W��5i��B�i6��ԺS�Չ$��t{t�1�܄h�u��Ȝ��ǉ��;_D1�.|�<f���1T&�D��mn����LB������;�GԸ��D��tqE��ϬFd؊�C�y�++9��_A��MI�U�0��9s�G����ltr`t.�rdM��M�	���wt"cdaQ�ƙ�C0����E�X�@w�s�� L�d���J�]SW�'�[�<7B���G!�2���1θp��	|��$!x�� J���(�<{Bz�ZNc�.�>�`���7)��.�����>�(A�p-k+˂�������L�tDh�k�������fg��j��Z�Ǜ�E���oG������7��EC���_�U"B���,@�A3Pk��Ցl���QB�S�AT\6���Sqv�~���z}�����ks� �E��P�.������F����a�-9��L
��W2v�>d���$8�~3/,�8�K>���rr�3���SF�?y�{߫�;��~���=�ߪ��,Di�b,u�!9�հ����b�i���Y#{<��黮�����Io��� 5��+*~��ۓأZu*��Է��`]AW����m�D4���Ǉd����*��j�fT����4����wq%����B��������۫�L�[����]+`|8��7&]!S.����6�%�ի�sa��PU�Ls#��L/*C���y��[�M��M�Zҳ4�I�w	�]��N�mcr�"��
�N9���*&*�?M�����l��ѫ
�d�ݻ4z7�ǵ�1y}�V�ǂR�h�ޚvw ���m�.����1�Gk)�N3A����{Q���ͻW��>���
��蜻(5�G`ծ�n�1�t�ݛC��˗����N���P��;��>E�h�]�5�웎���gY���,�����9Vʙ�r�����Њ�������b��3�t+���=`������Zsy�4����pV:�ԕ�*n�4�\��P�*K������w���!^o'�G����9�y���e<*F���3c��'�w��|0� ���*1\�!��c�:�J|ebys92�r�<�Q��~�'!��
���t���*�p�y��è���|L	i�*8�{�M_Y�5Φ��ɪ��so����������*�N	NBu�W���+7����Y��ı4��Ȼ�j�9�ў/k���wd��F�uYR�sqw>��Ω��Q���X��d���Q4�A�:�TZô$�f,��K㹙�*��t�����&KNan�\� ��*϶����ZPu�X�idc��]GU2����<��s��]P�΀����۱�����J� ��O���F�'��.[Gc���l������p���Ӽ0:5���r���Y�\��i��yhO�E���O���$�c!�{GRT���2��=�8��`��jQ���{���^�w^v��[]7\Y%Y���a�B�%m0����O��X�"��W�[.������7!���w%u���V`�\J��6�p�pVJ�8��/1@�����i���=�o��s���74f��4���i�#S����Spv0p�)FT@����ە`$�Ὅl�7%�iet��9�����FM�R�n�5ê��Y���v.r�䷸�ӊ��9Yڥku5.7'j�W�Rs�/�A��1�r�>�ǝ��y۞<�y�ϟ]u��~�9P�%+H�Kܦ$i�)�Z�hOS��J@����)V�(hi���hF�D<F�(ZD>��{�
R� SPJ�ЁE*�H�p�Q)U��@��U�Sܮ��B��y{;�7^%~'�S�ލ1, ���Ǯ�%�z�+�s��=LW��R俾��l%Qߞqb���=�z�u{����׮�wCͯ�=ψ;�Ѡ���A�M=x�u	{����H�4�#=�|��~�*r���~�����={�z��:��·�{�}랤:���ܞ�r���{���w˪���*��r|�q�㿼C�{Ć�G���#��C���S�w���~� ��>!׿��׻�����變|�����%{���z����_!��<��|�>��}�� ;��N��&�}�r_���9��|���z�����(>F��-R�y�A׽@���[�(X�`3=��(���?Dy����d9>!�r{>��ѡ*��h~A�2:�ν�>G$�:�it��z>��C����>�Ǫ�C�����C��{���xP���ȧ�;`���j���}�Y�c����O�	��y� 5H]8>`��!���y	]��h�%>��q�̽�#�J�!��O'��y}��>����EÅ��~s�LA��`���Wm�|矿}����I�MӜ�����<|�p���>ç������uA׌����-׳�]�Hr���O�9}�BS�]�*_:�uG�	��2.7��f��{��W��&._~�������x=a�������q�%P��w!�)_/O�ABPp���u�4r����4�$�v�����G�䜹�!�|}���̎h;<f��D(P_�Ssf�������t#}���|	�HS��t�^�����v��=p��0��{��r�����̚�'�9=GPx���]��=��o~<x.���߾����h={�S�O�:�C��Ϝ{���=��M�|�#��z�
|K��=G#���y��t�!��!�J�=���;�����_2�y�����A��ߖ��ϝ��o~��}�_p�y}|�9{��_q���N���������~�P�9P}�w�pu	\������R������:{�x��(�0��{�����n�Ȁ>����{}�L�r�˞.�fت��]�yvl��X�\��eY���۠�RG�]��̜6�6�{5�;�;RgS�ھ���a�c;��
�4�Bò�9yR�V�lۉ��n��ʻ�s�c=xeX,1����È���P��lL�Ѹ�7�p<
�;��3VwH����ꫀ����|�����^�C��O�	_d���������~� 9�l�=��y�x>ޮ�)~N��C�|���R�@���o��w���=|=}��}uξ��0��|:��)|�׌�B��������g���=O�=@i^���I�����=ϸܾf.~�ٟ����a�w���,��b�]�"}���>�_ݸg�׼}�͡p��@ig����M%��W���r���D�輩^R����/���޻��՗M[�dz�#>��ҏ�K"��Vh�������N������z�Cr��к��	�ki
ј&���߇���q?
8�j�
�? �2��_&x\A��^H��6	������y�2���0���+)�Tk�GKc6��$�c\wA�?z�yɻ%�<�fe�u�L�����/���4���9 ��ǧ��ڎ�c����W�٫�v%��u������30��s;7HSs�����P�w��s�ݲo<u�vt��9�-Ή�1�tC�����V��r:8�(|}�K"B	��"U;��	6zۣӎ�7�I�}z/bP$Nl�EKX�PL���M��(B�$l�r��8uI�M���3ę��I���WWv�X�p�C`E'9U�9�!D�nj�����w��x���n���k*�Rh��/�g�R�/��'��ߡ����uSO��<���77O�}�%�̽�HQ}O-���0����&6͉<D�7�vny�s�����~��ƨT{��4$�b��"�2��:K�
�;{���k=P��z�{�Q���,�F?r�2����ǋ��u�IolG����������*.���b��z��~�r��6���_��k���ҡe䬃ד�d��V8�A�L��^��$������r��TN����o�ӷ��E�T}���v�WvU2=V��Q�t
'��L��s�{y��k�Es���y}�}7�Żox���K+���6�y�jR�˶)��Q�~Я|b�}������j��k=l@Q�%���K�&��'j6 �BЄr�JS4=z�ծ�P|d�Уo�T�l"'�W4|p������v�60I�S>���w�L�u��o�t��k������\'�>�c�l�Z����J���!k�9��<f�]�Z�����U��U���]O��-p�Ű����76�saG��na3cݶQ�D�Ox�j.�l.E7<�էR�zC����d��s������ANThħ~���������F�S׾8��o6!�<���WGl���u��8v�n����N^S㬨x�q8�P3.-�4P[:Ā�[���w�o~�1L��P�8��;|Gd>�W���0 'q<�ں��J�;˻\�_"��]��]��uy�0��/y����R����U��D�K���w�gc�Vo����_��Y�6�r�Ց�2cԡZ|���'锪�Ԕ���1�S7�c�-��yf=t.�d�z�����۹��_�3s�˚�ӼK���11~@w��S&W��s��
��mԑY��3dw����uU�I>YY��W:C�4`t�3}���M��c\z�?�ҿ��^kVe�X�5�[�b�q�����K��,�#�������r��.W*�z�n-򧓢�����%�<�g����f�zQ�7�1�������X��ţ����~�_��`��m�^��:Vz�-�?b>~ս˲��ۈ^/ֳ�E%����z:	M>��y)�n][�w�s>W�R2�]]Y�/p�����Do=Ү��ڤ����Y�[Hu����|�G_.��?G����|��7.�����xehG�u��9Z�o8�|}ՙ����<��޼Vh��v�9=>���#�_*9wC��T�ey��A��W�q�Pv�Õ��MtdT�1\�1��
-��wf~�[�%iVju蚍N�ؾ�R�F7ǂ�g��fG�������O�t���!�]_F��;̈|/��ì�I�8�gn���b��5r+��|/V�c��R�͸����|#7���0��������T_�����K��[��H�d�����Dč�K�۴��A�U�f��G���vj��Ս��轳ɪ��Y�;N�x�u1׊.}4�ښʭ�ɞ�͈��靋T��A ����\�����韜W�cܦSkg�*�;���+T��@��A��,�s�q4W��x��@{=�G��W{��u+{�ºإIۨ�Y��m����V^���O.�ؘ�%��zk�+v#��{��S���j7ѝ^�އy�t|5y§q'��j��(�&�[��Y1K���'��F?j�NWW���er��L1���ӗ�X��_W]����|�/��k��b�F{k��c��d��{ջ�c�vsW�#�vk��^�K�Z9�@��O:��Ӱ�h=�j���i���-ל��v7�r]@��Q1����K�/1k�sv��7��~�_V����q�tm��ѬL�^	3+���q��W�c�by�^��r���/˱�s����b�f߶FHq�f��C��DGL��]�p�ĺ�V����:'���'k�����Q[I��Ү�:h4d������X=���R��f��P*`"��9��.$�/���c)շ%橱{#!6Ӥ�ݵ��%&�'���M��WPnbK���� O������|�����qa��l{�T�`u�����J��.
��w��*�f��9�h���`!��H���r���Ts�|=bN��W(�~�fn`��-�?@��b��=�V��F�ĝ�Ύ�ng;;�3�����;�9�"o��5�v�xś����[��5�U�ǲ��J�R�D�f!�`Tu`}��]�W��EE�/Y��yp�ݡ�����F4N'�����"��>���zi�0(��J�ݾ��+[؈���T��ȨNYa�.�SѺ'v�A�z|79|�H]?n=��k��f!���hQ1���͙7�5g�^��y�$j]�*�M{[R�����gܮ�h�f�{�mggt[����{һd����dF�B[�0��E垔�;�2��lz�qv|�hϝ{�2�䅙��c\�v�-C�U.�}nP���7]}:h/��L����;�~_��Ot����H��縅֓-C�O<~Ou�ٔ��"�A�����3�ɓ�������� 4�8�\�yp����9������}(;���,�����͝[��rН�k�G_=�쪿����_\�W���H��I���*�z�o���z��7�ٝkS�ss�f6~]swҿ{GG�J�a�bn��:��H�Þ�:9����'�����p*.]�;�?@�7�x����[�o���;��Cۂ�J7\�T^����R��}��!l���{ٯ;����FX��+�zWL���W�9���m�y�d�p�����vd罘���k���}8�t�� ����p9Y]��}���OH�VVw�������S�*=�#U���ؽt�a�/+�'Q��[Q�}����'�cѢ�(�/qP�8�m��,~p�W7����䧚��g�߼�3�R�j�0���R�Җ}**9h��P'�2e�<
�n�J���oo^��닪:�x��q�#s2XtE���X��U����lxe+�n�"����sx�*��1i�8���=�����y)�;�ٜelR�f�y����cא��U�}}xi�.�N�A�{���W�I�^a�,�b��s�Ռ����E���Q��G��rUԪ�ӝ��7����k>�L���G�{ߙN����&�>�MM�����WW�0�xߞ_G[�S��xQ̥�\/:-I7��e�^��rQ}�*7�����=�ޚ^��m-�FS���+��k���*][{Y�����j���w���gb��]����:�N�'���^�m��Yѣ��+��\�z�^�5��B�z�8��\KT\��Q��%�S��+�|����]��}��P�����}�S
�ī��W��)A1�#�=q�[���w�ӝ����ײ������Y/5�Ş�뷢�P��EZ��sj�k�������������V��=����/���ײh������و_sޟ�e9Q�̙��./���<�Ŝe��휘���[W�7�}��b��N��x]Õ)�|vY�e����y�:]��V�^M�*m.��6p2�p��С�en�\��"�8b�]X���-Y���ɲ�'���
����#��[�����^���"�%��ܺ��gy(t�''���S����b�O�������s(K���l�����K��}U�H���C�3
���O����[�.�G��-��Q����B��>�h�2����U:6){յ���:�:�Ww�tΜ�3QPa��ez]u�{�p�7��^T"u�~Γ���oݷ�7�{�J��h���ųU�܇� a��<u��h���nЎ�Y{���7������WW���/�HN�/L�ΏGLY͉<뻠�ߺ�%��yp)�~u�&9F�..93dG{|d��9v^�5op��6�8�?/ﱫy��Pa9
�u�u�}�/s�Z��rau��輈���`������|�t����e����j��&�8
�)��Ibxq��l� ۃ���� {�
__!E_Æ���3�}QP#�,�!��7���_�b���1D�xξ���N�Β_���o�J�2��o���� ���7Fcb�/;e�׳���LU����i�8��>�3E�I��	���9vf��4O���(�Vr�ޮUl��3����s;}pn��k�_hs}��{<{|��̕nG
u�ȷ��)W�H^�AM�ظ�sAj�B��Z5�T�yǞ���c�i��32�\M���T�v��	�:�h��w�T	�\�b��a�*�v��`� ~���(<�@qXǜ�޵�[�����'�]}�)
�r�,~�{�;��԰�
�22�hۡr���'��\#L碳��0�}f�;;e6_V��9ݼ����uw��~Ӗ1�,��$����z�<��evC��"���XB��Z��/�eɷ��-5�f�m�sK�
��s��
f�o���Yu�*��)�t��e]� �=�-^,;.�mKZT�ۋf�F� M�D�u��0d����b�uk\W/O }]��d8�O�儀L��Vw�w�#�xn�P���sQgVV03��I黢�<칕�j~Ե��
�+^N��O\"p�xx��91�=����2���w��m�+7�q�D_�<嵇���1R�١k^Х['Uo�>�" �Dz8$Bq�L�Z���Y�0!��A���7�^0:P��sk=Z�٧)SʰV��o���{w4I���]E^�]Zqw�c�]��2�:ܳ(9�}ݳo^U�B(T�3:[X�'.�FV��l�hJ��yX��5�����̃����#����t�H'5x�\X����t���w������Ű�flHfJ�L��w~r��Ȣ�8��K�+����<�޼�/[c�r��MRŬ��P�2,�u��wº���4E
%���;��?_�j��y�k��VK��ӓ�q��v�s�a�\ꔧ`s��}y����p7�D����3՗��޳M#_���\S:�a�AҤ�Y{|��`�:����=���[$�r�$�hai��ωO[k��$�i�4��u�p�1g�C�3�5e9��5Yt�v���^N�h��Ъ���ú;I�x=��WI��[q�T-E�_l��P�V�a�f�}�JI�9�e���Fq9�B6���NU���-���	�;�M�4�6�ܝ�JlH�V~�Usݽ�G6>��e!��^���j[%mmoӶwz_{�J}���N����WѸ���nz{+(�ުT��d�P:��w�>��c*�@i�_��P��ZB���}�_wP	@4� 4�L@4�+H���hB�h���h(��hJP�a�@�$�SBRUJST4!)܆���$�;���R�4���}�����!��(%�d*�edW�r�#U��Ε˞����S�;��ő���N+]�����U��l�������ﾪ���ƅ�鋜~x����"ꛡMw�����[�i�����y���sF���kM(Z�kӽj����}��>���7(���oj��29�������.����y��J�俭o�n��r�b-t�Hj��Λ?^7+Ӑ��δp�%�����'��M�u�g��Q�U&E�(mKE�a�l@��;1b\ރ&���D5�l_��s�B]i��3{'�T�����R"ՙ�e�x�!W���;6���"�3��J���T`c�8�9��j�;jY�}�6�zow8���jv׳Q�	;��kp��r:��K��y�Y#�����Dn��36buT(:��B�)�����U����)}D�er���m�W�f�U��_B�̎��-����Tj���+�����kL�2+P�R>2�uE�Z��O�۔fܜ����7j3�l�AB�����YF!�̧^)TY]�d�p�X%run�T�˚w\��fP'��<�2�@/�����J֕Pw-�����u�y��}_W�U}]�s���T~�~��*n�(?-a�v�3���㘪�em�K�<��'�hם��u���ru�g!¬���?We�޵�Y_d��_N	�Y������F{�w���W`��Q�{27w=�6�s;�R��W�Up�5�OGM{d����Ó\��~�����Yf2�o���
������ңE�>��lr���7o�Eٴ_�i�~��Z��>��7w5��ۛ�D�w���$R?�1k/����&|�ַ�u{��M/>у�U���=Fԅ����2;9��L�WR�s�v���_�й�34ɾ�r�u׹�3޷G��ɋ�z�F;�1�hX�{��Z����O8�SU�����k*@�4��3��c�)�zɘ���UyJh�� muۡ�BM�7���N�su�F�A�$��nua�&^u��t"�XF��7\ۡ+67�0�ڪ暊[�N��[�\��/U�#O�~���m��|^z͊���{ϽgT�+�������?H<�l�0?�y��$���}O���J�ό\o��C�4�~�S�6�D�%�5�B�֣j<،������z����$��~~�;�ntΌ@�C�]�:t��=���mC�A�UO"��22$<���}�5��jJ�-t���ֱblq۫[���\��}R���1
^=A�d���˵���B����ǒ�C!���-�e�1/\N�uU�����V����U��rM:y���)9���)J�Qފ9��H��o�Qh�w�����T���F������j��X�T�]��&p
��Dz�L�5_ ��m����k~������f�B-�&�EX)̺{s*J�[��{�]��}ls�6�j���S�H���W(��?}�}ǯ*m�yV�B{azf�b�;@id] ,��04��Ч"Ā��x>� ����b"�3�R�mW̸��m��-�O%��h�]�:���Ѵ�w3�2�$��ֲ��6YS�+i�������\jI�:����b�� ^��Į�;��<5߯��nНڌ�/RUժ���o�;�[:�e����6�s�7��C{[�S|�B��O����c�~�w1�o��Q�_U���$Q3��-��5���SwZ^��~�ח#Ǘ\ƪ�>�ke��N:��˖N���#6��z�1GL!��_n�Hr��-D?Wz��_���3��}�r��mv��=�}�z�a_��ܫf��Ȥ��&;�r�z�t{�D���1����'�Q$F�p���꾕���f����O�/�B�B+��ĵ�9��/f�g��n�n}
���yAQ鱖Ʈ�8�};0X�N>�{h%v�㾅���8p^����2�\KE��M鈴��P }r�w
�y�Y`f���(�����'>�Bš��5٧!��<ej2c�tZ���ڷV|�"�;#�k��G>����7��������u}韀�e}Z|��+��#��k!5rJ�9G:�m����2�iJޢ��)*9Fb��C�����������5�[�x����Q��ޟ�:5J_/���ħaa��zl�_�Y׾�\n����G(��N*5'P���oP�/����;�c.�{�A���S��V�=�c:1�G���#yI�9߾��3�6*OC��Eu��k������햑�Z-	X�O1=x�3�s�Sv&wa!�ݸ�ھڌq�־��1^���ǧ����q��J�륶�����k�蹻�ݎ�CU�ݯ�v�u{F��%�/ug8������<��j�z^����2���M���D򱩈������p�Sܫ�΂����~�Z���[�.�`w/v7��OF̮��k}��9pg$����p�i��9�l�:��{�{#�H�!���sݍ�Ã�W����o�|w��~��ΰ��1��U5qU�&�!~1����F��uf�S�2"KW�/�v���Dn �����V�%�ի�雝e��u��4'ط�(CQ5���Z ���5����V��$�M1���j�M^�md��G���>��thI��6w,s�U���ҿ�d�J-_s�UR�v�q��d��}�NT_�Q�q��{�9�T�`�����9�$�F��۪�%vc�^?��B�WF� ỗ67�)L�Rm�v����zK���^��$��~�N{���]�ý+����*}.ƪ�~�=����Zd���bT�7�H-��B�R��R�*ʻ����Z�Ό�`z�இ�n�f�/2�pU}Q=��������1��NL�MA]xj��,�c+����>�AJ����S�j�Oq�/�C���?#I>5�ܹ_� ��.����y|Ì��3;.��*��/\T�9e���������O���Y��ݞ�
�t�W]�Y$NOB�u�n������8~����utι�z�J�����l��~ƽ�ӹl��V��a��k�we�c'�Z�MVlA�2��,ѹ��u�zu^{��5�ck�b��!�rE\�V�MJpٟ�o�<��V.;�V'&�c�2j��2r��4�v���W���U}_WM�������"����^��xS��ټw���{|�{8�w��\t�m6U��Ӻດ�֕�<����-���O�\��<C�=ѝ�go��g\`��c�)�t6�{���<"�_���^�~���>U8�ԩvL*`gl�m������J���q��=޼�T���W*��k�����CW;<��4F?M<��#mT�ܪ6���:�N{��]��8/�ĥ���W/���o4a��lmwX���_ǚ����<|�0�k���I8fr�_G�_���u�Q�R=��=t6���c�{�]i�ݧ����}�����2${{x�w��fK1
�����z�hb#v�p��g%L��kc�{˯b:�{��uf�M7[�Ph�߮0��7���F�)�>������s#�3|�r�N읓;���]}2�<�vzro^q�R<��]�޸�wi�J�=Ԗ *��[|���@��Z,�;�&�WսZq��Gw5�wS\]p��������޳_���������������e�MR.R3.���/�Q�r��;��k0ĭ�]��s�y���\��^�ժ�GqX�+�}�5�K�&J<���/o<��?"~����s�5��+M9��O��Z1*y�!�A�`~�m֭�:-��p�#>���ߟ����UF�U��9�]�L��
�i��u1A���8���R?���-���l�����kY{�ǵ>��g����.¬�����f^!qZ�n-��s��U}��k����D�?z�fĺ��ł�y;�G���Kޢ;��ku��5��QG���=<w��oE�z�9�{�Ԗ��b�7��Qfw!�W+7�S���z��e�Sǋ�}�X�4j�=4��9���f��/ި�������X��nX��s�-P	���mج�3��CdO�ɸ���1b��P����(����non	�`�;���Ǳ{�Jyn{=�ŬO����{o��M4�E���/)�=���Mbb�K9)T��y�p����������J)꒖W䩡�"�����7�l�2 ��2=ܓ��������$��8���|b��:e:��xtS��o�`e*�z�ov������X��Ӧ��u�r�vq=��'o��*؏��f*���;��Ѕ��K+�5-z%3�C7�P�r� 
ޞ+���Qѷ��'���k+.���򁥆�S_,�~l�Ɏ�ka}+W��������U��)x�����.��{�'!1�u#�Sמ���^.ޡ����MڔfY}[�WJ��)�c�M�.�����~��d�?A�z��*V������H��=ImM���9���+��-m��{�JټO��8��q���;!�9���jR����t�S�t�[v��������^�3���q��-���W]��
A���;�E{����Ղ�Ú�>N����k{���T�se�á�S�����o��Qv�E�n�]�؉g�AG�!�����(� 0U�x�1w�-y�%z.�}�U}UT�t�o�rS����Jn>w�)���˽�����8c����܎��~���9�Za�&�mE����nby��_yu�S�1��Vs<�C�F������t�;㶛��U��_�a�J���9����-�Q�����#{� ؈[��X������3���9�g����^�Rk^z�Q�R�w����*O�7*�މ���{7���KpB��z�F�Ωs����b����9s�ϭׇ��r��}��l���͚�=�{��]�_�F�Y���L-��_��r���Z���U`�gO��/DP]R�<&Y���CJe߽���?�������	����,Ur���p])ɩ�e�6z{ON�x�ޱ�0�1ڢ��N̋�s~��w�1v�~�װ�}����<��sv{�>�<�!�473�]��`wl������,F�����Q���+fw�yR���L�tv��[�&����>ͷ�O�W�r.@�/��7�og$�{Vy����0V�
[��Ją�}�*n�BX�~��ػ�!�����Q��̂�ՠ]n��N�3����Sw
��|��!*w�{ZH��=�����6��X͂6�~�`3�҇ݷ���{�&-�vk���bE\o�{zF�xR+v�\.Wj�	6�;s4%�@���i<�D,-��,-�q%]�v����z-y���(�bİ�cXp�F��y��l��S]J����҅�"��⥦Au���v�U޽�=��v?��ܐ7���i�S#�P���}�5Y��M��V6M���Q���N��e�f&�������M����x�Ng�����]i�{�'��p^�\=�.�y/>SE[��/pQѐ��#rp0j@��V��/BI�8h�6�"U���,��n5e�8�d���>��kAx��{��ɑ�^]u(�֩*�Ӗo U��{�6���WѲ�Muy����Sj�E�i��6��h��B�WV
<��l�M�j�n�S����Ƶ%F���W��5��s���9N��K	�9����[�]�Y��L�7����&Tb$�iz��*�#�xu�x5���-��n�v��Tmvs�)�k�˕C�^�f\�t��kJ]�[���Rk�JX�v�Y�J���G�[�m�*.��y���P{�Ml���is������ڮ�k��/8��O�,v����71�q�����n��S�g"��W�ǆ���E����^er/u|�cT�2��<hļK}��!Y�y��{=�޴i��*T<�U)[M�&-F��^��囓����7 �#J����:13�d[�3^��^�vJ��v�
�\͋�P�:��B��wN��*{��-N��?.�2똫�U�|a���$��2	�����C�?����;�%F\{`g �\�f����
����q��*�<
 va��	H�n��6:�q�6j�][bo�1�<�o=�7�mp�Xx֩ܖ��>��WݮN3כ᷽p	�T('�t�d�w�V"
h�$JB���">T*�h(i
�4�a��C�$)X��]&�HP3)��t�4��B�E�(�
P�\��	�)J� "B��A�a4��tQE�	���N�F��ALLU�~}��}����u������Z�=Y}�����3��m+�u{�u�k�I�8.sۮ<q�a�3��������{��S��T�����S�T�f��k����nM��]���[4+\'���.��ۛ�'�[�,�g��!r���W�ϧ뽚�9Td��"�[98��r��z��og�o��$�����8ey�V�^�u)s�"}�I�IdK����ZUQ��ѷ�q7;�d���B�~	��D��;W�_O5���WVX�y<.��t�m,7i@~b��l�S�3��l�E�x[��~3����ݎ#���z��!���M���gc>�3Z���<#�r���xg���Lu�f������^Ag(G4��2��y~}� {���Dڈՙ2��2�O^P�8�Wv���b��2�� �γ�ӣ|��w0&�S�;��k�;���.�g�k�S�4�<Ԭ�(�D'�E����H�qa�7]�-���L�3���콐t�z/+����Ô�vCX�*
�{:�3�S��-:n���C4��b�]+�1=�I������S[�܍ʯ/� VD�?��3�/_�OV5p1qX�E�U&��vEwI��'�Ns��뜽A��t�;)��'嗢��샩�-ϫZ��^9�~��+���>�x�}x�go���]Yw�^�liUu�������:G����]O6 M6*���[�z�@%��i@e?+1��3h}�{�])uC��8H@{wT�nFj�W���+c���T�c��x������>���o������\+Pȳ�,U�x@�4/�o��x�}�|eb�����":zIggg�u6�+��o�Cc�m����5�K��ig�mž��sw��w=���H��]y��G���uZ��h\}>�҈ܢ�{//��ؔã�����]@/r��@0�ߕ^�/޵�S���7X�o"f�q�N�GI��H�[}��'C'�ۏID���ۍ�=��S��):�56q��>�1���7��'Is�.�;-FF����b��u�8�SwI�N�<�Fv))�c��CU��tK��YFּ��ea2�NIo�����꩔��:�k^�FEZ_�]�����L�����\m#�A(�9ᧇ_�G�0'�U�7=��Y�8l�yJ�����w�Ri��JGnIb�����od-��wT��x�L�7x��0���_n�=f��Dn�pg�.s��������2��f�t�í�w�T���.wPّ}˶��PPb5Jݞ��1!n.9F��N9O��ļ�e�%_I�9�����զ}�������A$.�s��;��*=^J5z^�
9(���5/'eZ��r۞�3V=�o�{:L �}]E��D�a9e�%� �P�u��&�8t��f"�/M5x�)G�����otu�D?c�P��]�S�<K�ԯ<��d�!i�:���KޯH���D��x3�OuR���~J�l��4�#��/r�ʦ;Q�M<���7LF��@0{9�q}t��%X��<v�����j���h�SZ�u�ٯ�9�S�C�8�rz���ﾪ���1?{����*��+�J����w�:����JD��ˏ�[GyxG˱��
�ڔ��ll��p+��^���85���]�s`;U�o��jGT޷\aVnG��M�࿥�t���O�o�����_�aB5�����PyH%��.�0�ן����R���׫�{�ڥ�w�{L��_�&�)�.��.��@��mg�Ƴ>���=�޳�k�ժM{l5w��k���z:CV�B�sү�0etV_6�S����[�]mx�����{<z��_�s�г󫧔�+��Ӧ�{j&Vy���'zƈE�#�}����w�S���B�ظiJ��0"~pc�	}}���j�]зoTM��hA¡yz �i�6#����]<��S~��;|q�LE�WCnnLdFh��]5}M8��l��r�����v�,Z�s�{k�tK�Q���m�\<�.��rp���Bb�}bM��p詓��ö�̶-O���}s�΢�a�J�:C�/���r�J֭h�RO�O��UU}C/��FҼ�(���1n�N����������kQna���q����P6�`��/���bFJ�˪L˨L�2L��{5�����Tg�*���S����Fz���'�`�7&��Q�E�ʥՆ�1�Y�Qc
��y�J^ъ��Ƭ�F�u��2?A���i�]Ak��K�,�]z��_*�is=�Q잂|oj-��n]�<��tw�6��}�a����.7����ұu(���@�8c��ҿ.�а{������������'ĉ��͑oo�wf*����}���u�򣷣����.<�2����:Obñ|"N��v7��.<��e�v�y+��S�r��a���ʹ���g�A��z��&��qz��w}�ϸ�1=��[�]Nm�b+c�����(����61�ᢏTw�N+�6����mIɽ�{xRb5�6���x�3%��,�7(����1��
��B�E�I�#N��|Ӝ��UUWvH�y	�ynV�}��Ƥ�]��C�w�{��}[cy'�z�v\>�yP��t��r�ܱ�y��� >���C��"u<���~�!���=��;QͿ�7-�>0��������}�� �o�t����Vm���}�i��\����~���Or��u���^������޻��~���������5��[^1ԅ��sj$����jDs�m3(��l��}�MI+7��m��p��Ͻ��)y��s�h��WCL�Ǽ-���\'�ұ�-ze.ܕ�5�Nu��L���w�y˽����R��]jG����^�f*��ځ������{bՏ�J���q�;Q��#Ξ��GSu`�6 @&l*�~A{�����+�ٜ%������W��d��<�:�@�)��R��WtȌ7S.MҊ&��1"��A"�]��!��OR�o-���k
�S�J���3o2��  �x�Fs6�D��]��t���]�g��r�4��f.e܅�6�)�Q{���P����XҪ|��f����͙F�k<���xu1v�j�X���}-dۉ悈o�˃/��fw.OH�(O����b����##���k�r��^���w�-�N��k��>.r����T{]m�⌸6�y/�p;亮�߼��Ù��Ƣ��V7Ѵb�`������ɯuw�
������U�׳Gn��
���Y~̕���Ǜ�K2}�.���yI��T]o�.�v�Y19����54v�;�Y��t�㋳p���$���o�7�വ�U��v2/}�k����h]_�����z��l�F俽Q����"FxB���×����G�7�t}�LG@��	]q�=Ք��c��!Ay�S~H/�^t�{v�Q9����\.l)�U:�:������(��=Cʲ̓a���X��a�ҍ%1��H���z�g���5ӋWo/��f$����޻���K��;�n�W���˙�8t��'I}۹�ˎ\�6�]�}�}���.��Lvc���|�I���5��I̟�6^�Ȫ�;�5.�Y���.��γ��!�m0�hA�ʥ�]	y /ݺ�F�#X/�|w�@��0ꇸ�wݮw����EV�Et��ȭ�X�W�rv,�:�s��߰�7�'�=�����r���]�T{��]�fj뮦C��Q'lԂ����=m�
���J���K۽�]��^�]�Tc�ݹ=�=O��*��1^q|����;�!����������qk>�4��ʎm��Sᓐ�bvȭ��E����v��W/}qI��f����e���:������|��nFb�����jU94�Վu�����<�c��{�wh�gl_9�����w�ޝ��S�wغ��X����T�F�4���1]gay�2c��Edl���X\�J���V��L��U���v������^�û�r��3X�&؊�S�O���s����3�s@j�����(����-�;��ޥ�\�O%����UUnjK<d�E���d��Cj���������u_���~V"�U��!��ux]���h�j�G��{qdP�\��-�V��n���������� ���5���[����P��Wo��PcMoy�I������kn�Px}^�"�c}�b;1Y�n�|�̹H��$��}G�p�F�Y��k�D��9Z�p��/B�}�k�v����T����q�#���V����q*:w�Y�����#7D�d����@�����FK�9sZ�Zc�7�W���p�����j�J�"cp��r�̋��*n��������W"9����m-U�/�/�i�W��-�LF��V�ݾ:Ҫؘ]]�׊9�R�5�*R㚽2=P~Ӯ����_
������ĳ����^#@���7Bʃ([�vY82��Q�j'�!ʀI���E���y#'V����pH��
'\�X���n���$}�k,����x[��+\Pq����Q���m��&�B��!O����q�}=���5�{����t�;��{妓~.l*�M������_��+o��ӽ|z&�g+T���f�b��}�'��Z]�R���x��=��]�د.F�璇ϳX��>�o��3fa�{�s�qE�}�Ʋ+��#�0:|U�ڂֲѳ�����1޼o�ݓ�*��=O������ܶ�=��F�(GY�l��\{8b}{���.F��}���Y��{uz�ddnn�# >C���m[>��{����I
Ru��O��{���̎okUrs�h��I��x�v�;y�G��":鏎���T���Ҟ��pڜ��3�r[�W���S	\N�x�2r+]�J��Q������H���؎{7xr��*8��Nǝ3j�?_�zM��l(�(��$Ia2|L��Df�����`�^4�Ċ!�9�9�B;�7����Ã=G=�Ē.����a/D����Ej6����ս#o�9g<���'�L�^�Ѿ�,)�w�^�v�T�1o:��3����M<1r�GI-{^vM�ULV(^4�ݰ!j������+N�FbU�P�^c��[7s�f�x��PP��v4[j��ð�1R���Y�K���I��'�+�M��#���&��IƷ��<��K��kt`�䡪*��rr{��\>8���RO�o���.<�w��
�z��^Nn��:m���*͏���z}�ݭv{Ҽz��K+z�.��s��g,(�9�T�O�jR��+;c~�l��ew��1M�O�e�z��E�IR����O<0론Co���T�˖(���kY�Q���Օr�i 5��YR�f�k�~��4�dH��.{S������*׸�m�Q��QRw;�(�ݴ[����>Q-�X�9.yK�g��_nS�.J�,`aǅ��[6�k�7�D�s-�B^�m�������LN��mɸ}:U�M�T�tc��H�����/�֍8�w�
=�})��7�-Ի�����s]��6�N��p�q�Xe�W�?Sű�BEC0!�"
(�H$LC@�`�Q0e��-4�澱	�(K�[y�~RVp�x��Nb����7�H}(ƈ����؅��������o*�d�<�[��������z����b�;*8�YpYc���U;�z�ޞf\�{��������_����Ä�m�0��P�[7�+z�s�أu��׻�޴XB77���{�c��rj~��qfG��S޽ͽQ6ߪ��X���o��yyDr�Z�A�Ӱ��n��}$�s�;G3�_[4B���|f�Cx��Nu"�W������Tx�}�9�k�[PӱJRt�s����o�o7,oN���r�cT��:��H\\����;�"������u�R4xi�Ξ=�߱��j���֍�>�2�KC9:�}�!��R���oX���A16錂w�������ǥ���Lg��)��΢:3�;͗�܏�۩�^+gzs��\d��j��lzN-^R���1��Hۻ�C�2��߯�R�7 `z.���}�T�tN�yQ�ѫ<��.�p�'5<f/�%ª�i��U�J�unV�x9W����'Z���%�t�!��%�9�N��t���PV��,f�BQ]��ĩ���������ؤ|ܒ������ל@�y�7%nS0f�8e(�� ٓw~��rr�C��AkiM	�(m�����4Ѧ�@j���V�Ԇ�J�9RS|��l��EW (:
lk.��N#j��)1j�јѣc���������UE�΍h���,�[1��%�!�j��Nc)3�yri�mUo�Д�/6�㙊��>ե
�P!���9�/�|H�O�	�u[���ms����x͝N�qOL�x��t}�nX#��{�u,�L�c��k�Y���k>����)���Uۯz!?�8��d���w_mu_��]��Ef
�=�y���RpG�fVr�����)u�ݸ:zw���%�-�s.u^�f�r�j���,���*5JJV�Gy͕�ч�t�"�32-���bݍ���2�[��j7����^j��D�6�My�K�Q1����՝C�dR��%���tL+�ة? �g�ګ�G��m��ӱ���ٹ}���W��5Vc�p�"r��}kx_m���ֽY��x����h('�k��*<�ٓ}Mz==��<2�����sC1���]4*����,eJ��'|Q��n��&��6?bƋ�~��7ַ�ƃw��~�'��u�|�,�2��eݙ�\
o����+{ba��߫h�ߐ�u����g�j�/�(��Yy�s�=�N��v�\	guH�I��nD���-t��v�4v����݃�K�@����z��u�ڻ�&�'M�Ko���G~�K�u��.�헛�rA̫��[�~�@�Ik������ڿ_i�51ߟ� ��+���"j=�޾��۬S9��q�Z����A��^������ڣ��V�Tvvb?I��!������J�r���=��Y+nӧ�QU�v�e.�.�46,C[C����=m��{�r��7R3�TSxz��Wܰyx,�F��6�"\>s6��x
�4k�(�o�{=�e��f�����5������(�u	��^ڏ���"�{�?~��D���/TN7N�㔺>Q����B1���>9)�ײҍʜ���2��|����7uy=@oW�9�|0�[{&�~;)V�I��y������]�t]�+���}�s��EK�7�֩)T�ƨ���L	i�S��M��D��)_\{�y���v�W%]%������:<ڽyzxYX\���.�,�Z&�צ��1V幛��*<���yC����{̧C�ڕ��h��V��U8���Kt,�t�=Q�1����/y��|�u����V��䶔�:S}�W7�3}���'��c��yU?�ז�t���wN�HƿIK�:{73����Uq���v�yV��o�:����3��Sv�n+�{{Li��]�Blr}��6ǁ��Y<ݛ�d>Pb�R�P�U.�_%Һ����af'�y��9h=�}C�Z�vt��B/�U����&^.������q�}s�,ߌˬq��UK�\9�9�w�'�W����]u#��r1Q�5i�.xǣ�z�"(��jy�u�q�w'�4vEMtW~�C%АL�I�V߫��J��\a@��e���em�n�ם�Á��M�.n�,�/,F�tk�/��Gm�S\q�;���C�Uw��׸^CF�ެ�����D�������	��z��H7�lפz��DA��H�	zH�נ�)�t�	�������;�r²���\��4S��r��n�yz:��y�V�a.����u����$s�87�d�v���V�LuZ�|#�v�����j��rx����^���j���Ʒ�R��qc::��A���?���� �����Y�iw{�u]�}�v*6������Q�t&�M}yx���N]�V�A���<Yا�ѝ�|�[�w��HZ�tQ��Fo+GzE��k�{�\��kt��:v��R�[ldWj�=�	���㵵-37�>3�^f�P�ö]��k�=W�����6x7��lGtT(��Z}aU)ǮR��Gt_��9ss}�!D�y�h�v�զ�����d��v�.F:�ͮk���7��QQ��z�G�㓴v������½^��a<���F|��o��q��iK�E��Ɋ���b���uE?�v^���濺0cJ}����^i}9��x��;7E_mu�;u���,�s�_
W����bW�U���w�"�xs}�����DB��E�e��~=��[KJ�|��53���SIj��o��so]s�Yd}cA�Q��oJ�Q��T��Y]t�c�8!�e��-�XvV%�ղ�����z�#�������=��uH��1��Y�c��'|�q�޾��:�8�=_C�U��]�`���ɸ����*hX�4���YO۰��y��S���Ͷqק��㼭��"Ľ{���#꣒>+��H�N��(x����{�`�%M@���$�%��S둧��,�L#1C����繇z$u-��hJrQؐ+~�-��NU�Q�ۆ�}���a��� Cx�8�'w�-�����wd��J��[�ءh�D{T�z&<�j5�&܈�P8��g��TV��w��1Dmƴ=Y�ߺ��}�y��B��s�W�/=
��4b�y�����̒Lޫ oz�zwk�=e���I�s�E��8A��ǎ�D���P,?���0�mܟu��5��ڱ����VT���-pַ��H�o�te�s�{z۝)3��l��f�ld�4�]����g[�e���j�W��y��9���S�>�A� �B���4[�ç9�[��{���������o�9��;bگ�bU�3׻�~����{S�p�ȳk��{���j��?L�<�m_�S�Ӽ��]�����˂�O��Mj�9C[48tvm����#�����k2iˎ�j~Ϸ��K6�&wfa�X��'q��%;&���9��/C�<#S<��qtN]��Cf�Pt�Oڨq�X{U��Y�k���չ�9$F�wbW�q1=edUY�*�b�W}���Iw�F�v���Х��y\xG-�ex�N>W�D���h)\��ٖ�G�����{!8����'����C�+z��a�oǎM�&�w)}$����V3���F�T|�$"�k����W��Z�z��0l��ҢF�C���:y��>&�Ќ�r�m'sd֙�-D�EZ�{q��y"��2�g�B,5-!G
��'_V�[�]+c{	�"��;K%��ѭ9�C�M�����Um�q�=|�Yޘsc*�(����׃d��&͏�˽�tǛ�c0��!�+<u}L�{e�/w��Bx�-ӝQ�l\#����T����^�'���Cͫ�Z�שɈ��܉��n��m��eg@:��$��:!ow!u. 2�R�w;�d;;�T�{���ؿ{�s�����a���5X���]��x~_@�b�Ծ�MtH<�^��y{�w���~��K�cv�쀴S�h����G�yԥ�����ѣ~E��\k��v��u�}��Nu��L��v'vj���s{e���i��I�q��W�{t=�}����N����W��o��wT�w�v�Ů�J]E�[��
��{�{ׯmײE"ѫ����ǖ��='����\JP���|���wT��Vx˧u��YϷ�Z�o�W�OW�c�c�i��u]���V`Dx��䪕{�]i��\�c��}JT�����{"�gX���d#6�l-��:�P})SJmb�m�ݢz C4�u� �$m+�o���ɓ��<�����Uk��e����*�/��lj�k�^����E��`;��K���̻Yl��j+�#Ɯ�$_:ܷN�����,S�C���)8�0�ޢ;��ш�ѭ��-뛻����(�>�ƅQ�u��Pyu�j�m���j6RF�e��W�W���]�QyfE=Q,�td#9ޝPGo�-�6���d�����.\�������=ҔH��0w8�+��9�D��������=k3��IQ�cBU�J_�B!��Y�������.�f�$_��h�ty���.|ս�h�@W�8���,���Bѿb=��B��z��]�3��D�nn%���7��g��k���B[sm�G�'FM/��U�1}Վ_�z9�i���C�ב�N�]�'�n�@D�Nb[��""�,�"����O����ȿ�tv5��M��h�"�8�K��+�k���!��g_��"�Λ1�X�Yy�_0{nv.f$��mweC��+����qf.�n��ō�7�J:���KLl��y�ʾ{<���2�c+[8��A��l�G����ģsN./�7�e;��k���4�d���^�)xg*J�cM9�jC��^H1<�y����X֣^�7��M����u�[�V���u]Vي����`N&)d���e��$uz��;w��p�����J�Y��C�vF��y�n�M�|��}�����On��d.μ�$��t�t�Sݧ)�.]��(�����~1q�L���k�&}J'�{{������V�.�#�
x�C����zSx���'q�~SѲvsi(�Mz���=�s�T���A��	��4���8��?<� �y�j���qQzvV�Ǐ�'s#Wɂ�h�������1F>��<v��Jw�9�ٍ��7��t^I��V6=��񿁥��\̏b��[�82����q�۔}�e�n��_��)���?s}@;�"��'��=;�VmZ�mHU�#���C���L��y	9���(ccv��cq[qg)덨C�m�(u��v��鱅J�����-�[��/�'y���2�p3�
7�\����}l��/T�ɮ�"����:#��>G���*[�7��Sy!�orΚ;q<��M]\�OJ;����>��F����1g���������Msؔjvr�q��'r���"��%<'�h/��;=�؋��uv�g���s��ꚫWhs����VB��U:�t��*�l���ll[�~����SƧun��!�Uzk<�ߟ<.��x��|�uE^�|� ��Z��
����}]�ݘ����nq��#���w�vq���}_XO�o�cy�s�ר<��t'��ܛR�v�]�s�$r�z��ﮰ�utn/ms~Œ�3Y��zH��E�Ygm��q�uľf�{EH�B��:�t��;6����@lq�F�{ˎ���D�Vƴ&�Ey��>��f/vǳaK˜�Պ�}�CL�^�k�C�����@ι
c�ب�����q9�"=��&"}��nl�Nb붇m
�wcNN�&��Bt�f���[�Ӯ{g^:^6@�_����d�g�����2v�5[���ݤ��{WbW"Y�9�\~9��)4+G �8|Pg����g���F�f�|9XW�*�A�:��N;]�g�C�,�>�	v�Θu.K�����R���c��5lą��I���m�v�\[��A��N�kЭ��H�0��`u��ED�AU
;�]b��jČK�̜�1�'d/kk�<�\@��c�ͧ�$�r��u��4��A��1��.:ڷ��>qثͪ��ۥ���h
ˬ�T��|�>5iʝ�[��ˇ�ٮ�Gk�/p��8��^W�iz�,�{u�x�Ӕ���i�����Pv^l�s�am=:IT�DA3������-��=��'8��^=3}�U��:�����Y1�8��5svwAFT�W8L��
uz���u��1/m��\6�����ˋ��*uv��i+��z��^Ʀ��dR4"�_��k��on��^�롴S��Qg��U{4�h���-�l��	_W=��'sǛ�6�[�cs�����ذ
f�f���i�a+�v^����-!�/!���MOzk��\+H+%^1��
��2����ͬ�(���l��C�H� &l9�;�=W�h
����֒(3�9^f�헸�K��gw�ݽܭ��|��gK��	��n��NU�
b��k���T��j��=x�����`#hh	��ۭ�Yv�k#��G!��й�ݛ9�2]�,��:�N���e
�
����D�������7A�R˴�f��9� ج����W��י�� r�ٯm�r�L��h��cԔyK��N\�mf^k�0B��X�O�]̉4��J6�ܝ��oZ<p�J�.�yg�ۭ�$P#��8�5{�a�Tn`��<\x�:���=�i<��$���{�'��	q)��7<�7��!����{��AT��KmU���s)J�-��zi��5��b��$���;�l��
�l�훃Ni\-9;�/6�9e�s�+�Z8��c��;5�Xu�������Ǯ^���̆Q��\Y(�2Dl;��\V̻�u�NBo0�7qf^�^m �M�nW��-�޷��׃{�>��\��κ�� ���i(���kZ�h(��.	�55:�>lK���k��h�oV��j�����mRMy���h�jMh�lF��X��\�G���
�Ѫ�j& ��\j6B�47��d(��Sݦ���E=Z�m=l�MkUL3բ���MD��DUEDP$� �2��0�#��Nzuo;!��{�c]�=�ѱ�5���� �%�Dl�s�y\���Vu�̻dp��y��?�N�沤^��g�Ο���ꧫ�~j(�@���*�lD��^5�*����o�ƶ�G�~f��u������w��5�N��\6J5/5��3�SX��8N�9Qcj�����(��UD �(D�*���jó*�mH.�[��ȳ�@�9JY����U��Q����++��oDB��Et��X�⾯pCy����fK�{��C������R!*��])J�z���K�7����<��I~�ć����v97�Dʩ�Lv���"�\Ome��V�ǯ�*�.����:�}Tk�w���Ʊ�G+=�fJ^,]D��I�֒�%�F���kξ�y盝��],�_PŞP�L12���n����x{����Lc;}u������z~�>bNҒbz[�N��j�{r�WW�G�/��i�t�ifY=EJ�Н�a��?E�I�J����w����&�;u^�Ό�S�:� 6e�� �s묢U:�seb S]y/9rN1B��E�*^��n�.���k!�٭��ק���ߦTr@�ߠ�W-���0�A�uX�ֲ4T�s�Oz@BUgd�6~��^JvT�/�;i���Q���	��wYg�V�KO�f�ڿ"z��7{G��rU�9;�P�*�L�ҫg�K�Yi���.�`_y����
�ܚ�<�on�:����q����H߫��n|{Σ9�.&��8��n�]ײ�.�<ڻY�=P�+i��5��}��ۣY���\w��(�izjGw.�ݿL���1.���!0cp}�x����T�E�E�p�r~�w��+ �*OqdyP7��4�}�����N���0%<��F�Y�_i�7�bZ?	��R����O/��3��l~�N��wԣ8d3�� =o�	�Bt���+����17}{��3�w_?��g�{6n�n�j��|Y������Ƌٗ=�����y���us]�ݒ"��y��'�z	�˧����!,:�̆|�s��,;8��C�Xn�`�p��v��}wYO;Yo�5�Yjt��3�۳hE�*SSRT�4���Mչ��׫��gW;����/�����5��$�~��+���k;��OЌɐ��TZ&�-Tg���zG:1�0ͯ��&<��̽��95����p��9�Z����.����{6��7��W�
��-�w�����LJ���a2��x�yTX^�/U�WZ͚0J�W���|v�n��/_�O�S5�v}]gh����R�j��؆kss9��n��.ͬ�S}>��{v�?]�t'x�r�܅�5UM��ފko���7��s��n_F^��_��U���k�:�*��{6�9\j/�T���{��$��m����W;�䬯�ʃ,{]9��в���P���;���_E!��^�}�.�D�J�2�Y���@U�E�<��x��GC��_]���iX;���{0ٙ`92�)��;��K���%)��-�<<��&S���v����2Qu�ڬ�d6g�ާV���$�4A�
�w������;B2���a'ۏV�pMO
ٶ�n��l�<��~�۞ޢ�9>�{����/�����~1��G���js^��y�f���v�Z��A@��G��N�[@��B��.M�o����W�i��,jݕ>�l�ج��"1J?%�m�K�|�r���.['gd�?\Yך~�h7Y!�ߛ�ϧ��ռ���J�NE��E��D"s��[5���a&�D^��w��{��ھ�A���S���v/�7|Ϯ�o���S��kA��8�4��{1��Փ#$ե{��.���P裧}^b�o���2�f,��o{�>ӓ��v���9徉ͪ��z���*lNM�`���|T�O=ɳ���p�(���'���������)Or��[Z�y����\2��~����)����31�������]��eV�,����{̾��٭��K4q��Q�2�d;��T�m3D*�U�Wu)K��*]�-�Ε�j��}W���e�fM�	�¸�&j��7YŃGj���)[�w��b���n�(�Uz�;�^Ѫw97)����ݽG��r'��o\�s��$5�=�yweHqYC{�W��=��.����ό|^��^��d���B�O�_!���x����93�����&Wߍ�����y�W�=ն�z:���MՏ��&Pq�2*��w)e�ZԲ�=���;�ӻ���1�5v��Q��}A��C�����эj�zwy��骞ߢ�Cci���j�e��q0�  ]�Q�r��;�7�d
�n�ywΫ]j1=)��*������)�[P����5��a|��s�ΡyG��r\���\eP��}G=y]N(��S������=��(�ubh��������:���c�^��=��@t�^���S�{�"���*��d:�BU����2��pg��\y��]��5���5�o�M�Y����"I,�Y���w�r^�F9v�i򛽻���8>�J�`7�Cn�Rh�{�5���r*w5�U�M���<�����ެ��'{�Q���C��c�(���3x�ڷ��Myky����/o|�s��#�oc��ɵ����;<Ș���{�p��VU�g���f���]3��k�p�ۑj��w2�N*���;;�z�:q�h��gm��j���2��O��q�r`�m���-��|~Z�)1�=��d��\��]z�{)G���zl_u����!^e&���跗e�5Jۧ�e��k�mG�'��۝��E@}�\��+�jym�X����
'W��m8=��X]%��S�K�Z��{�wɟ�e��r�Hg�L��Y�?8�X<��zf�|pE���A�l�
�X��Wi�0��{�L,�I[�U��yW�7�Wu�gWOP��f�՜�ƻb�coj�D#�LDo�z��ܬ�C�n�YiSF���@U
.s�1�s�F�]%7'`�����������(�����(�?v��c�9O9q]�[b��[[a�C���u����*lW]W�#�
�#z�Y�%���v�Ђ���ԕ/ߏ���؍������g!8�T,��,�ڳ��{�9�j�q��4=G��Q�M��9��BURy)R摫]��E���T�]+�W_ī���}P�c��Z�6�,Y����G���T��qo<ţ�U���G�#����\�������Z�B�Y��|_�8|����a>�J��=���ܛ��B�=ԡ�U�	Д؞��yQ�����{�ף�L�'��8-�{%�ɾ��v
`Rk��N�B���n4�˝�3�Y�Q���m���m�ڗ�z�����o��W�=��{3Įh�3Y��*7��k*���^��.N�]��<;`+T�WX�S�N�@ci{��߫ǧ�Z��̺r��N��T�{DY�D�9�4���3�r�2�5�ޭ����\l�MX��n>�Wx��& 0����1K{<r�WO2z��\@�dN+�RQxWFD���`��鈩\�V��;���ʺx��k9v��V�^��}�Y��̘t5��k���b}�3��P���_�3���p՗_��ҫ��uP��a�[u�j���G��5=�����L����^F
\�zd;͇?��S���Q~�����Id�wQ�x�nɪ��s�hn^�%�� )��攚@�~�;�I�/<�|x�!�pn��0�j8Y�����
����:W�#���0���1�K�މ���f����\{Ti(8��Jbga�\�<H��`=�c�Fd�':\^>�׻>[��ד�$Enj�"�N��uS\Kbf�-vH���U���v�Y��7<�z/�Q�8��rD�.A���H�dk�QlK@��u'�|�U�\��sL���n��G$��Usxc#��f�ʞ�C��%M�Ǒ��o*�]<�_�ԍRD�6����E��ɱ|9�Q��N/!~��+��6cc�V���͞f:=Qq�>RXv"f���[#*�l��	R.<�M�#�nG��(���?�+	�s-�i�a-��_=�X7�.��y3	�;/vzm�ݯ�a�՜=��B�l�5�hT����:*��5&��T}�el+J��ѭ��h��1��U�s?���[>aQ0quA]t&����d�|UL��Ux�Ek1c=h:�˴�lmOis��2�������	��k�2���R��{*��_�Epy���Y��2{�F��a�ZY�"��#<�x���J����\��[%��/���+��ٵw��G��'������Z5`H�Y�"�s�L$;uVM�Mp���*��p����Oz�S7�J2էu��e��\N�ڌ��D] R�}������c/��T�c����������ᘞ���G���.LC�o��"��/"���Hu���zu��f1ld��l�S�{��������Ftv�jtH��b�F�&[����p��K��ڬ��[
c��:V ���n�)��y�!��0sB9Q���7�sfߡ��s�}��K�.���E���N2b�`H�����w3]�jfo\��[q1��a�ո��gK�Z�`u~\d�k�l��>Q���pWF��Y��ꙇ�f��f�	�\�Fٹdឭa��R��y$^�=�5���}\ˍ�"�7��vwk;�Jϵé���.�z�C�S2s�K1=��N��	�����t&�vg%Z��a�P�����IZ��f���35+
�#�7ʷ����Uy',�=�r����l?&��{�JQ�TQ��mL0���9OD�<ɏk��I�pȋ��nv>��*gx		Ҟ���v궮2�� ת����Bj�1���s���G{w5�ܖl?�l���f�(ɯ���c��{�I�o�R��a�雱�
8��:�����q���B�ga����Z���6�ϫ��V�SP�T]������ك���o��?��3zA�@�/O�=�89�P;�rK�g:���Ѯ{<�ޠ�c�R��3}f�C�:���v�y�L�r.Ej����Gl���1�>tC��z.�d�����
��a���d:k��R��>9���c�˩I�����[���t+�j�l8��C�s�lI�sL�coꅥ�\s�B�N���OX��)�mON(��r]M�s�#X��Ӓ��9��s���3k"&"���[+IO�H>�k�MB=�w]�D�z^���"�y������O�-�zN���D�����";{"���I������'�$@���&��B��x�	Ad��::�3j9���Ό?�����>G�:]l�4r�����tXJ;�gn�n�H
��m��ٓ��l�nj<=h�r���O��l������2�+����s�x�����K�W@��>#^���\8;�i�Cq\̍���D1v�h��I�����Q��a���(���WKG�k�iV���?�UO7����U���c�R5H�=̷���)𢋝n��]u�t�I��[��1b�I��¸GR0��f;D�(J3|��L�>}ޕ�mGO�?W��/f�X���<4f��)�)�ʶ��:i�k{Mm.�]��`h;'��B����xCFw��󄴂3����w��,�KstԤ�]�ő��h��3�����|���n�>�2֗b75��b��%'7�a�������|X��<�;;�֌��n.4�� �5����ݼ�gk�x�mi�3|����:���%<�z����`f-6�ý���$���u�|�*YM���4��CM?M�c�l׈퓰{U����3���S�GFlڏc���w�,�gU���ڧ�Vm<�Un\�;�)�y\���2k�U�%L�)J���ΗNt�..bK�7cV9�Zty�o��hW�J ��&�Oa�N�#��Yǀ��\畠���}�����Ş�^OE��V<h�	1�a	���C�`�q��,��6>Ri����g�nb�Zu�ү��^�G�8�ݯu�4��y���^s��� )$���e���|�_h�wWfߛ̏.Hc��v��Q�.��	j�{w٨d>����f��:�Pgp�g�M>�-t�c~�5J4����v+Q������������Cˎ���n�j��r���78��W�=5Ԫ4g8�^aR�bt�q�|E"�-�CObNA����+n�02�h	���C_���u;���U���	��>k(�ضv&I:��wK�|��j�]"���Q��/b��Um݅�>��V�؍M2"�-��5ʨ0���/��7ܗX;�cn2�)��֏����]��L �{΁:n��d	�M�;u_��®��:QsV���:��*��Sb���nE�����佶&�ʳ�@ܬ{�.���F�>�_0����ޏ/�Aմ�0W�9!�n�ȷ���E:pG�V���sfZO�֬�ʂ��ģT`D<�3h��_M=��G!`��"�O
8�jj��W��� �+����Ծ刍R�]��d��:�XYX�;�(̤ ��/�^K׋on�m��6�-��vn�!��X�#��r����k���tQ#�[x��^9���`����ʈ�*�
fB&H���)��*�Z�)��3E1rն(&h"JJ��cL�ͪ����lĕTE	�a��*)���DHD�PS��lj�J����&!�����JӪ<A���������D�HL�IDh{�E��LSUDEAA1ATQDT5UQB�T��l�!���8��i��k��CThqT�؈��lU!U�к�T45UQ5Bw�F�Q��}\v��cb�f@�6t$g1[�9/��%���#*7���cU�����mu�`.L��7�h����f8���0�0�y�+}� $.��2ߚ_�A��ލt��<5jJ��s��TP�Dq�}wbN�-�=�kȋ�Vd*�W{�J'�}(.7t�"�~����?�v����/�DTR�v8�X�;/A���Q�p���]��^�D���~-�����`@��F]��`eȎ�L)1����R�B�5���ܾ�w�!Y'_����zQ3����:�S�fKU�{i&c#��4|����^��^���*)�%J���2�YX���LB�L��!���j��NO����Y�V{"�e����Y/����U
��:c"�:�ӟdK0�����S�3���?�2��Mk�����j'�����]�H5Q�;�<��B,2�J�N�b�lɏ/M�eaLVNd��A1��v�UkS��$\q�N='m?$(w��t)l�9�萌i�/��|7v�,>������L�4��*�W��u��g�y����+����O;�5��Kd�Z�������z���r�6���q\��,�7�]z[6B����y�7})�3�cn
��`;=}bsfKi������N��I���3����MoB�ι�(��h�j>�^����=yr矪m�g����(��ɾ���T_󔐆b����N~b�|�M�J�)�-/������t��ϝ��l����FDAF�z賳���GLu �"�[t�@ܼ��\�K����Z�z�|�c"������d�2��w\�I�;�|{�>��}gbϩ/H��RXt����$��}m��~��k6=׃i�_ʇ�{���f�ʋqg�Lգ��1�n�������r_*���fkMno�axS��A��,��I���c���
iʦ4�yY~J��g6܉1�=�*���z�9�{���׷�ù��yTN�+~Lܦ�'n���7oޯ�{f�7o{ң(\�j���E�La	�^�,)^�S��G/�D���ae�ՇN/=Jk�w�����Z��-�%�S=l�v�:&R�cz� qY���^2�6�/�7$_����*��xXێP=�̉q.3+�dGAߣ]��f]{�H�]{+��:q�C���!l�9���qİ4��݅�<��z̔��S�Ä��יF^u55T�	~]�GԹJFm��ו�7��Eg`�(���D����ھ�[Ӧ��� ��E�^���@F��1�]K粢g-T`�y�
�o�����4L¼Us�/*=Q<rA���&:S|Hb�`=��!P���V컫��~fzs�pԑ�������c�6'-�H���.$�~c���cL�s��׷���X����"��d��8lr����r6is�<M�W���T)r�N�9�#���8����\=)���+�B롃'
9*��7��w{=�+�T"���:w��0�ϡ��|*o�}�ž�/brW.u����A�'���J<��K���KY���[��l�crB�4�U��Y7�t��Ҳ4����_e�N��c�{/�n�3/l<���-_�N"=����=<��C��nzZ��Ge��||੡z��Բl��f���f$�&�VH�X�/ў��Ӿ���nG1�Ǥ��|cr*��=?:]g&���j����m�n��\M�d"�[�zh�2��X�E��c��&�q<��v~3�m���$Z�ύ���cJݮӊ���(v��S���)���o����A��H�1U�W�ԙO�֔�0�ڍ蟅�������)���>�N��{�u�@�1����U��S�)_������^��ؔ��}��}>"[�T��U;Q���ހ�Rpwv7z�,�E�9��
����ccz���Ș�`�SC4��Z��
�T��?{��츸���^Y��㎌�x�x�TI��b�'�N?zG��\a$��s!��xnew��eA�a�l�q霮~7F_yf�912�!̿j��+<������p?��k��C���6*���6�F�	1�`��M�b!v�<kA�S�x���;b㹓���/�s;�P��n�~0��؞��".n���cNK�~uGE��1P�r�Y��'���<Y�
7X��7�����y[˱9 t1�'�[p�As3\�b�R57�����=��W���YV�rYU�w{u{Fxd�0>�Y.dw���v�MDoR``��������.�IA�;�Pе���z%�N�?���&����&��z�q'���9I�5x����!
`�������O��,�a�c���{���!Ξ[����ޮ范�Gz���^MET_C9��}oo{4�S#����p����˸�_�&�eM�Ev�fd��GWb��,���qޓ�{_���nz��}�ih���.M�v���1]ټ�Nv���O�#���,1�UQO��Mir�1x��.}����������y��Â���fw�<L��rDgE�Tv'��&"��#hƗ����_36�\/z����nl��.�Ǝ��l����W��^k��c���[*�s,@7٫�W�)d�+ޔ֧�,��9�$�SM���~O�FA9��v�{��-�S��~��ڔ�G'� �3�
q�����ppu��ת72:�a��`�������F�r6����]�K7!-�}�M.�����+4_���C��c��n�d�@���.�z�tgD+e��}z��p�V:U3���t\� "�?h���Yl���:�S�иy5e�MoE>މ���w�2`l��qt�z�fJ�o���t���^��D��n��gT��IĢg5��|��u��^PP����r1�TE��^���}N-֑��"w���-kw_D�:X5Q~+bĿ^ъۆ���H'&���^A�����5O/Vq����ڞI���[R�6a��|��\p'ywn��x(頰3,@疟)��V���ҷ��",g��ؽqyE��/Ō�¯���DN��v�J����J�UU}�򒎽��ޑ�L[&���\L=�C1Z๤K�r�E}�~6�����T�����޾�O#�ukfvΟD�ٟ�VO�c�~�v9	�%L�P�B�3SO����cѰ��q���#�@yP�6�MX4.<����ˡ��s-K��l���z�	��T���Ⱥ(dNF�>�1Z鎫H�ը��c��٬��k���c4���D�5�ݍH��q�s�K���'/]Fy�Fg2��0�f�(���s��/��|��ٱ��sP�hf157	���3����l�XlZ���D�\T����(����M�VT�tO{e�^r��y�S���͇��1��1>p^�(y~��&�g�^�����ѥ਱�鿜xfF�]lA�@��^,�vd4��^(>ж"��Q��NZ�&����<��"���F[�ELNGW��WO�Ov��xܧ���P7x{�ar�I`7䑓Am19�X)����1�P�߾���c�5��^���kf�_�ܥq�v��R�Ve�b�WJ.ѷ������ Α]���E�_�
ՠ��-}<ڕ��4WJ��W&�n�s������y�,^��a=c8�t�ot��v����Bs=���D���&0��ޑ�.�t�9���Sl�F\X��p2|7��VTE�G�9o���3��d�F��Z�C �-��L�ш�����ԣS�9~�7��
�D!�K��>��ݣ�j5C�D�
{��η�$G��2�v�M#��.�+6k�ҌD/9R"�7��ȇ��~����\��3!s�D]�>�.uK�|`���l������{�M������0��=���q�ø��e�`�b#���%L�d��.�9���A�t@|��I�����UyQB��u܃��
K�JR$�>���q#.٬��h��󨽤���#��+�iq����S��'�(Ti'�aݘ��Y�O��tmu�8���j�C� �F�胤f�3��}Q}~�[�P6��.A�9��J<�w3VZ~U3H[�x�5�����`r�Ѩ���3k����/�{ph��fX�w�Wrs�s�"����2u�4��=�h��~��NԖe�˰/��B���5oQ��W��L3�ɡ[Q��]z�P�P�s��8w��.�C[��2o.�n1�qHL
�����Z�AW23�6y�x�h\k�i۞~;��}]N���@���n����7��\�}B�Z����D���H��YyV��G�6���}<�ﮖ>�Ҿ�Ϧ���`QU�5v�TZ;��	S�MJC�T���|�R|�<΍�1��g�v�������Tg����i;q�P(\آ&�S蚍;迶�wG��Zdش�kw:g�eE��[9�	<l෮z+샚���Mq=`��`���r;��Y�4{1q�F��x�Ūɦ�Wצ.YF��Ed��/������W�-Od75�<�߁�"��o�9�8c���<���Tv])���,�6h;�}P����ݽM󊨤�2dDYl�(�Eg��5tFD���6Ǣ^�'ٷ|;kݫ�I�1}�9i���	�^3 �-�F#L�-���ﲶ��y�÷���&'���ڈ�tF�t5�������2X�P��y�=ί�q��=�6=�g���b�2�|9А����I����1����ٛDtKB^��:�{*%�Z���091D�4�ֺ�v�\�}��&��X"qll��')���e���PT#��]ԗ������8)��1=a�- &8:� �J>نo/
����Z�|��n���*k����B1I*~���?q����d1���W�G%��8��}4&����L�9��u�⢷j�z�y�J[��J�'��md;�vfk�Tc*EBus��!l��2/�.9��m��};e�;�w{�	\]D��_��q;�'C�bw�ar!u�Qz�o��Ε�D3.�G9#��;3��h��w���8���q�%o/c��s4t�Ww2N{4E��A�^���[��Eꪈ�>�o
�nR�D�x���!:=gcK��s^j��|.j[g�"7&3�+���^�,eE��^�¼���:Ƭ�jQ�>)�B	?��l��n��	�?<������;,M+��BZiYɛ���X�&�ӝӪ�}�JجbNz�Sф�t���Q;�{��#� X'_MßEV�#}�7��b��ܦK�:c�Vbi�c��q��p������㯲���{�4w{J�þ�%N�T} x�.�bw��P/o>���%���)}T~������l���`��)��6��ǟ�:>ײKb����<��V���N�6p��T򕸐ʅ����O��++�����.�p�!��5���8��4��ې$2WT����i�S��t>�Ǳ݋����cG�i����X���b7"N���D(�pH���1�B��w��zY��r�5rC@���\#��J�g��,�ى}Ly3%�Uk��e�b���\��y��҉����|��W��������*.�{Ǔ������
�*�&Jީ��Ĺ^�
�r�dz��c���\b��6�J�T�xRY�|Ѩ�D�~}�� 3{�"\��f�~%�7�Z�Y���ě�gOrى.�8$���lJ�E�~Zad���<�X>�o�_�4"����L����2�P+�ˋ�-�m�Z��R��7��q>��C��)�sx׳�ICS��z�~$EhE���=~�?��`��Z_hR]�G#b(٣���*���3��=P�֔&U�:�%�}��ק<*=���c��S��c�	�|��y2f��t��}t��k^�t��'���9p�F����থd#�~�3*��x�[�>�x��A�}�'�ol�����iU�����.����ջ� Fq�Y�ϼ�^��LΊhR+&��PeV�Z�-F�6wID;��m��&F�Κ�v�1>�Y�6�P����Ε�R�o�4ק����q�=��<U�ԍԫ��;7j)��{U��!�1�8Y�9s�,Jf��<�����BD��-b`e���#n���UA�Gj}��#i��i�����x��{k2��V�f3���l�I=�-��v_L��Lo*�2�f��ݴ޶'v��/�;���v�G�������t�5�Ku�;�}���}�L�w�����F\�NZԏR�.L�hf�� ���V�q�_�q��î%JϦT�&.�@���:�z�9D5i;Ä=I�Nks0�[G�4����FW-���^f�q�i�tN���F��p,��M��sx�������c~y��N�!r
��R-���2���F�^��mN��pfک��ގ���V�wՆ̌9y�N�
��ۅ�"t쓵А�i\3��.Z�<j�-��� K�(@���w�H�NOb�0p�*����YЫ�#Ǖ�7^� 9����,��E�g_A�^w��/N��İe�&*S��;��N�
� dY[�W�I�wS]FF;�d�.�����N�w6���נ���k�8�ІP}t��FP�O�3�jw���wt�Ȟ]P��2=h>���^9^L��ћ�u{�͎h�`Ij�~5��V�ɺ�my.�}P�- ۣϛ�|��M|��^���$�G����� +4�Ҳ�L�)�E6��	�����Z���u^-Z��)oi9���X��n\��(Ew&{�̆�}�PD��=3gDe��W<;����e����E��缷R�X1Nxr��qs7�|���K����1�k��_I1.��T�>�[�.���m��ڳȞ���G+�F�yN�q��K	õ��o��]����떳*�����jn�+�={�p��UDy�,��}-C;<�^�<��I��tC�+�fk2�w�v�"!|c\�\oh�iGR�nk�=퓊e���<#�y�#څD�}`���X� �I �H�v�$��Ai�S�j�I���!Y5M
H%elU�B���0�웮�l�p�pq���f�{jFY��ĕ%��Q�RHf2܊�ˋ<��y�
�O���β��c�HUP�Uu:�bb

H����j�+Z���

��JB���3͠ccAM�EE��RQMP���Phj �� �MD�!9:v5!�G3�m&��1i�'�p��嗓�Ns�0mY"j��i���ѭ%CZ]m��QA�s	�u���um��ES��E͎p�Wl4�1`�ABi��PkVɭ+�(�h5U�O1����4DQ�O�yCA�˖!�l ��R��(���A5%G6H�F�hփ�U��-�@D�M�c`�Di
Bch#4Rm��Z�N���LA��k�W0i9i�AkPb1&�4i�b4�V�>:��k�{�Ǐ^��s ��kiAt��FP�q
ų�������}�|����\ŨӒ�������oU��Q���=���b�٩Ĳ�ݥ@��l*���{[�ޣ�Ĭ�u����M�۽���2,>
o	n"$Zg԰鮆kb�0�u�Gv�Y
k=�F�z��^q)�D�[�-l�4)����hHu���9��Foxx�a���~�s>sWn;���&~R��z�F�[l0'��Cq�q�d_�bЕ��v��^���r���/�1��#��p�å
.3qP~)�����;���^��k]�Y�|��P~f:��Bb�z��8��-	{���ף@���V��@ѓ��r/|v�ɼ�~p���ƈ��ˈ�G�obDF�A�N?��̲�uؕ»������6��G��Ú{������iEߩ����cn9@���(������!u�l��9����]�?Blz�kŌ#B�a禀��򙞸�̰���Jx���Z�0�k��G�L�m�	��/��&_U�*�a^�
�lKW��&$���UF������zg��zv���ܕ���M�P=؅DT\��P�qV!�ֺ�
�pw���4I��V:e��7��<dk#חW������4�,�ު��ugga޷��-\���ǎ�{`N�@��q�B]<���~�u�>���M���~���Ele;�w>d��,8њ&�R�&�7/��y��N��Qs��j)�F�v�~î���\{��}=�#_�MF��_�l��V`.1k��ɑ\��tp�+�WB���
��n���C��b��P�/.<��#��77�������:Y.<Y��� �̬��ߧ��
o�B�>��eV�,����c�ܖ��s��q>�^>��*���ػj�"V�%�Y1Ƣ3c).;��6�)�*ro-��uj2���6�����o<��x�}_E��ٌ��fK-QS+r\z&����B�+�;[
+�=,��]r���Ъ3��:o�X��.;�w���"����Wq>�n;�7wn%���l�љ��>�w���=&r7m_\@��&�F�)�+��=�yFi����X��w���e+(9C\�k��B�r��SH�C���)Ƞ"D�*�2�����+��&.�_�d	7&�r�X�-S�.�����̹w6����M���l�ܺ�]=���:�8}�8�=KU[��JƼ��ܽ�;4G{�dO�ފ��餺Y �]�������rΣ��[=���6NLK��I�<?�#��e|ؤ��1�(\O1P� Od߂,����v}6u#C=���c�L1���)�T}��!v!??�}rd.���B��ȶ��շaw'��pFL�BW&+��n2=��k$r~pt�D�,��J�Xp��N̺��=�������{�4
>����g#f ��Y��#��V�^V� �5
�� 0��+%�B�1G�Uçfzo�}N}�獦nMq�U�[��Y��,��t��������R|�I�� ���H��z`g�r+V��g�x��b��J��Pм���L�UzX�Q7�1N�
]���"'-�m����z%��d�&Ǚ"j�:�ƅ����&�8ǯw��P���Y�I�4&c����%|�u��0�צ.:���u�Du�&����)+��+�9�l�Q�c��k6�KWT������>��O{�������#���gc�zE�t���/N�Bj�/�Y����\�0AX9���*Ru�.��Q����3�Q�o�y�0��m���)t�~���\N�b���V�植ud����_>nmң�ne�QU۬�bq��+����EO'E�?�ݶ�1�9�����x�<����la���j�{%���<B�\ �p5�{���g�=C��{���ܕ�'��A�lD��*��{�D�U��`w��_{�I�5�g�Ȧ'��1�*cM�c��Q��/��:��<ę�	_��>������d�5�m�٨TrҲ��bU��S�cf�7�d�x�on:��F�ܺ�=��|�dp�fY���f�sL��<�b@���-�>�����Ԧ��7O��*��n�p'Q;�Rѱ�'�I���n<$�C�/��eҚ�~��E��Ѯ�F`q��`,PeOL����bӰ ��u�7.}��f�b1�VO��ߪ3�FcB�F��e�_���B��%����ZY��"�{�f-P2�Omn+Y��{{��r���T�QG��̱�n�,Ér�rԳ2��٘Vtx�(ӕW� /��N�Y/�Fso�6Ԝ�J��<} �W�U;�<%��`�k�0�+w:z&��b���Y���(�� |�{��uR���p��[[�)�n��q��3���&�7�i��r���F�F�Xl�;Y�2�9Gg�w;��g�5�֟�յ��2Vo�o���Nj���v;����f-�����m�Ǹ����6��c��9Nbo��+��%�~��<�]�:&�|J�'�|�"�,��^=��|�C�����-d�|���M{o���o+6�/5[33ͪ�=��\ �:�ps�(���e85?_<7���&�c���D���������gg�*_�s���Pz�Ш@���V�4q҃݊���Oٵ[G����x����>q�n\,6�!� �-�FB�{��XȻ�ƜoC�B���O�-�ȼ�UJ�~JL�;a�ec���.6c&;Lq��B�k���[{*o�I���α~�YV�v;ڥ[��w~� ��ö�{�����X�1��F½���p�5T�j����1�d�1*��P�V�
��]����h��dΎ`��U�mʽ����i��b�j�#ʏ`�2FK�+���t��D��H�~l���AӋ��u~ɍɪ��]G{�_CHk
�Ǔ�OV�7�/���q̆���CF�r
����.ϥ�f<��,��Bi���AҊ=FM�{:\T�� �V�u��^�YؼN{߽@�8���F;<�^G?O4����]e� k�ք���/e(�I���<.�fMk^�S�*&s�����}~��}�zx�GX�����+obDF��{��l2�����nw�����_iS+C���ܣ2P��˜�'��U�阰��,�A:S�� E�
����x��ә���D*��H&酴\�:�����@B��������k8w��s^"D�9�q3�@��8Q��aݑ��.�F�>0�wg����a�[: �lt �2���TQ��hK�j�2�a��Gx̡yUcp�'	�'Z޴� �Y�*fLC�s]7����ca�dS�s_/p�P3Fp��GEF��U5���ۻ��#��F˙�v48�bf��m���Y��I�_��ܸ���6��>���᝶���|��a[&XȒ��7���Ǽ�OqL	��z+��;ǫ!�Q���f�k�����Ǽ�rlTc���:<��~��7=��k�$��Ss��ν]{p��vE�ao�@֫b'�ΉO�yQ��3bb8�؄*^h��p�k�,;q��I��2n�d�f��<�}W�gv!����|.]�^/��n..����S���Q�7�2��.M�`;�ݯ��qD�SXT�U@b4�ɴ�/����<m�Ԙ�}���fS�ރvd�-��w��?�������.7�#�ڰ��a��`1kzG�9ЦmQOI�[K#�E}	���1��Y���=;��r��ٕ�2��������͞�yV�yH�2�O6�u��0:�A��+=�D,��+������C^s��6�9��O����ۃ�mv$�0���v�G����'�S�s;4j�q���V`9CX^��q&7���[�R���*��5ݥ��6O,5l->Ԅ��z)%�d���_�(���f,3��Bq��1~��oc۱�>��:���MB�%��Dƕ�ؑ"��gG��
n�P�P�fp�����*�0�>'�A+۷������bluW�Y#�:x,���]��:Z+^�9cɩq�'&���A1�N�y��bg��bm+�* ����"\N�~<G�Z�@��5����ba�~ �eF��ˑ�TXs9:���&3�Q�MS�!�&.j'��>��]������۲r4� ���Lm;���xҙ����O+~�jq3S��A�~��t����,���D���lG�]��ӑ�z��+�3����]bcɵ�8:M�o@��>2�׶�E���f���N����i�ɺ�̰E��}5jp�@�^h��cت˺&�b���\�q�  �dv�N��/Dba�#�����rk�Cή4)���&]��Snp"mU�%�y�z�cUɹ�jd!�Ao���]��&��z�Tzz���u�������N�r'���2rn>�Wf��XNNt�p�,JU��Nk\ �Å��:�5��y7:Ẃ��Ԝ���>���3�Q<9p�v<����N�J ����y�޺����<��T�YG����s]�%x9�}����(��n�.ey���7/,�w2�e��Y��P�3mu�K�ފ2+�\4������ȑc`ND�o-G���$ ǝI��bPz��j7c�h��X���D9ά������%�d�~�����T��0p�V�ۯ�K;�s$V�/�8�I��=7>�4�?d�������i�S�-`�Oy�;���Ι].I=�Ř�ˣr<'Y���a˛���}e�//�9�saz��7#��� Ϲ�r7v�Њ7 �>}����fr{�.�Iii̚
�m:ػ�X����Gx.�#_ؑq]~��Y�9��:�-|��?�ryo�gr�/�ȃ�.�5ᠦޱ2�w�-i��evp��r"��=ϓ�%������D�Ұ�U��Km�}ó�R�~uȡwz<om>��Vu]����>�D�V��F�C>8�3�x\VuZ�ٮ'��h���E�0��6��l���fe�6��#�s��u�<�L�Ũ�~Т���ϹY��������=�>��P�*�F)8.k�r��h�G,e�{z�Υ�P�s>u(_�~��G�%Q���	�Lw��<kQ���1]n{>��q�'�GFZ���פ�- ǎ�r���=U�qA�}Kxڵ��Kz�]o���1�q 8�"V�:�)5�̸�X�v�H�l�96{:oouW{�,`��3��]3>��d����><Q�{F�h�dM�{k���S38.�lim�����`�(�;d�ˏ*�;ǘ(E�Q0.Dr9;�D��+�L��/�wP'�э��'_K'�~Ci-�Y!��usO�)qqp�&'#��ϰ��CsA2�;ݚ��xO����7D��+GJ�����zTב�ʹ3-Z˲��ǹ ���G��ݡi�'��@�h�~y���������=��Q��귔�3�����ae��kv,oa�NV�ԙ]t�>��s��uaژѪ��22��/��	�}ں�C�&�ަ�\�)�n=�VE�m�>���a7�{蛹��L�*�g�eؙ�G������V>G��3y���w�{��o����z2<��8�5�J���f� �T�}��.�2t��3Xy�9u�3���Ӟ
|.�|)���4}/��,������H�y"����_�8�c�z�oR�~�ѝS��$�����CHk�z�>�1����0QS@j�a��=;1���w�ݽ2�c=�*kI�,������oD���7Nj��{<������goq�f��=7���2�&>\���~5_k��)d��u!���7��kǦ�����-.��]�����I\. �Y��k�
�9�wT����QXj�j���"K��i��pA��%�L�rzd=��6"{]�	�٪�+T��@���t��]�����>2��.o�Au��g�z�?5�:|T>�߼�s�]������uZ �S3�J����#��z�y���ve�Pe�2p��m����&S��DD�DI"`�	��!0�D5� �C����p�� {����
�º�@�Y��VX4��!���\���e�&�C�h��ѓ�n�}�Eӛf����4ď�]�
n%�sC
�D�^"��<އu��3Y9�-k��5y^���n�e�g��ng�S}�-N8kU�)�I��np#�g7}�.���5!�þ6��걟4�`� �4�!صn��8��ɉ|""�-��n���u{�-)�eZ�G�:�fhUv��dGrk��.�f��Am���7���j �X�,r�s���nFO����᫶lW�S�}�uS��e�>��w�m�i9!��Q��;�G}��G86��Ue�VA�s�R�ҷ�_E1�n��
j0�X>4u��93A,�-�ݣ��t�YF���t�*���c�3t�o,�4ro�t�֗�3���Q�Y�P�V��"�r�8��Z�w�d)�u±�6��퓕ܰ�ZL��F��@ytX��Λ���;#�U��������Cݚ��]J����S�e�UdgJ��Q��{���{��zq����N83�.:(�V�<�i��R�S���K�|��v�❛����b�ό�y���xnCG����\�y�h�l�����H�V��1���^޸c���x��h]�fW쾴�M͍��O�\(b2!�f�PD6���Ʊ<H���W4xsr7�y�l޺[B�(��lS�ڴ��՗776��u�U#�Y��}��Ʃs�0.w7T_#�Ba<�7�/��Ks�T�� �n�U}�c<I�����Ļ_�}O�J,ênC�2v_!�6����y������w�M�l۽Gr��H��p��/7绹X�T�]�ʲzf��X�}ŷ�K��  %�*7��2��o+M2�n�QR=�2Hw���]� βY�p�ٲ2b.�Cr��hX+2��M0���L�卌�^�̵�B��s���+��]���.��F��[�t)]�eE|�t��^�kkVmV����Ym�'�n	K0bڇ�dK��p�7D��B��s�۴NdE�rE#z��{��7�^�挴h���G>���:k���(��U�=��|�$�q>���4r���q�����:�cZ*"�vNq��� �inֽ���drZ��J�ar	��be�-Ba\FwV�y99	���ȏ^�s�" ��s�j8��8��
��x���%sgZt%�+A�q�NI�ڳ�)�֊��9�Xh(j����&&���	*�V��*�X�l������h
�+lRQ�Е���O#s�ZJ9f�����1�gDELZ�P��Th�5Z�h4�O6(�H�mوCG$�E4r1�JM�EMld(��d+O�C�&��GU)ː:*4�J
��ւ���y��Kɡ�9&�"]bJQ����0��� �%4rM%�T�< ӹ�<@rh
N��h)q!AJ҇R��8J\��
F���ꀡ�B�Zi��4 j�!ki�M
�B�dMR�#T�}���z�jP4�-�}�%�k*����"�v��6f0"=�4�}����G�Jj+L�vf�kl%�:�}:�{�5�[��<�h��33J)̮~���M���u�ں1�1~�#�_h�����=��㞌�y+��F{�6߼)[�đ�'���v}@%&X��ǅ��5��V��B`Np��S<�<����Y.5�+f�*;��C�v<&�펉��|��|�H���񒃷�0�����D�]�՞���e��VX��.�K}��[�����І ���98��W�^��N{��p�}�{!�6z}1^�WϹЧ~��<�C�}J�We�lT����_��3���^��8�=��P��+��:��cޟ����S]��Fyq;�]�gl,�/gg�aǤk�z�jΠ*�w�D_��́Q��)/Ϟ�]1��~�5"�_�L\\����ݗ�0�����s��fLq��)�������t`�ޅz�!��0�@�"j�$]��<�hW���423��2�8�:鹸���R���-��bM������Q]�wO��L�p�B��r�GKӾ���"����r�<g�S���kr����8s�ݙ�q,��U�[q&�d�!	R���Kk~�tt#=�g��c����Ν��-J��N�}o�8r�:^�[G+��܊0b�`�i���wzY܈"\�;99jO����Y�"%L�1\ظ�$h`����&�O����(e�8��FH���Y}���M˹�.}�	��r!������r�����JL�hV5�x��ol�mp��$ǆ�F��D:*k�&&C��<��d｡�{�d�>}�%35K�^?��Qc�H�]jv,�$�Z�}!Lğ�!����{���/ى����D�;4R������*ߦ�(9�Ԯ'C�bV�gЭI��C]����`$zc!vMdߑ�H���Xg�G�^�3�ڇ��1��(;�{��V�k��ߞO���T�E!����Β���TGh} �?��3^j%Ne�[����zv�3�q�eO�����Sʎ�Vk�GE���9�V��j��2(�����5_��c��
�e�K��EZZ#gk����4�૎�}p>�d_��r�dd�ܟz�
�q�93b6�M�I�ޏ\��i��tt�Ä�	�����L����Z��r_9�Z�k�ܨ��u�}]}�_l~���o:��ᆫٵx�j����R��`�QR�lV5�yTL�����@j5�"	h+�0o2O����T��_�/��w_b��c�xy��x�TE2(�UIW9u�p�m��yq5Rj��J��Z{����{�=��E9�$�nǊ�Zriqd��V�/�3}'"����ڱ�յ��37"�s'������`9�{P�-91Gno2}�%��Q�@�.�!��t�l+�Uq��K�27�=#��ZX������l����;u�|���ؼ^��u5�N��"[!�OT-ϕ\��i�N	�X�'tY���}�vCת�.������`?���prc�k��S�`3;M��n���SM���y��;�~��#2 �c����+�1�]T�/]L�-��c�����V2�z����D���1s$l�6���.A��[�����Φ�Wɴ�8ʏ	Y��6���pO�߿J��y~�DG�g�*�/U�Xag�wes�ގ�y��Iq<��ZtݣR��	�7���P�)���מǧ�v=�
Y��n�.�;��l�[gf'��f�Zߡ75�gG.(v����K=�M3��σ�m�*��;�g�~uގW�պ �/Z����1gm�;wJZ���g�{Y�� L�Ot	�vF:Ǎ�������ｎ����,vw��F�T��z��D�������α����f�I���L�&��P���K�Bd�t*���#W�t6>���,��KƼs&X�Ih�!Q�.Lr9/\xtǛ���27A
=Øv0`��9�j�;6c)�E�[2:i+�$
K���~lἎ:s��סƊUʰ���Zp�0�u��d���ї}3c�m�B��VGbOlG�J����r<���]��o��|�o�}T����b7Y;k��ZP_Fz/����P.�>��d��XLV�R���cNr�Fj�[|W�#F6�7�o�k��V>''N��^v�/C��|���Vzii����L�����WNu�Ǳ4�l��/uol��g.�l���b�O����R��.���o��a��;�z:0�1�扏�,9����$�� ^
K����A�̝�'�cp�L4�*��޽�s/=L	���.:Ƒ3�r�^�C��,y����
H�d�۔�3�v��Y�:������<���f1N�(����v]bV�is:q"Qc^���7�%��.�J�%��q �P��P�"y1�YN4a�r�"�߫Z��>��Ε ����h�M>��������|�v�٘��l*$�ŹIq��dl(قk��	v�0���T1�C����\sk?����=A܉]�~PN��팄��-��+���s
���`l�^��u�*�Dc�!��n/D�>�4Æ&f|ܑ=����y�Y0�/*�(eɠ��<�#��r�[*j�t��B_2e!,�{$K�b�e���^Ї݁ju�^׽n-�*�	��YS3�N��z����rX��p��G������c�����I���?Dq4f-A~�*�mG*Tx��܋��(o��7�x碦P�ܿY;�n�����~�N�D��̙z��~Bo��S��<.5\Ox� M�q���3v�w�5���;�f�VDs�َ"�JN1Ƹ㔖z$Tn�Oؑ믝��6�c��������:��n�;>^+)	{�Ⱥ���5�؈�hJɍ3�%���1�ީ�9՛�vi��g�gK�:����N�V|��Q2����NB�삥��PEM�^��2~p��>�L����8��j�'ތ;�Z}Z��5������3}@~�zh��%�4nX���'N��L�Ė�h.�\�UՀ��ݬ��Z���61Lѯ�ȋ�V�/Kc�%#S7+YԢޥKb�EV��zsoOq/���j@[2I�����Շgy�v�\	*Ly۾��gJ��֨9k�Q:<�qN�zહ���e`��,#������v��9s~A%�p~��D�hG��p�0��"5a���(����=Q����/�>n,����M���,���D.�3����Q�̣~~�=��~eբh��a��E��Ӣ�{m�Kz�k�GE�Uٵ3
ݼ�a���}��Ľ�X6^��N!q����w �1)���n������=������������O�lpp�ZN��?���Υ�&<��ށUҷ��Y�t�w�(�fë
	�̯M�2�����)��)���I<�Ŀ����fZ���kxcU�6���0*+��}�� 1����>5C`J��'#��FG��51[���ۗ��[�01���>c0ĸ��_y�@ȿ����i�Rf���cR�ާQfErɉ�D߫w�l~�i�}��P�o:�|%��)� �b��}��r��R����}����"@�[����!��uO�zg{d흕(��y/��n���h�0��';g��2�Xm��w�K��>�殗,��cy�����ͻ8��[�G�gv��S~� �T���z*8Ư;��h�=���;fn���cՐlR�m�Wo99�r���=v�#}CZ>9�B�����G_+4X�V_�AgD\���褏G���;��ߣҠ̸ͻ�5K�R㞋���>r^�l1�����C|��n�6����QJ�߁�Z5�^�D�;L+���#މ2�N-&�!�p�`M��͠�W��4ݞ1~4W��q^�O�&;Y=��~&��X����=;QT�������}�Z����U���q�`�J�����a��-d�X��Iȏ87�J�S}\Tmk{�zT���l���$���1#�X�*��x�w��6V��v�?K6et�8�;����<_�ʩ���xE��
>��j-\)�<�&ڊh\=�%���Wf�n����=
�қ�5��C�������,�.$��a��ۃ����xs���ٯ"`,PUǸd�>�Qq&;ȗg�Y��,�2�����){��Y>n�fS0�ŝ�!��id3���w]���[O��iQ��:v�j��D"���Y��ɫSh��
��7��4e�-�>���V2W�����ϫ��f~5�}�Y�)�?G�M`R���*�,Ǟn�T�[�w��K��'�N<h�w��7��� ?�R|�Q��U�N��Xc�=�7��q6�gA���Y�jb��K���8Tꇜ�������AY����;�-R�/�hB��}�� ���.��	B�^��}-e^��t�n����~}��q��e�3��:T��yU�\�=9�E�7"J�P�(Nu��=��3ݰ|&�x<D��pǬ
J��\p<]����3���gC�6}O��h���Ω�$>��KȄrrC�W�U�O���_#��ʳ~��9�H����}���fЬ�������w���*V.:��x����Y�a�Sq��4��>0�rY30i�۠%������g�\xF�s�w�;8$P��$�ɶ���'��mϪ����ku���6\4}5�\��-;�C:�B�)��t~����f��� �4>G�|��_u+�][���#��� ���8��nfM/>�)]�\h�M؜�~����{ü����u�fC;bg庢��b ���y��Ѹ�PQ��{����aN̑�N�T"�p�÷�z��.
2�g;r�	kX����>4evvh�K\����:�7�x7$SP�*,j�:ii���*zD��5��8U�Ta=}J�M��Ͻ�g�.+MM�m�"8�`o���C|�k,:�/V�;tT�\b�ڼ�(b[����즼w��~�!oF(+覹��$��3���S{�A�Q��w}��ށ��\&�\�OTF�5A8�aE�/���j���I���8S^���Ql]_2���[+�dL�uI|"����P�"n+DB�M�Nc��6%߳Q���	z]E6g���2�˨�)�54�����é�]�=3qm��>�����J.k�[��H5u������SwLd1�[�ײD�j�Hq1�O�����t�G\U@�*�/����M����DOA5x�+�����|����>���͘0����
�7�E��x�fW��NƓ����s`�Vr��#����1����m��1���G�<*�_wK�&�D��Z_q�ay��F|�ƃ/��&�O��fz�p$|�`�ظ�Z����� 乵�l,r�����[��g]�.�]7���c�9%8���4䚈ʾ�}�t@:�N�G{��}����:��a,���y��	2@��s��,Q?x=��{0z=97{����D�n���GҨ��*Lw6'7�;c� ���D�h�F5J��l�ё���.*�	�VEN�7�k8��ɚ��:o:P�/���ߑW��rVs�c��6֚��a�����35�SGL����ݝu}��d�qq:`�Q��6<2���s��Ta�����v�E�G�-{6��0�<��Kʞب>LԀ�2�ވr�\1:���e�m�s�M��_ٷX{Է�qy�Ȅ_�7�ڃ��)��s��&d�=?R������M�d��^7��y=����ٯ򈌃c�	s�!�l�r[��i1e���騝������>,,�e����Ftq�OT[�u���f�5�c���Dҗ��"���lLU�+�ﺽ]c�i�}Q=sM�	S_c4����7.g��D��͊��S^�f�{I��tF��7�x�c��	��]b����2��>-��l�%�7fO��/��S���"�~T!)�A��g̤���O�0m�C畟��ufi��:��ڸNA����`@�9��{'"���ش�}Q�+�lZNb��۱���E��q3p@�ս�4J�k&s�g
��2'/k7fuZ��Ľ[`���f�༡AM�ꣽ]Ρ��]��I�[P= �軔:	W���}/����^*�������ϛ�f�GG�E[��2Ⱦ^���Z��m(=c-a٤�F���؅6�j�;�*�p���I9���뮵٩#�&��v&��͟*�����_r���G�e���Kt��8�<&���ᴿU�� ˶�Y4C��>��=�����g�/�kÅ�����JNu�d����$��h����r$1��N�D��Wzj@��
u���g����NsY��K�qGu���y�I`�35]�9.��1��8{8稍j�Fn�w��+F�4h�ГJe�������&�v��v���{^z^��P�C'�o1��j��i�B����j�x�����()���e��T�͝�~��x���E�N>�]�+���,���� �H �ڦ_w�:v���O��=�3w|�Ѣ�`�d|��zˮ6�V�"�lս}P��#{t�叱��$�F�s��8��7�-�j]�8���5�q>�*��E�e�vX؅�J;C�yj�������n!�Kݹ52W�(6��%Vm����Q��ֶ�j4���d�ފb=�(L��i���dp��ᎪpOl�qn�f6?>�;o����fߩץ[�X�?	�����3ֹ�0��,��Oy� ����w��M�Z}�7���@Yצ��2Ȕ�=hL�9��Mh�喖�'d�Z�7E>K�Y��&����#q��b�B���v���s�%�����d<U%}�ۚ�	�(и���2ca<l�%������%�+q���9��}�'$�ϐ�ruN�Z'�b�S��7{��t+�;R���P.]����{�u?[�@7�ow����d��I}u��w^�������[=چxy*THk@K�]O^3}2j�Kw�Z��'1�iƲ�.錧Ƴo��O\�,*�b׋o��]���լ��k��G-!;��۾ݾ�uSlȯI[q,�]h�����V\�{}��)�����7��C�"ȃ����:�7����n�(.����k���Z�땢pg.����H� V���q��n�rY���M��;��7`w��H��M��Z�	�/�����
B�h
�c̦�hF��(���i ��(������QT�J4"D��IJ�4-5B44�P�AK�44II@�PP4!IH�UP�JV�R�i
V�
� ����)�A�(
�B�)h(N�@� CKI@P�RR�-R����'p�F���i���" �)Q����+Ξux_>ּ��6?3�/_V�%�]a@��:Y�n�;�_����������jVm��w���#����*�g�L�� 5Q�2�XP�g�UNk�LI�3V�;���o�lM��z\����_��m�
X'�����HS3֩r����П+,hq��Je���D@B��xf:_�î*��=�=��>�qZ��_��Tc<~����d>���}�s����*K��n&!���4���&���'
��8�hg�uc�7�c�3/�w�����qra#�"��Y+�`���0���(������z̿��ί7��0�u)"�d��f���H[4�9\��p�n}�}9���n7�$Y/���>6%/踍;~L��B�*k�ÓU��xh����Y��5��am�q$�jAbT��}��5��x�>���*�J�o�ƪ��{�+��s�w��pz����Х���]��q⧬9���0�ۛ�y�rNtl�0�{k&��J�G\j�����p�T�����}E`�����{�����,�Ƴ2PD��mm\ô�Kh��(�w�4�*��n쨩Ѩ�g^s��j��P�KN�����k�Yp�~���`B�⪥����7�TPj�c;"6�Ɛ㲮�Nx�X�q�tg�#3����
���M�;PONMBٿ��y�~�1�q%�,�����{xL��F�����|g7�n��p�`Lq���,*\X�Tc�k��q��j����Ts�iv]w�bO�3��;���ه��ub�WR.$�O�#M!/�_�{�S(�C�\K7*}����&�9���]c���D�@�=���#s�T<���3�'�d���}D!� �7� ��n���ˑ
]C��k2�"A�����E́���\��Y��=��^�d~�������}��*�(�E�^�(���=N���/��p\r��tH�5Ui�)2f1��r�=e����)�ɍ��y!;�1��g�M�ҙ?q�#]�3� ة֗*.z�E�TО�U�l�W��j��Ò���08U���8*��dȿ"o�-��yȝ�S���|��]����S�c&��U��z���9L��ez��~��
%MF��5�s�:r����I
���;�䏞��wI\S*��v�����z��jZ^{�g!�Ռ���?G�e��=s��S"�.x%�#��!Ƒ�i]D�BȊ�܂�$�(�����J�yw}��+b�� �Z��H%LT����rܜ��׿m�$���h-s�����v���;6c��Eֶ:�Ԗ�1V�b�g�K�|�����6���O�=�o%b��g-ț�-���/T��V^w6ORۅ����x��Vl?l6(X����:�?->.�I}�`e��e��.��6v5�a��3�����/ez��3�����!�}Y=7=3|�f����a�}�
��q8'<��<(����k�K��pr�K�M�z��K���6=��H�����E�on���6%�9�|=�µQ�.ש"}�����m�wۯ����`/\����.��Ϗ��38�ɴ�崚,��hq�x9��y�tfz)���ك9<u�^1�	��S�Ԫ�Kս����gy�>�UL�x�Ĵ,a�#r���Gd�}��dL�C���8�v���݇F�a�ڐ�ˉ�f>�s7	�"e��txQ�����H-mzs�7����גZ*r�� �{e�6'�%��&v"��4&�h�MQ��e:U72ߟ>kn�f���B��� h�K�Oج��y�`=m�Y��"�k�f������r���.�r�.��x�^\HSɚTg�b쮢�sN�aCN.�ͮ�v^\��D��ԕ���w�ս�w1�r����WNT���z!�c u��Ub��\��1�Q6��<(O��]��_i[3�0��.��^�^*fLm:s�ZØ,8��Q���g�{^�+�����}VT�"p��&r��%V�|���TH�WXĞ�����:�s��3q�^c5�,��Ty �ɘ��>�C/��S�B>��ŉw���O-������aľ=�&��B�#QʼX�U;eI���I6�,��Q�b)�{]�l`s�[����&{ȩ��ݧ��"�j��d[��3�AD�Dya;�<�:�g�x�L5S�Z���H_�r�6�'��Rv�L�Y����Vj�y��7#|3��խv�{2��]Ǣj�̚Pu���W�(k���\fF�4_���U���E������x/XqF_*�Q^�@̿�\�1���#�9Q��k������b�3t��m��^��*r�˰��Nlu��O͛��93 �=4���H��M'��������C��gM��A8Lu�i^��(�S�)��J T<v�7Q���>�\����/ws����N�=��cU�x����*3p�+)��oy��ؒ�X����ѧzW��cɻ�7Nd��?��qQ�������oF����lTԁC���Xg��}�4
�~��~uA�(�#$��&�Wq���81+�+<WlH��ؑ!��7��Z������>������MÞ�j�A�o�� ��މR��'�+}�'#`/.��}q�㷌�q�%�x��)ɥRT�����L���V6(32��Bb�dv�Vg����'^�S`����״$�� �eJB��C	��ǌp�yA����ZWN9���(�
�2�?,׃ʟ�^*ۏl������㕑��v[�Rꀗ���_Ȕ��D۫�C� �d����3�;=Vrk��Y��[��<�������p�\Llq��a0�m9��&�>�3���uQ̋5��{Ӡ�zߩ�3=}�5a�$ߤc׋�;�/�7�5���(���ў�w�bFW�z0:�����f3Z��1q����2���r�Rm��F�����^{�����L�ꪅQ�2&���Y�\��K����t<�z*Gf�))��ь����Z=�}�}��p�u�/��Qn�/���P9���Â���n%�����Ffw�o>�O��A7F����8{�={�v_w.h8��%���3Y�p��s�NN��'��]����
Ღ�� ����V�x��q�m�+?:�h. �n����m0}4�~�G��e�=7�v����[%���>/�>����Li���®��u]�2vbDw2{)��A�\虍��X)q�x�|ZC���W�U�/%�ӳe����A�����7>5"w4v��>���Nw��4./�o��^<�����E��WJ�J�G���,;S���8��.��0�>Y.OK�\�Q�SG
�C$/OT-�P��:O"O���t35�������"_��
�"#��	�YQ�.B����ě��6E ��N<�7�w]�2��p�pύ^�ab��7�D�qCYC]�f3D�.�s�:O�<��F�F�^���ja�q��<��6�uƞ��5�1-]��u;��{�n@�"!�U��s��r���~���3� ��r�,����H$�
.;��6]8�J�1�O-�r�y�}�]�R�j��2[\��ܫ��4Vзr��ls+�P*4�+���"Ff�{�b�f
q��Ζ!���K 籖�57��Cz3+;E̩)k��l�{���Y}�2*y5ٙ�* ����#��V������⁔�3�\&�����&֘
��bu^���Qn��s�a�`��vt��L���Z����ޤC�f�I�.it+�.g{<2}�m�����b�N=n��͚�>�|ZJ�f�V�O�z=q����c*6����'���Wx3.<��cHPΈ,�T�LEy^����3_g�+W }s���7�ۼ������T0rk�(K�rrBߩ��Y�p�#:��B=4�����B&�e�ߢ{'�p��z7ѷhu�S�
ؼt���tM�+j�ऍW�����J����9�+%OK���eB�Z4���]*�z�T��EՏ}3K��@����}׼k�_!2ߋ�q���-�v|����Σf�Ԯ;<	�N��^���:Yۥ����{�+a�2�Y,O��M!����c��6dv
znl����в�U��=5���p�O�ش��b^AV�e�m�Ё�`lJ=ʌw��7N/����&'�5KOз]���Z�{2�W�����i6A9��;�c��y~�y/0�e��ll�;qs�V�ed;9G���f.o��?
��:�\Xɓ�>��[�s8)�Q�2�<�����������T�ۭ��u���1���D��Òb�,De�H��9�ȉ��$q�j����9�$�33�9j��7�^!p��b���,�_B&3�:���T�rpe�hj������&)��F,3:��
$�f[E�3ﺤ��3U3j{.7�z���������>��e�i��?y��-��Quߝ�����5�y���펉�pK��~�N?	��M��f;E�?O�?�+�yt��t��2���N��Ǣk��J�}�`�pv�h?1������$Tw��$�����=㺜�0��]v���wC)�y*�-;ڨ���Pe�2p�����������4�>epq'���}��}~�#�����.�J9��ـauA��Bnn1A�W;lNp:=ak1�'Ź�8ì&��Z�v�S�ẉ^)1Z3��H�JY\_Y����)dƞ��=Fh�s�y=�JÄ7�;�R�����){�̵=�b�O;"����uV�{X7`�{(�1����~��MpԖ��������n�M�{��<�0"�s��:gr��;�{��:(^A�L��eq��xk��U`��w\b��������-����l�e�*W�Ox}.�w&��5�@���/4ެ|���?K���1���瑵��F�v�7���_O�3��wQ�c��܆��}d�])�Ѕ�Bؽ�_���+%b�����(����t��w5��w�E�}[�7?xhr��>�z4���%3Q͂�xÍ9q.v��=ӝ���5�o�!x��n۽5�ϑ�R��{�ג9�`鳳`�s�w�B{',�y�$Ξ�♺٨ax2{!��*PGN�;L�">ȍ�/��@Հ�t�:�zW�}�vy�M��I�-����S;��~4�f��T���[�����d�k�ٳ+tN湘u먥�!w!N!2�=��03�9����L�6*%}����4v[����dx1�b�~��e�[�ud�ei��Q^�9�����V߸)���[Nf�k�7#z�ɉ2_�(k���B�ގ��t�#�	�r7��j�L�'�J0{=��?2���c�c>��C:��|��A���{+P��������K��x*�w���B>��A/DQ���Vi�J����)5Sm[��y��5�,�E���Q��[��Z���9
�`��s��֎�S= �2Lz�j&�7=M��?~��s�ߊ��zh��D
�a=K��Y����u�qmf�Su62�����	����K2/�a��S���5�qFpTq"kU�y [�{�n+&��j�_���G�����&q����S2y]96�N�&91]�5���u�Wz�=]nζ�s������7Ȝ�Ə��ٞ�C��c���&wmg��#N�eON\���#����r�q~.��5�u�+���Ρ�'����p�"�gq�x̔�9/w=/�Ӆ���r����n��J����W)���U��}#*x]B��f�	j]K����T��P̝������A슉扡+v<W���xoz�O����.����%;�8��^���F�ћt7>�W�&;1#�)���匞���Y�lZ5���!����Vv�mcª4�	Tu�O��С�=!sv7����bn3d�ӣ�y��^s�f���\��܆&:�I���i=�&{V�D�s;���N#���UUU���&Ȁ ͏��@@��ֹ=� �?C���5�>�`s�������PD��{�;��ϣ���_dP0H*?`b�C����!�B%b@�I��_|�EN��T�̨�% G�J��U2(�!EP?�Hc���k��;}^�	���Y���@y  ���TC����z�������<~]���?�o�Xt���~�Ȫ��&�*"��"���"��������(�*��*"��"��j��h���b���j�j*���&������**"*"*�*	�������&*j����(��jj*"��"&�������	�"��*����**���*�"����&���"�"���*"�����������"�����j"��*����*���(���"&h�&*&b�����`�"������������b������:}'�/���4Hp��/���������P!�,:'�X�4��8'��;?�RLDET�Q��4�AHA0�CI%%4$ą,CCB�K$�CL14�5S0�MK%$�1�D��ғD��1+TL�1$�+0PA0��LTH�0IA#2LLTT3UMD�UA!L�SIAA44UT��PSQ>�^��� �)a�;n�>~(o��(#�P@@���UUA���� �������u�����a������_��Q���8X�o���_�Șj��9�����?ݿÁ�O�{���@q@���O�C?�{:����B"�����D�������0w�����'���Dz����x���%�k����@�����;����s�:4�*��"�=����[" t�(�H����C�hc�{�Cq��N����O����?����� @�<#�"���E��C�(�?f�n)T9�E����PV�5����J�2Q@��>�r>�}�<WtZ���1�� @��d���~���~^?z�����_�	�Nx���o\!М(�xyߖ����[1!f� ^A�2���T0B�O�p�}C�� Y������2`�.�	
����������d�F�@ {�� @�O���ۿ��5��8l� ���*I 1$#�	�PHH�x���f�q�~�$����G� G�DQ��E��0�ȟ����{���s��	<sZ���n�؟x��?�d�;/����ק�����P�
�����'�|D���� �������
O��� ޘ_Հ��yvf z��h��d,Ҁ������d��?lA��G���~���?i?�����D;��(���h���v,��3l�"��vr�����	�/�(���U)(P

V��T������Qh
JJF@@di PB�
E �TR�h��D�UJiP�� �A
��� �hUZZQJT
�JV��Z�iQ�� i��E))
QA�)
A�TR�R�hJR��@)�Q����V��hEi)(JR��/��/������Ec��A����H�/���_��!����|_��QF����A���A��pŀ�p���R�S�
�o�Fn��Q��=��T��_�"�������� �?w�!����w�rB�>�X�q��?���{#��G��������A�c��xߧ��:D����'����,� ���)���� ����B�ٿj"�������������~����I<O��O�������OD�~y�����;<	��L	��?�2'���"}�O���w$S�	P��