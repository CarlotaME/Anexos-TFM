BZh91AY&SY����ߌ`p���"ߠ����  b1��  '�^��M��[IX�UjU��3b�"�E�j��h�mX��m�͵�����%��PZ�i�kTl�0-��W���Y�PRJ��"62M1%m����BZ�M���f�%B��#m5MV�S�}۲Y��T�Y��ْ�H�U��֕l)�Y�5��y��ڪii�ɶƥ�k)5�ɱ��R�2m����Vխ�j�(���!��U�*�إ�2��LXj�KU��4f���j�2����n�i� �x 3^��i��X�ܦv�w]�j[�]KkZ�j�n����M���;e1�l�U4l�Uj)���nc�]�f���mi�6�1*Z�i���&[�y���+����NT�/N��JP�K{X{�$T�����Y�ڨ+����y��^�U����^�E^�z��R����4{iK�'�}�4��;��/h*�*�/�he5��vݵRR%�� ��|�m�s����}��{��ީ��}�J��_��k%�/�}5
�}��뾵RN;���b��[Q>��`-Y�G�}���II{��B��PѼ/,ѢT����ֶ�JkU|y�R������7{GZ�v�^򛮲����W9�=*�:t��xn�%R���ޏ<��wMއ]�#�
�)G��ǃ�%U���V�h�xӭ2����^F��hڶ���i�V�"4�#}��E9*���[�E�IQs�^=J:���G�m��.�]�	������6;M7��s�=*�̹��oy�z6���W@QR���^�z�s^�JiMR��l�����J� �}Bm�umw�gy*�R�����������{J+�+m�������j�w�7��v���-[��{�Kwv�I�z���SJ�΍ХR�i���z���6YsԴm�TiYB��[�ƶ�� �����V����z���U���E(]���Ӷ��{��*Q�#q��6ґ�w�������*N�i�H�欋�yy�F��z��StW�ɭ�KL�bWl%j�m� s�����o(����� ^sӀ�{ޣ�h��� w�M¼�:�L���t���Ѯ�7S������ڐAf�C=nՖ�M�mm�| �ϝ}ۯA��z+���.�QU��N�F�*罧�ocѣ�]�+C^��`�v��S��^�ޫ۽(���q�`��5M�UX�J��X�EI&�� �} ���z
\r�Eǯv��������=�z 5��k�Z��L�X��N�U���.����        50T�Jz�@4   � ��ъRR�0�0 &#M0i�O��JU5M6� �&a1*�	*�4 C@4  �?!0�R�4` ��  ѣ@��D#IL��Q��L��4�6��Q�z��=���4�����_�d���L�/���ϱr�φ-��^����~~Flm�o>����c6ٶ�6cl��l�~�ͳm���{�o�o�����o�lm�k?��UU�=�fٶ�Ym�ͷ���ɛ��m��?2����2lߴ�7E��D�a�a�0�����F�{,f=�0{&0�X�{#0�Xa�e���`�C��c�67��c�l1왰�[0{-�d6���Xa챘�L�{,۲��le��{,m�e�m��f��l��l=�ɰtA�e���c�ll��7�fm�c�m��A��3e���gDٳ�f�{,1����A�ə�>H�ɇ�m�E��6����m���m�ɛ���od�챝�g�f�[7������6�[oe������?Kuo��o�y���~࿐��ޘB̬v?�����9JJ�D�ɖ�;�+&�F��tR��]CQ�	[�F�v�L�%q�e�֐b��+�,iݻ��#��6�c�L%]�;���"a�%�:XW.�vWwA�fMJ�C�W2c��&N71���c��[��Dծ���m>%���hm�	5�I����]gR89���a�sT����P��:7	g#�|�+VMn�6N����7�5C���QoZ��q������)R��泤۽�w�K����75��1,�^ (���nʺ4�T��Yh���2�B5}��Ƶ09Դ�B(��y��`���l\9L0�ܑTp������[فU�q���‱��|wή���{��ц&�`����/st3r�gf���5�Eaml�ݎ
 �(Z��5�Wu�mCIQ��)�RX#ц���G$��19A���Y۹���m ʔ�#�A�-ذ�D��'E*�(^
�,nj݊����p[t�#��2`�CV����0��u5ҥ@̺޾�짶�<Ҿzz�N�I�
^5=��49n�$�n�7SS�Z���D��hri-��AG:7p�|S�}'je3��J´�u5K��+b�)WWH�b}�4��LC[6�Wٍ�kt_:�(5y��1��qP����V%�b�e=4��-�'t�X�K�(�ًe\�V���؀90�vM��z�D4w��ƅG��,�J��Yo9�k@��a]��mOC���Y�AX�^[�n`�S�4�GJH�����]l��y���
1c�CD�M�D�|��	��K#�uleH�4���u�r( �R9�0�����Y(��S�V����Vc��9ӣ:�gS��k0�Yԍ*	GvK0	(V0�^�H�-���c�+I�P��A�ҙӴ��[MGn��i�<�ܽ ��ҵvh����s}����P{PS#!�Vŗ��%��n����`���s.�a[P�Sy{�Kz�1�&d�NѼ�S˸R�]M�H��;�X霷�H;�^�`<�B�,QZt��AP�b+U���-(���+��RX�#�HN�#��2�5��9�W��|�9M�U�3%��u9�}3b��� ��J�е0K���Нw��'zv��N�A����.4�,��C%ֻq'��W*)�ĺ�Qp*���[[��Gre
?k�ކ���5uU�2%3ib�B�T�M:�5e��#���C%�)t��k�>�F+I�e��X2mb��"���۵s	8�m6���C	��`��}a��x��h�b����U�NZH��2�i8A�ځa���go	�]���i~Q����lVSˤ,�X���6�f`�7(]2��+��xpbk��U��,8rJ��e$*m]�������YPSmQ[�2�_%�V�]�Yn�IB�U}c0̱C���	H�t"ذ�^<�.l9Y������\�;c�覈/���
����U-n�j�u��N�ռ7D�w!�C v�hO�sr�#ʎm$����3#�k��i�ڼ{���������{CMCW�l-�Y���o��{́w|8�x�\�.��)ˈ�W�u�l����֦���Yf�z&Z���3x��F+c�V��i�e���
�"�O]kٔ��5-��V�i�kP;9l��m7a��9IӼ2�*�b�sE��KV(L��$�W��3.�V� �T��+/.��e$5�n )��VqT��ՌIf�nb��(�<(�goTA�Z��_oa{RH:�Sp��2Эӊ���{�^m`�u�o4�ui�M��O�n-��X[�q�:�c2��%]a<�aR�kVcj���{��yA��H�b�
�kD�sи;��Rғ{F�4�I��`)��[t���I��3��w���3b�����9����XC�+�Kॶ�6�:�Y���"T�0�4/6���)�-��,ă��)Xj�G�bp�%�djKh�ZJҁي^0�̹`��&�YwBv)i�Ov�i9A��*�k�Y�mM����dɧpcn�)�f��R�*r}����oZT݈S��"����d�n�9����6k����z�f[m�K�\� !iEm�f��~sGpa�K�ՉWk*��r�;)�׸���Fc(Q�Osa9�(E���rW��J��o0�-���ұZ�T��p��0�0B��X�x�.-�s����Ob�"$n^M���d�t��׶��!ʃ1����a��zK��*N�R�zӣ>�8�R�YÖb���<CpԊ���[w�&�7�a�̛��:�F���C�YO:����\H֒�g_+80�h)�|����3�r�*�P.��P��7�Aǈs��Z���̣f���T���M���r];��2���C�-a�"�����nn$���J�M8d�h���Z�]�t�d�(�ݎ�2��_!�2�Z�xʇ���%I
Cq�Y��Q�論���OJ����G��Y[J����㯩�CZgPy2���^[��ǲ��-F���ӊ�k3&=;`î�kOg4 *:��컮�R,ժ�Ɨ�nS94>� x�ְ6�S�ip�bn����n�&+S����v�`6V9��OU
���g�)*y{�J{Q��ы5����M�j�n� `�V�m봝����..Ы#VR�En�k	A����9��v�q��{/m�%;\; �h����z���u4޼��ǹ�!����$�nV�s�sUi0�ۭ,�s4̦�Ա�6�J ��M&�^�V��� 
���IXS�L\{B��\�����b��%]���#�Y���$��x,���n�ǲ]t#�+Ǳ>\i�	�ۦ�MT�SɆ��B��V�ʫ����f��ꮥ��j<Ώ�k8�j`�VC�8�7@��拔��	Kw�IqF�w��C0n��5�q��WH��'n-Eh���e���u��&����/#8�Ԙi㬱��*���;�:��L�˘���n�²]MEǪ����n��G��-��tA�����0H�*��T�����U
��u5f�ɧ�_$(��{�����4�:� :�":l!�ƻ.�g�{�t3/i��.�h�#�f�AǌʗJ-�mk5$o&�(W�>x��x�`�-{Wa���t���q���yf,R*5$	�94֛XRUV�e�-Lt���W�COD�Ov��qG7dn�5�.�Y�Y�$�ԁ�JK �n�PS�z��L/l�o�i/�����{kr̷+%�Q�7hS�'R�cq�Hw�]����W�-,��>p�짌AY[����a��D4�ЊZr�k��p�`�$�v�b�SJ�Zm����x`��tˋ�Z�{1�&��4���<��0��C\#����m0���c.*��wR4Jқ+\��ۮ��=�N�ŔD:R����L��:�[EZ��M���*j���)`���� Y��_%u��f�앵�N�?�U8�^
�J��h�V���ϙ8�*,����{)_i�0��A������K*��94Jʏh˃-L�3��&v�G&$jf7*)q����O�E^IC���&�}5/�iX���sk-�{����i�~HMe�ܲ��nR�X���e�&s�i��P��[���C�IK��G)��<	�(�����7(�� a�{���=k:�qP�H���`hojb�B9�H�`�{z#8�|��uw�R57�S+:j�u��[���h�T*�R�D�o&�h�ѥ���&&r!X�g6�bh�5�S�wa��痶��#Vز"sG�^�q=�:�%b���"@�=6ZJ�������87Ob�7V�J|RO�,ņ���������	K�mlඕptp�"�I�T]���m$�o�kS�ư��v�l�)Oo7�� �ܫ��V̦㚧*���X6�˴:�&�P���`� �W�%�=�Xԭ��.�;�5�ܨJ�т.��	ԝ��]�8����}j��!��䣒�"� -9�*ĝ����HN\�A@@����h�AJ��v-1A��G8�e��>f�#C1�n�X��n�Zu��|���n�r}�M��� qL�/pk��$2�J�9�����L��+l��5��GU��̤�d-��'̀k&*{˴��w������׉���j�"�!�C�1��B�H���Ԃ�x�[L5���	�ŋs�j��xs��̖3{n�g1^���5�G ��	u�E�w71�Ћ��1f�`-���	�h�WU��S͎S��c.��;֡�r*j#x�V$��9��ۏ�d3�)%I���� '��U�o�M�_ma��Au��p�Z�/�Z���
e!�2/%Mm�6��3D�v�Rȳ(% ��+,��]��F�Y*(������8n��\H�:���y��
�K%X���^s����iM�k�:��2�Ꚑt�V�
j�-�Rޖ�1On�n�tKyq�Xq�6@�V�Z�ʹ�}���5
ò����Ǧ�-�l�].+�e�b��PU��b�}FA��IJT���lt��:�q��b�3�,��6%A��v�,w����`��b�VN�
���b�z���vq(J�Wq�S�!�#������p㷒�m��ZN ށǵ��~ԏؓ
�Z��7���ܦ�a��)th��)
'%,Y��F���\�[G�)�UB�����r�� ���m�w$.�8(�{��	N��z���H�=�c�$��M<+q����*���(JwA���fb�&�;�sv
EI@��u�sU
	����Ӌ�^�<��0��j@Pov�V���F�R�uՓm�a&`�y���Z����Q��z����V�}�|��ʳ]<|i'Z�5`⼠;�G��Ů���aG�[۪r��V�T�|o$9u2O�����{oq�z"��v3nn\*�#��X���s@�Y"�ڷf�d����Օ*�CX#�G��u���� ���`�� �Qۣ�Qw{�9�����%S5��h�(��i�/� WD�t���VY9&q���m;ȇ5r�_�mXl�5ǒF��_^,L+e֍�z�wm�|w/���v�ޥ-Z(�T��.�1��̨���өik737G���[*�:�O�{q�Uu�gt]*2��(3([ak0g	r�nj��ֵb���p�M����C��#e�ԝ���\ڜ('F�Ϯ��4iܩ1e�l�R4���]E���M]:N�l�@�����T�V�ھƫÏw ݃]�&^� ���]X]�,��C�6Mb\z�JuەИ��ɍ��l8�� W���a8o*��i�Ҟ����ӊ�6g�؉�m�ٴ�]Z=Z̝פ�b��Y.��snP2��1�e��&�i̽��3t-��޹o����n�.��Z/B�ӈX�M׆(�u�:���P�vl۴[�sE�yOc�j��hŵb��]�P��Y�.���#eh���~`%.�[�ш&�٫Trq�{�^b�*J0D��-��y��{i�M��m�$%o�Vf����)�3f̤�c�PwR��X��|D�� �5�̔�.�f]⧭̠�B�*vαDĜ�7f��d��a:��BcK�H��0�V73D֞;��C�f�h�[&��[����5V�fԮ�ޟ�1�A'��1�=�����A�������Xg`�E���۔ml�qix��45�d�iE�^K��J��S,��bM͘r�s)d�r�ޝc(���r����j��\��"@!���-n��ͭ{3�k�Ue�5�CJ�ٴ
��j�Y����;qK���$ �SL� ��f�uf�ä[40>�z�����<�����CH2c+@L�
���if�ـX�j���Jb���f�l5��'*۴�U��oiڈ7�t�TuhD�[��-�N)�^X�jn�R���ߏN�d����Q��"��=��S���Zmm5#��Z��ܒ�̫Ɖ��V]��n����&C��Oya4^	냷��d��kNS�I�k�ܽq����s�4Q��ƈ(��W�WBh�:X�0 �I��56��6���oȗ�!ʅ_E|�u��ft
Ҵ�l����G�$Xc]iF��v��FT;�9�6�v�<�V������sB�١����f�V*��0a����N����^��ըP���_fPˊ<�O��\�ň�k�ۏn��a�έX��y��IOT�2Ź[�t>�3@�ݦ�.
X�2�5��7��0����:��̸�à�8�-a��ǚUZ�X=��XO����n�+0���k��hU����-ϡ���\`��2J�KSV�0BM�z��0�0�-��sfՓ��ᩃ�k�EJ��CB�P��~�8�//$X�z��G���v��[�(�%/�������&9F��4��v�Jz]i5�Aѵ(��F�oC���a�;�n�[�r�AhB��7��wv�и��s)��w8�H9�!ʚ.�=�Rh�@tG���ݡ�b�DP����C77*u�Zs�N�K���,��ݺcx�[+C�LD�eaE�VL|��.;e���1>�C[4�H'O������]:F�ơ�4���Q�����6NM�\�:EJ��.�kro�	;3HM�P��MN���#0=�3&�]6�X��<���>��#/XoOεV9�F���W�FZ�d�i���_n��A�Ǵ������ $b��˼�vIb×��q�f���R�2*f u2�d���7a�]�x�*��AT��J&m1a�"��sTխH�{05X�'+/r$�銏c���u�VCM#uh�F�:ӵ������B$!��Ņ8�*���/���e(B�#*+����6>Zr�J��9L�r�%R�Se�)зH���N���0������L!�� �T-V�Je,�	F�T��(�K����)T'�
�*��GQ�\Wn�����<�g^|~��oog�ϻ?>�w�>��T��:��~JqvK�u�u#�VI��)�7/.pUĳ�|�f�����}�����w����WW�]���$�I$�I$�H����OsqIrI$�T�I$���I#�$�H�I$�&I$�$�T�m�rd�I�A)�KR��G*I#�$�$�I�$��eA�6�S�iǕd�j��pWuge����������@"�=s��
���M�S"�5�i�,۔ԛ]��48�s�iA��p)��+{���Ra	���������lBy5��s�;����B�
v�&~0��D����Y�jU��hRάݭ�%��=�&+��uz3b����X���`'N��oleu���s{���c�P�ЃhiU��eopU-����Z엞�s�P+g����53�ݬ�3��������7�.δ�I���֓M3��&���O'�MN�i��bY��1Y�K8�}�����}b7jU���`
�U����O��kL��c1q��ۙq�z�:\7]lL��E*�a������G�����-���i��;`�Ѹ�v*�\�{A�[�v]���-�T�>j+q`:8oN�Gqh��|�0�q��q���<<v���K��w��v�3Y��	�n�r�mL�A7V���e��C�i����hQJ�t�����D-�'U�]&���*ttn�+I�}�A�ՙ�a�4)�[m�7��=ڻ��Ij+%c��m���%��.���zGy)И/$9�kPK��@
�0�ʻ�q�Ⱦƹ��(p�=\o'.-�Z��x�Ϭ�[���:aVC��>�ޝ���@}+&R�-��ُ�p����R��t��>��wnU�V �n�{1CתU�"��t��%>�ۭ�X�����H]����4���1�܍�U��re
��.>�if���U�ݭqf���]l?CO'�&�lε�YkWIY�d�����`w���(�Fc����ّ]bTS�jr������4L�0l��@���|��5R��t��۬LA�M�r	ٻ�.���3�pF� (eYP�#0��r`��m(�uA��]��r�>�2\_^���;,�ŝ���y�@�ѓ�:�q�{67�u�2���H&��W�q�*D�۫��\�f�'�)�%�G4Q��"@��m�Δ��n�'N�6�U���d�#=��l��?,�s��,k\%d�S̒��q�먎�
ʦ�^h�ar��"Â��a�![e�*��0�Lո2$�o<.�47-��ԓ{�>ى�W`�xS$�\'�#�o;��<Np�M�9�]S.�� �U�M�M����Vj��"�����v)�I_7�.V���@){��5�ҋ璎F���lT�v�2���'A�S��Z��R���ڸř�v''l��?K�=$��+vA�*�9uҶ��۲���8t�/2V�q{X�T�lx�Gc�����q�YŲ���9����Y/�}nN�B�)h����\�3�>�u�����(f���5ʌt�L�ұh2��/�{K�
�Um=���)����P�0A�ѕ�1h�t�jƷ���
�d�,�&�^�Ȩ���ҳ_)m���)�R��m����%���跏�4�H`{-P�����S��H�7uČ&w����#�m[�f�2�bB�:��_�����ux�һj	c�c����#��ڜ3
�4�Rfr���6jK��e˭y����]؛j�gdrl��-�EV�v�
��㙴��73���*0�4�EK/� �b�{��dg�C��ݦ��Q��w�ڹ2��έQSH��i52:��ݢ�N��1�!|6�5U���ج��0]��э\�3Y��em�`id*�j��}}��XT����<o&7WY{f
Bq��	�W�J�]��.{����ᰤF��j'ɮ���ӬW�2�`!�W4m�t��Z��B��"q�9�Wn��z�M�$슆n�zr8(p7"u�������t�F�*���s�E�i��l��]Qs�J�t��l�p��B�BD��ʡ����h���t��L�c�B��2�Y�5��xn`|�%�7���87���;��=xԨ4��b%Z0�t�N�4�f���F�Ɔ�]]E3mる��*�\/i��:L���~4x��+����$)KK,^|�j��3��py�v�ې��G� �n���P�l�/.Bt��=Z��1
��P�yKV���Nm�����v܅�׃�B��v��;
��mӨ��Qo^f�c4.����FN� �����A��Jk2&�%�Gc�x�����Z�7zk@�+M&��ir�\w:�r��qo1^쩓�^T+0KҴJS���+R����S���پ�SV������
�wk�������e��2tr0�c3�������^fl�$#^f�1"�otRE��f��|�Ҭ�$)Z͙B�����uj���着%ŵ۰���J��E��!xo42���2��Psz��=fva�V�ތ:[wM���W��Zx� �l�"k�����-�Q�ێ(��ҶD^ٙ��wM;n���;W`����&�y$;ܮVJ��V�9y�HM�U��U�`������f�����	+{�����������ǵ�v��ޔW� 恵i�Qe^��)-�y�c*�	X�iBˣ�9���]�u���u[�9�y�	[cxLr�S���҉FwcE�V�K���釲���V��aޜ)0�ڶnʿfR��C;�P�t)f�k{�d��nNN�jИ��ܪ̎�H��^���v8.+T�w����icB�7p�B*����R��ɥ�
�u7B�ɴ�g1�1ͽzV]�����-���pնs9��/���M�]Z�Q��������/L�{E�����Ӊ�z$&b����[����Ǹ��3 W���C�IA3o��"0��3�=�1������g�G'1���g��� 6K��ع�]A)s�T.�F�n��{�І���K�ǲ�	b�����9g\�i�;3F�hw h]��!�.�dQ��5�9�]��V2�1��l�k��}7�,� %�ֽ�+�\�]�Ϻp�D��s��e3�Cwq]Bp�����[���Ѻ����MZ$���Qn�%fn�]GB��N�u�.�s�jȻ����bd��X�u��y��uB��wCc�]������n���l3�20����Y�]GN%yL+����S�aV��_(�]�Iv��x���|��>�2��.�������z�5�y�g��i��ż��h�dM��*?'�&Wo|�l�>6ŷ)E\�id����r�Uq�[e�;w0΅�o/J�V�ۜ2F9L� ���ªN#4�@���|�C�C��@�ܭ�iw�(��y�ʚ'D�'a�9|��ߞKH-�QQ�j �g��J��~�:BhoNe��4�R����iи�E6��,�@�c͡�ױ�я]���5r�3��)�Sv�+��OR<�kGm�����^�u�_SRzb�-�� ����Dރ�e�1��C�1�6a�̢����Hn�=R��N;1(+���}`�+�/�V`]u��e��|L�֓	�M�8������l'h5��I�sNGOF�x32��6v9��](WgWG���Ս#�hU�V��A�� %eb�S!��VP��^=�� ��$�t8m6�Hc�M��=W՚���v��ۖ-@�ZM��hV<��/x����@*c:��W��h�o�n���ϯ�9ӚA�糾Vko�p���R���Y$k��.�[�GS�)�K�s���H��[JT�s���)���0"�ZB�h>�m橹u�3qLo�g6L�=����Y��U�D��5$�]�q�<GD�	B��k5�4s��l|��Qt�/�]�#]I9���^�e�W��F?Hn�n�A8R:2fS[�l3���:�����Q%7�*�{bT�����K|�U,����ف��A�5k�I�̠��a�<����t	{�D�f�^�)�^���A����(ls��EvuN����W؉���7�����P9��ܽ�J��Y�ԼܮE`e[L�m+Ș�[X������fYW[Ĭ�� �n%��n�%�؛�+�[�e�;m:�f�2�t�#�-�1j��&��C����7$	+w�C�]>݅f��]+b��o(L*�F�R�fY�����y�I�{���A/(��s�M��q�`�Ei�v0ɯ���[�N�����DE%w$�9<an�&t]=�G:J|p���qwg8c��P�+o.*��굯U��hɗHbhVJ@���1���B�8L��[*��^�G:���,�G�E���E��V���6{T�v�,eN-n�&�ك3"͉�Q�5K�u=�M�P�9�5N�CH:D�\ݘ,̋����s�Orv�*m���iU�"5�V�u��sE���ERud��t��0+����VY�P��+T�"/y��T�NRh KM]U�p��4*@�g�׮_�8���f��&)A]�γ�[ւ�[v�vӔ楇�rN#�&���+e�	\p�Lq�Z�4���G=e��hr��J���Xq�V5 ��*v3½�h��{�.�
	�v�[ǋ����oҕ���}�1CԹvI?CG�'"�U�`�r�\i�R=h�Z��[S��k.��/�S.�b�Co�^6&�S�+�Ҋ��@.�]��7�����)NZ�5����BocK�V�艭Wn�*N��z�-
���k�[���,��z3�/"������L�#�G2�N�,���;9(��EK2�9�n��7$GR=r�5$1<5j��+[��t���e����`&��9��`�ƩwN0��[o������l�|6 �Zg*⾰�=�:-_VDҾRn�m�O^D��#p���^v�U�ѭ� ������o:�牭p�8V}/.ɬ�u�H����K�T�.�R��Γ��D��u��H��2X�B�:���5w�9p��P��c{�$���/4W^2#�`U`��p�ם������zm[���k!�mL��0��֝3� �������d��y��׻��Cn�T�O:����2�	��]a*��E�B���%Ghj�Ut��eC�K�p7��Z�/)���fg0^��Vt1���80����l�]��t�ʔ�1��H�⯝���7,[tؕ��19������m���:�q�����'�����s�8��8�/���oZK�2�ǽ��_&KM�r���ov_jޤ�ȥ�VX���	�."T	<A��*R�DՕC�n��x�kR�i̼�S���jђ��I
��ݭ��x���1^m�a��vq���a���9�0�O����L ��[��-���7yE�W����L��i>�D>Nc[�e�>M�X�xZ��Q��1yWd����aJ��}h�Qj���ya�|��ZI��L�������� �:�*1�Y����w"��g#�	\5��n�Z�*'|�9>cz�
Tç�����Nt�=�3���6�un���Z��tָ��m���Z���iۦenc�������,�k���c�f^���n�A��a[q�vܺ�7�-�!�����1��� �թR��Y-�W���)�fRW,`�)*Ɓ�9f��Xj)O����X���������Y�rG5��4�ݮY���U��m�&0��U����}I�̙�����U{"�+BY�y�7:V����Wo���1����s6W)Zq���Sxi>o��Q�\��n��ʝM<�Xb��Jx5��9���u���d�ܝ��˘�Rs��MPX̔ puFw���a�6��ȳyW�L������m��Mi�p�&����ʶmZ�w��������tǳ~ɻ;h/�IW5�
���k�4�IF��TB�^V��}�o�t"��TЛ2�W����8�c�?g'|l������A�����l9�8��Z>GQ|w�EW�:��ٱ�&�ȭ �����5\}x!�7�� �5.��9
����#U�Q�α����v]i��R�Qa�:n���7M�\�p�b+���
�;D���:��O��M@�92I���
�n��znp׽{�!�AF#��Ni|�!�u���RZ�͆�Ӕjj������-�Ү@ ��Xn���,����k73{U�1IMq��Mf�������cX���'�v{7��ָ��:�f�YǱ]e��ⷍ1Yǚާ3u�X�Nv�]��ڐEl�+��뾎,Xo6���I���,�yW6����]u@#fb�v�:�%7Z�%���L=Cm�έ
U�H�}���F�p<��Q&���Wk��pEv
�Ab[�]���789�CF2�!�����RQ�)yx���C3m���(hC ��/{.94a�O{�Pf�$�#�- ��`�-�3��\��|��Ҹ�m1@�=��N�=�1�pX�����&����vb�).F�:��ѳ#��:(��Rr)l��ǯ$#.��]�N����]�;�-okI���f���gp�T��i|Jf]�LW�`�4f�Yf,���C�i=��	�)��aWZ���t�*���:�e��۫�j�8Fch��٧(��o��z���5��]Ռ&���{��-k�A�YCR�7b�W�-E������H��L��{9R�kݾ�H�z��u˒�ϵѩ|�a��Ֆ��[��YL�:i����.����ˮ��˅gR�) T]�)F�G]�e��έ��ry��z7[qJ�̗N����U��5Z����T�.[-Ef=�H�T�;�>̑˭�)�TRJ9.oG#� �����Pʚ�5(Kî^c��I$�%��fv�+�M�+��.�V쨒mI$�E#��$�i�$�I6�$�nI$�AHV�2.�yB���a2J�c1\,Q4�UƝ� ��Tjad�ӹ ����uD~h����ͻ�V]��g)(����G�Ō�Ch�f�2?��32�HKmO/�Ml�`}.���uu�Ϟx��w�n�qw���l��m��<fm���{>��}}zf�9�o�A�W�������G�4k��C�6�v���¹_�%���r����n��
�P�vL�tŪ�9��]J��S#�c��ƭ'��weI�-~Z��M
�E�)���椦@�jt�ڏ��<M`dZ��$j0���6M۩$��Ve��w�d�*Y�Z�(�$fZq��.���j�9\k'_uvv�"��P�@_C/�bJ�<�ً\���8\��A`�����SKA�@k"S���[΀�(�fUo)�X�	wI�ᱏ�,���%�l�%��x����r����2}(�t��c�=�lcxR���`m�vf��X���|m<��Z{�@�3���L��X=SP|�e%#Z��"U�@;�����av�q�ķq��aV��-�N9�((�N�:�VV<b.�\H1�+�+iU�^m����'@��,�ӹ�p��I����:;f��Us:-����%��jS
��`{F)h��Y�f�L��5,*�Ґ�)�u��H�3���(B�D=�5���lV7�n��HN��ˏ,7���X�ޫ�P�W�������O3�e��ɶ6��x�i�K]vН'»�Ϩ���9�;�N�&OM[\��*�6��7+�c��`�4%��ǖ�D�ɽ��F��b��vd��Ŵ��(i���n�oD�~�o eε6���G��uoCH��c� �[M�9K����[Ω�_gWq;7��w6�c����oSU8);8-�}'�š`j������0�n��w�hݬ�+P(�W�Ҧ;<ݯC�-�wRR���0�p��E�dy]�>��Cz���.�7�H��V;h챓�l�/5���4��E�c]u�8,�+N����	"�v0���ٺ0,��6oՓE�C�C�#���wz�ЩR��3N	b2�jL;�l��BX[u��RVdw��v�:�S�c_��J��Sg�)_j�R9ܔ	�د	3�cu^qtx�/��y1�x��� ��٢��Z��.�b��$�F��ʎ�D`�q<W���Ed�Nk��e�lCG�������`�::dt�WX�k9����#W�l�"��r5vîpҔ�$;����	qPF��z��v�HN7�Ivǵ�9=�[�Cb���6��u�_L�{�hm:{��lN�0ɛ� ��Y��}�C�U�4�F�w�gN�fU�h�:�x�n�.��))�٨��N�;n�����c�d˾;oRϭ@*}�����o!��y�E�jbj �ok'fs�`?�Ù��mI������q�y���]j�8r���f���Jw��q]$В�T{Y�hfJ]�Ǘ΀�����K�,������������ss�(̚�HL=��Fh�p�m�KV+�1�,;�j;k��a�D5�Xܘ��g%J͡:,�',��R���G���{�]4W�ٵ
4!{�P@�d��U�n�8ƃ�-ׯ��Yθ)�u]�׃I��KQ�N&�y(�/�D�D9N����<୧�:PMwp��Y���@�üi�`nV��'eNh�{�V���8�d��w˲����$㕢��V]CmQ��ܷ��rZ�᭾!��:t�̝�Vbմ�: `��̻{0��`6���wjG[�r�\/6R�X���f����E�A��d�E�K�YQ����6�����n󡣮�v�t�T>��I �oE)�#J����K��j�A_j��ٰ�al�[+�^��:��o�|B��x<�˕���Z�Wά_S��x�k�-Ԏ�VNL�K�SVwK�-p�*�������Uܭ��V��k�W+��F�9V��ӏ�gJ�/&76��K��f��V��m:�U�%�ۻ�����}z�*b�*N-�[�AJ����RnKM
r�
��^�8�Ӗ�f����G�J�Y	�^�ҹ�9�*��"A��-N��`}𒻠ܬב��BbEֿ��m-&��hY��ӴU���ͺXͫ7zEl��+_FG'TP�Ԕ���YD.�n*RT��%!n��>F��Njؕ���RnN�T��(��S6�摦�JQʐF&v�C�eͺU���b�$LN�k�	.��⍮�T(fVU�WU��/f����N��&�f������+GB�.�Cm����%,՜�v�\ܨK_}��TX�=(c�X-�;m�qhv+)����(]��:��死�,�?5�^Y*ɰ���"�i�#V�ҫ��׏�;.��Ҏ�E.oe!��e��5��ݚyw.Jv�S��n݈�<�9�[��W;ܺ���4F-N�h�x"��9�1����/xAf�8i�ƴ�Z:���/j6�JCog�H��81P�$�f��-���B5�Y�	��֮������ڱ:�4$S&��i�.���F�Q��n��T�|,V�L�؄��Q��}�����`�T��4�^歗�ùлc��c���I���\����.�Yɂ�6��!l�����5��1�0�G%�B��.�{+��8�t	�6��ë�\u8���1�/!��lV�;�s�n][Y
h�tu�r��]�>�Y]/��
���Ȓ�=2�\�p��i�cz��QH�ڽ�p!9����9�o/f�;���݈o��M܂���,�������*�U�������Tϥj��}��ʠW��|�>�;e���Uë�1����u-�Fm�kC���2U�}����m2;�,IQ>�Jق^��J���Q�o���Z��ŝ��Mо�"�Y�47�aZ�|�����d����ʶ�Y/{UI�����h涬����(��&^�r�_e�&:��-���v�r����8\�\��-���m>�a׌�T�&m�U�2�ᥭ
�6�L�-ӥ�K�gd�J�;KsH���t
ǟ���h�Eh�Ba�[7�f*���P��S�5�sV��/.�\\�̺aQ���vl<"�$"���V�2��zƊb��c]n���m�G���k��X�W��T�Kc)���(����Tw�d�	%�£��=Y���x;5n4��R�AN���Q�<P���߯��e��v͒X���9��C�s{�E[�	Օu!�%���ܠ����.r�@�ޖ�F�n2E1G�s��J#��Z�U�Vvfê��[���.l�V��/�Ć�6>3�8��p�K7'ה��.އ�R@]<g2�V-
2a�T��C�]�[���յw����LY.���Y�)�s;�҆��PJI�����Bi�W�9�&M�X�aP�Y1�XM�YI��k���crd(E�5��A%ٳS&�x4tE�ܢ�&1��7j�]��ǘ��jTE�yB�
�"�7N#G)ʚyC�ftei�0޻ݩH�A�&nZX��{)�8�H�į������Fj�\֊K2��z��8m�ڲ� ����c���wkX�!�hus�<�^�nG�]e�FIr�Սm��nWL�g�S��.�.^��w����K46��Peu`��f�-�YF��1:F����������(�,%`�b�k1J)�
ķ,j���	U�#��=x1c�i>}Ժ��˸{^��IG
�$;���Ց��K�:��ˡ20��j�8��`�o��fB�޹d/�v
�9����HLU��(C;�&��,Ӿ�y���w-��E�>V��$�W'P�nѐ�&�w{]��ҫ�*�櫯����ͭ�b���D���ZuAw/6[���+kKu�c��F/9J׵̧*��9|��X��K���f�Ô)d��-��+'[��|!Aܹ3�b���d����gR��Kz ވA����Pme �,��@9ִ�mh��\��6����^]wSG�R4j��ҭ�t���{H�L�D�[l�$�ABn���E:�H�o��^-���'	�h����R��۵N�4�]�J���SV�:$B�3T��C���+>�ZCN��0^��!��u ��]��en�-u�'U�gwfUn�%н����CE�'Me�4��3�Z�{��ԩ�;���j�:U0G����!N�p��WA�A��s���9Y7ue��,�ز��2I�:�]�c	E+V��F��h�ɽ2������C7{p�=MR|�M��XѬU�GjT+m����:��ie�ٮ� FJԢ�N+u����}+7�������MӸ�Nٳg �wU�h(А7��D.���͒� ��vT8�S�)Y�`0L���9��i�f�rJ\�8Q�]����3v���	0F���q>��)jܸsGr+�:k�r��h�`�)l�w��q�v���G��3̌��i�4��!Za}��u��a�ԁ�"��V����Z���������G�Ć�qN��!���-�N��=у	y� ^ݻT$N���u�M�Xp"�Iy�t��QX�í���ٲ(�adt��W��N�%rF�t潜�i�Jr�δ[+���'�q���Т����y��~�[J�=�}y���X����΅�Iڦ����H]ɼǙ\,Q��u]������Q�eT�Ygq��ChWB�^e�K�\" �M�Y�8�ɸH�Q�ڍ���0'@�`}Sv�hS�
׈.��+}��u�Cflt��J�(Ss����X,#V���G�����а�A$�i�3@��ϖ��C�)�\m�S�����|-2�B:nhS�w]Ǳ�p�J��:��M�Υ!��#$mF�+.��
ee^#�J��F�c٬w �f~rMS��]�.I�:7���'
W�r1�n�{ZS��$�%,o@C�l���^�EX�����;X�L豷�1��y��P�u.p.IL�:��׽ǲ�[u�n�:��$T�(�ޅ��i�oK�)>���&#G�a�MΙx>��6�m
�֡CAT�����'���ٌH���Ð�bM�GQz�u��2�,�K��s����]lnբƂ�Sm��Zn��3��˳	&�'(f��i�q�CsC�R�"lɼ�gU�)Ү�X޲6T�b��Xk1�E�A��rC+]�<���CU��j�vNl�aD��j�Z-�*�{u�f<s������ܪ��X?
��(�LD��Kkznsj���gb��ieM(�J�c�x�j�����2��=c���t
��'nj��Qs��c�Y���v��q<��+*�h*bD��&��ɪl�M� z�'W@_�Ns�D]�]�f�T���C�4��+VrU	�|୹|j.ic� ��w@XpVnhK�TӼ1Ǜ��ɖ�$9���Z��p�߯�&����d��:�7�N�K��Gjef�.L�-��,��.���q���v���c���" ���Ձ�L*�ǽ��O8�� ���9�4:Q���Q���`�PrY�T�Wu0���G��u�4�86��n� �Q�	�ƘN�ݺ|#I��I�����ӵ���7�g]e�Y����s��l���`�Qݔ8��G�ȃ��8�F���wnmv٣R�(�����ٮ���b$z��"�Ơ���hhVRT��z�.%�[����v���x$����d�9S�M�:5�&���*�K�+lݸ�c�N3�uw���6��Ku�����i�|�̥��YܩQ���Z�e����qs�h�����& ӆ�%��.�Z�@ ��qK
�>5��qv�7[�L�]M��ۮ�TP*4I���'c�5δ�%Z� w�ْ��ڜ&cL1]q;%��
T�XV�}&[+;��ܤ���� ��	Q��3S �ϊW8� ն��;7�F`j�S��w޴�"u�M�O�̶;�f�)��hB��|�\H;J�VC��Y�]�C]�u�3���bX���1��kB#ќ�u��`գ��u�Vc�J�ב�*�C{��k��9�ƘB�<�>4��Ϝe�}du��3�$4L5�X����̟�ʉ��y��2� u�#K�{������pdl[�\�8�t����2Y�
�(�:t�D�6XM�;��tEA�p��7�j����qجu1\�3��S���wv�E�u0uLSS�1��%�������;�LX��Z~���H���m�����.��~|��E򼭧�ťK���ρ�N�_@8���9K��"�E�8��
Z�U��}bX���wlZ�65�]��e��m�(�֍Xj��	(>[B��%��Kq:5��#��fKm�3#���<�%�A�*�	�t�l�GVԉ.&�J\ǉ�u�҉�����#�9��Q:2	1vGԬ�AC�٦P=�#(A��ͫ������od�6�B܁f1��[��K��p/�b�;nr��v�p�;t��,Y��b(��ø���] ���7�_u�85�`�,���0P켢�+t�*x���9��� ��q��u���I��`�ժ�p!�	]2���]%��b0�]�����T6,���$�jC���_X�&����/z���0&��w੏�6��ӮV�M��U'm�A�=��ҋ��q��VR��x�QŖ�m�q�qe#ݚC��@뒔���&ڨ�8E=
(p^��k�	��л��Z�vf�Cru�j�|ޭ�r�|����ٯ-I�U����[��#�si���n����!����c�r�f�B��)׸:'yZ^۠*}�-N�Uټ;e�v.�ft�����nΝ�Z�5eQq�U`Q<�0;�ぞ�k��-v���=�!�U�Y�i4;P��Jm)W/�t��Ԯ���`��n	�0�zU����y�X]��k�����Qv���4�j�@�Y�v��f�:����\��L��ng�PN�j��٠JJIl���ԡ�:�`��	a=wD���ܷX
�negq#�m,;�JG)��v�c�-��_/\��_�������<x�o����f6ͷ�e�/������>�����~'�~�~'����fe���yp��ݺ|�=�'�NŁ���X��[Y�j��wGwV�]�oji���p�SI�ڮ���yCa�Fa�ʯqG�	c�)*��>sa�)^Wu6V����4��iG�>XmXh�t(�A�XI���h��Lsk��yb��F֟����"y��D+x�V���X+SR�ַQ�3-M��tB(Y��_7Fg����ٗ ���N�SB���MV����;�f�]�d���ڭ��n7��.t�L<P��ܫ0f��-�;���'fauo%�I^IQ?�R[\�`�rg�X��%�ozL粦(��I)F���lv���,T�N;�5�o7�AY(�Nlhԩ��Ƕ'A,�(Vx�ӆ�M4�У&���ط 2p/X��;S�YƆuKF����=��5��*ipf�I{�:�U��m���(�j�_�M��,+�r�����S��k�T���+��S��`6�������@����H
�F����1@l����t��,nK���+�)n'��:��Oa��J�h��u�Z�\�:D�%���䭙ă�50h��D0]B�f�4����ީ���5վ�z��毻�i2�^R\�A��E��(�	����
����*t�Z�.r��e��i.�����V�.;z�VE��o:���Lgdv!\�H0�t��j�E�x-Y�����*2�� � �������je���ٷ-Y*�&|G*�R�M[SV�(+g��Vejǉ�l>&g��)��[ea[���ղ[y�f���Yʙ�)�^y����P�����V++!Y����Q��V���-�-�'%l�ܷ-��Վ��Sn]�o��۹�����\���55
�55og&+j�Z�P+e3u�j۫���m���ۧ���8�8s��k3p��R�jV�K%`�aS@-�Z����6��*y�=�:�e���<H�hҢ�������'��Ϝ��P=�����Fv}p��V��ы���CWQ8Ó�ۇѻT�z��[�^�a�yG�/u����C} ^Y�<sΖj���1f4�e��}Ci����v֑�=�\lˎ5�c���>��˞E���7lH��t��.uyVj�2��E�<�׻=�E���2r���`��C_u�W�pr�X{K�۝E�v~ޞ�]�Q^Sf��Ǿ^AΠ,d^�O���}�=�w�9VtOZ��c�0��2�4e��q7C���Z���<>���y��ku�.���(*�<�&��#;q=4=��}2gϘ}&矍���^O�ֱ��I&���6Q;1A�o9Pϩ�6iŜ��r����;�,��M��_���{�9:�1���`򫽗�~p�ŋݦ����84��ڻ��}�������O���Y�'�Hr=��
�.��q^e�E/N�m]�м++I�0(�%���1�[nh5�]�q
r�k�`'��Q���e<��5�R���f�\p��[��f�ͼcʗ��t��庇���	V���SY�WkX�v������>���AS�mz�}-���c~Xz�y���uZ5��[t��K�-ɡ{!Ϥ5p���HU�e��{��������ۗ���k�u��V����}.y�z���ʃ��&٨h{������iW�`�kfټ�=+N�4Mӛ��^u�@c�F�T������C2M�{/�+��I{�3�����lz���ޤ����Sr�{�枯=��~T�m�=���M��'�L�x�踽��O�������d���+��{��Ӈ����K{��gվd����2W���_����麽���'c�9s�&	��7�2����>�-�Y倭�en���~�+��{>=�����P�ꐛe��k�~�:I�{�x�����wT	�y�cR�3����LȈ3��Y�3Ր��RQx�OW���Gc�l����{Y�w#�s�m�[�36�!�M�G8��v���/�s��$�͎a���h�{x�i��$�][��oD��)Z�9:���"��x�tz�=�Vi�t}(m�e�ǎT;��W[L+�R�ʘ�J�Z��d��4t�:�S��.=�����8:Q,"oV�ް�-M�7a���D��*��zK�{\Ƶ{��_g##a��W�R-�+y��I�Ǐ2s,wj�i�n��~U���y��7�A���w]/V���Z���#��Nh��f���Ĵ�w�Dq�����I9�z�B`^��B�P��5�Γ��±5�rGF���2��W���~���K�*9Dv����%����-�;���۱�"���~�D>>��W�c]+���P�[����*�%��?uJ���5�� �K@�'2�=]G;bD��c#�����O�՞��{�S_o��+���|ל�~�=�Lv5x���2h6��l�m�]��6�os�/�4�>jg��3 �H��hRs��[�/jn�}=�9�Nn�*�����U�:`�����+*qk��F7?]��3x{�WQ���P��4D1w�%�nZ����9�����iΞx��+u{tˏm��"����V<�T�����mMt�f�]�y:ٱ�_=,<�"2��ؙ��ͳ�".H�ͼ[�=���z&=}��J�FN��2���]����}Z��܂VZ��3��nB.e���w]��¢]��m�D֞^)%�kꀶ�Q�פd��Rvݣ�M;��_5P=�g�]G*��sԂRR���7�>��|'vd�����'(i��T2-�<z��Z�uh��ޙ�WTL�mvz����}��Cq��滸��I�'v������xm�b�F7��	
��\���V�{��T��X-���V�o{�	�Nox�d��^VsG]�`{}r֏/_k	ߊl��А{�J\ϯ��
��=\�I�`��f�sq���ru����ݏ90�>.�������Y�o����Rv���7���̳��,��gO^����e��d^y��}��y���CwG��EX��㧮=3��>;F���t�iƖ�����k�~Ċ�ŝ/�K�cI�T����cƽ���<���j|�J~�]s�6�'z�����2:d鈫��f�}�����z���c���\�v�ºY��e��[.2�V��>�i5c�mA#c1�ËT�
b���n�i+T�	�r�t�N�r���=�Y�1�T+(�Z�m�Ϭ�6HN���-��j5��u�Gx$�'W���}�(�1<�K/�7�;�L�RZ�bo!0_#c�|^N�~���|L�gٟ�W�Z�җH��г�c��E��"V|�w!����DU3V�){>�\�+A^]�z�z�9֪
7�0x׺l+V	Q8)�=<��u����p���3����WyVc̫ݦ�v��~����&훌Y֐L����a���C_C�������2�������z{d�2t��;d/t��:�a�|�x�Ď��=�o$�ot��p�T~+~����NU=�V�s̒yDȻ�~�n͏6�+"x8�1ڐ�-S�f�n����h��s0�ޏ��7O�J�^��9w�q��[�T���Q�������{٢�;ҽ��\�d����Ȁ�'�Ϩ�}ӑ����zϏ�,�M�?g���(P����a����۲��7o[�ު��^Q2so��ȯN��l�v�W�m{O��lX�oNK��Kg!)���;��'VC�	~���ٸc5�{GG1Q������i�^�� 	��K��h�.(��`��-��-�;��B�U��� dv {�rc�ی�58��xe�� �E�<A��+��B�Tr� ��mL1G�cVw��W����6���U�ƼӞ�?eJUl��3����!������.w�W��//��}&<�F����lמ�c���~=�ؖ�K����qjZ%z�ס�K*����}�^����3�;�/�/���M���%z�ͽr�=�0?z��U�hC�ُ����o�Ͼ��y�O�A�=��vM�(�̳JVߌ�̡�R�p/��֫����������	eJ�ݻ����� n�����a�L���R���Ӫ����� �޶2�s��~�G��X}"=^n��_��H'�HsDt��׬.�s���N�+qWEt6u
�70����u19>�B}��H~�3��zZ�sWj�k�H�g����
[�)�S�U�z�ǻ���z��p�^�@z=����䨥+�2ߪ�ߥ��|o\����˹�����	����v5�6���v[�+)��]��6�M��6�Y�$B�Z5\��E�z��).K
�X=/��ZE�x��MHK��ͩQŽ�^S��!cT��qr4*�#��Rh@ ]!c$۳�Я�� �9}v�ݛ�V�\s�1vG����cԧol������Nd���]�f_�޸���߱���Ɲ��� �D��3�>�;�v�<���iy������W;�x��3hm����]s�M��B�Na<�z_�,���L�g{ۦW���c��Uj�����ݣ7��.�c�RS�A8�{��>N/k?{�sx��W�^����]�������V�����׼�=�z��`���7�~K�>�׶b:����kֵ��s�!�����V�^f�}��|�	�i���VӉNM���q���$o�o�����/�x��������K8���y��{��{��N����,G�fP�{W���^�����JWa~)/X��.RM�o����>����}YG���;7=��	���ݍ�M�͓�f�ϽF�������>�:L�=�m�e�d��s4��Ǭ52�-�)��
��#YZUȥN>�O��>W�vā�R����q���z�2��'[.ʣ��6녡W��[ANu1Br���m[��������TS�Nɤ�J��5�e�K�n�L�Z�+zpO�vIb#�G�.JL8ټ=G{uM�(la��gu����f�*s=��5��\���>?\ڹ�8W��\�D|!P����P��RyWWLib})�͖\���{����v���>M��tL��0?U��5Q}uY`��{�R�H��3xuu>9�����k(�z���=��7�]�CU�ӝ�<Mj���y�d�K��,@����t��	߾���)?�׈/v]�� �Y��L�ʃ�/\*a��t��@�=u|G<�rr������;��b�)�7���V�\�۝ʠ��8��ᡱt;��9'h��o+�S������+ތߝ��!����L˾4�f	�;�c�����Iޯ����&㏒��Ov����$r�]��z��y򕲳=��i^��5�1��5���G��g�O�Q������6�� u�ϲSg��eS�������*�NF�V44T:��ݺ�� ����𹠰�^���U��w;���fd�1�������0���b}b���X֚8	0ѩN�Pތv�̮���9L�3�c��驥��*���Y����f�Q�rvm�Z��n74�?]v�����"���^>�������9��g��d����N;�Yf���;s�{w�x1�j{7y������WW��K���������S[��8\Fj=���&�Ξ��y���厽�|k��mO(k����ˍ�����~Kr����״.$~̎i[�ΒO5^����{�3��TLn���ݴ�t��hƲ��HU�]/]"�i�y�dO�������F��bnK�8�I�z#fn[h7H����]yvּ�K�o)�K����[��#4�;G5_9�P�4d7Pb~yj�_A�Y�:xw�4i��O��������;&�}��p$Vi8ȯ�:-y|1e�<';^>�o;������te�����&hqH�;N��h������=Q{˒�=��O�������eMmx��;1&�'����lB��9���ѹz|�ߧPc�h�u�0�i�i��D�H�U`�@�v��d���m���J��}����~�U���Sa:Rg4ҡ5-��[��|��H�c��j]3���P���@N.��6v���#!g�yώ�\�åt[��Ω�0wP����n`��w�	�F_wȈ�Q�5���k>�����A�Z��h}�&�q�nx��*��J�-O&-�^)��L|�ܯ����3�d���B�7|��6�+������N{�{ '?G7�ʩ��}���ݾ�V�U	�Ƴ�g�~/���;��Ŝ��S}9��#�����׽����;��9V6�=�.@R�pMH&�������W����x9���ܬ;��I�������ҠDݭ�vd��{�}��'z������y�ߛ��6k������)P/\�:�~}����fR���]��$��w����O%���R�æӓ}Cgl��_����9g«kA��K<N:Ś�}��/=ez܃eח��7��;j�����ĉ��rA�M�;����<�zD��9ϼ@rH�mpsCY�����3�^a�_��횜�9Hj�F�:2?��/����
��, ����E�N��j�G}YrG�ղ�z%�5�s'vk=nBѭ���]WK
m��Los�I�;��M����cL��E�+)kaִV��N�
w��^�7+FEu����*HU��Z�;[\�)�g��:۵rd��+�6 U;��B%����u}ٳ,<q3.����5VQ���P���J�T�ݝ	d�H�t�oj��ԟSZ.�k,����l�)�:��Y��e=hI�Ӄ��r]*ůHx�ܪo��Ą�4�l���"�t6�<�����a��1$5&f�*�D6�Æ1YYWe��F��.+�7�:���+vhH:��.���s�9�&h���"n���]M�D,�d��v\ @��3�o��D�zga�
\�G6�.X��m��i�٘B�6�HhI��wYD3�&�c^���N�1�����P9�����nP�?vPϯ���s� )���J>�ko�Pp&���pT�h�>������2��E���=�b6CN�͜C{�X����攈���fK)��]��*Hm��ǳ�Yl��3o����hPH{�WuH��K�ͽ�j����N��	N�D3z��	��%ƺmry���]Ad�"7A&b��.�1�
pmAL:WSt�vO�̬|���)�
9��B�3�5 :z�f� �'Qʎ��ΰ�l�d�r�+�=�2�m�sJ�_̛>(��x�vX�P�[��x7"�3���C�����t�w�pĬh��5�t[N����}L���^o8���$����5r��ZK���X;�e5�F^���\���ٜyb����W�P$����6�e�8�a�ٰ��,�C0ֻBS<�X3��R�e[��S�4�hɓw&oX�2e<}VH�]]i��}=Z���2��@���9:��d�o'��W/��VT�u� SD��l�Q��\�V�hŕ��դ�\��z�2����4]��:YC6�=��c�k	l�wՋ9]�e��˨�l7��Lk4!`��E邉\�=�{3�qL�<xj{]��.�p�����5��Z�ȝB2m�RU*e����K��["������6�V�:;z��+�h���i֓;U2j@�#�ޕ7�=T�9/U��Ҟ(�8�WK7ة4��h�o$A�?uȪ�C��m��]��V�]ER���]�(,�'K��-]�
���/��%�27��h[�t�c�3�Xf�e�d0�<��:�v+�Lt��T�Q"\�6�T�$���v�*6<�n^R�u��rGa�׻̪ږi"y�cJ����kW��^�7�7y�η�]�bƎ���`겦*�A^�jv;�"D6!����k3�= �:<(]nv�b�Ǫ<�Fִ�j@�\����%d�5v�3��Su��e�������1p�/1e7�a��u۲+�H������K�%vJ��S%)�R��~�޽��p�������6P�*�Sm��r�y�
�ej�MY[+VՒV���,�f�wm�5lVw6��.��Fۖ�M��6��
�w6;���CS3��iz�Y��Y�fr��7���6�++a�f�Fj��x��۩���7�6����u6�:Y�ƛ���G��[��y�J^������ �P�SJq�ri`�[.��7���t��O��*kr�Ry��a6��7�C���~��\�F��F4��2���ADa�"��>PM�/���@��\^1{�5RLK��ih݂�z\g�1��������������y0����נ�:ẉ�k"=��f휻�?�5���.$�?�`�#�?�@��c��^��٘l��v���Pm��e�[A���M�_�({�;�/��:�����w�S�HF�:Qw����f��D�mC�ӷ�z"�촚�ֹY��is7:쉷�od��?�CdD�|/���/�E��LL�@���mmo=!�Ԍ�׷�k5�;�_��>�W��dݞ[2�Ee��a�[�]��lnG�j>�����}�|T�w����O���Ǿ��T2�GyP�k�cR��"�Pnn�ZS��כ�ʫ��s+*ƴO��ֺ���e�]��]�9��O0�?}(��]��r�x�{]ψßoznP��Y}�m�{���U���?&�Y^�'��;M�%t�\"��E'��U{���$ͭ����+��m��F^��*�ʇ��^ш�*���韼��#=�Q����T��ܢ�{��芢Eʗ�=y;��}�/{8$H�%MdQj]8B�-[V��
��_�����ǋ��A��ɂ&!���ڼ�P�����8�i��L��3���[K5��qi:��)���;O:�K��n��\kL57]R�y�t��(��]�QD�-ވ.�]0g<F]�V��owν7�ra6|>��--,�)x�#L��6GP���K[�5X����|2,�\��[T�>�])=g�%�۲��=||��%/W���`��0����n���V��<����r�lY���������:~�|��c�:zfϮk��p�`�΢4�K _�j�o�w�Ϝ�Rի��z�u���c������Vl_�B;�@�G��ƖuU�U\����ȃ�]�y�\�^��ݾ'A�H���BBv�\}m���|�y�y���� ���%8�E�ڪgWu�^	������┟R�q��!V��?W�Y��nϴ����%���ȸ6]�in�ŉ���>|�A�nu��r���t2������:����}
Xz�YP;�n٨I�h�ٱG��|"~��>�3�:���ǉ���Ԋ}���ŭ^���k%U���\��-�F��|}z�x��>_L�1�eNBty@�8�r�\E��8|��*�t����9ߤznj���n��x���냏Y�7aƹ���q�9_l�+lr�aMC5L;�lv�Tj���G���׍ܕL*s&a|pu�ub\��U�+��ޮ�=<%��0jkZ)�gc�1P�#aP���X��4�A"ج�T��\&�1@Ľ���[Z,�fn���1���C�m��,]ێ��._-B���og���7�!��<<(2��ޕ�9��h�ϊx���d���Ԋ��;�S\pߋ�E�dQ}�wh^�U���\Z�vgY��w7w;
�ytE8!���wB����)���q.~۬<n6z���!�s���괔Ή��U�y΢�2�^P�9y刜� ��.s�jD����p7��	�p�@���쒝�(���l�%Wf>��)��`%/�WC�S}l3�e���\^�<��]P�^���*u�؟k'/�0��u2+�u,�V�K/��Ӵ9˴)�iIH�ѓ�UY�&wǰ_J�*U\yLBu��7+Z��/��2e�zͪ�2Y1�9l=��P��*>HY<�C��B�����춧�_��	���39�Q�����*����[�;[�{G9�B�z}+V�tV�z1�RDW>۸=U_&D�qDP�&uH���^Y_N�oQ%u�Ĥ����Kd������p����;�q����1l���!@8��!I�dL��C�E���ӭ5��LQre�H�[���~ �n�s�;���ϛ^���Һ�?:#��G�T�E��~�֑B²�������C|T��_}[Z�MLӺ�kg�/֚��L>8��g
�����Т���M�5�z�h�b\}C;1tr�|2�����M���w����uٔ�u�5Tvp��xP+I=�v�@.l�3�9�u;���v��z�P�Wl��:��y�3�}},����Z����\����ڜ�⸏s�d�AI�Z侽��H����X�q��V�ۦ!t�b�P�[
�͆������b������=�}uB"[B��z\.����"u=�,���5r,n��6	5M@�&R�s�P�$O�=����"*��FLԘ�Vi����Gq��N�+�x��._�Zk �ώ�˪6sX�bC�=\�c�!@3,��s*�ֽ��}�l��aI}���B��+2���|j�+��VMx��U�c��O�}�����,ʍ�����r����Y��U�YQ"�ƨWjBT]�Sh����[�|ɿNLzt�E�y��7a�X􎸌9m��\���u�)(̈��uq^}�i��l��MW��+d���,�kj�|2�2��F��wQ/~1�0Ja6o%Vv���[��>J�r3&#ġ�=�}/(����I��3m1����P����q~4����(�5�Q���c�)pE��y��&���ty~���� A/8�@���m�����E��Zד����]�������K���3�*+�u���a�Y������j�j�a���G��W�P�r�c�n�gf92�ۃ����	^�W�����F�m�t�K�r\xq�߯�of�X�,�.d�O�Ύ��t��ͮھ\X������JX��sP�v�'r������U��5�ө�['��ُ/��RPr	)�BTiD3��9#3�ٱ�Κp18�3*��S���az���t:���^���<���	ޕ��!��ʝLЕ',��������4m���ϤV�?H9�KNXS�i�5X�x\�ux��2"� ��B�r*�u_&8�5���{�];��"{7����!�kW���Z��=�T���1�~�)qѡ]1�k�̚��ӣ����l��=wHPK�P��q�Y�t�/W��䩾���7V�Y�o*l�1P����#׹�m���_	UX���;���M�P��fs�G���(Xn|�OpDP�SQ��y�O�qRד�)3)A�{�k����9a����z����	R��T��Z�RrpB����o��7��#{�!H�oՑxǪ"�:ۦJ�5����m���"m�o��5�5#HMWM�MQ�f��-f���i�o+�,m�"�z"$j�{/B1�9R.�"�e��S��:�G�Npw9Yf��a���|�,��y��9��+��V�q)x���h��p��8|����Z�\'
���� I�9����S�w�.9����>w�R
>��t��gua��y*�G���f_w/�=��:ma�X��0��AZ�t�;��1B�vw��q0�-��,h� ��<�N95�|KT��@�|�'i�w���W�o{����"*����ۗv���o:GltIǲs�o�R�5E'7�E6�oXS�!Wא�=t����dϳ�Bx'���贤ZRܣ��;�F��_!�t��%��T/�ecg�m�d��b��ި�t(��LfG��B�<�1�r-d��& �ڂ��s�W@|�-]ϭ��G�:�7/ �
�������Dp�+l�C�T=U+��#�9�P���09�l�(��TMؙz�߳#nk�Oe[(�r(lś��~���QԐ8F�a���5��>3$���KX���Y�Y�3��@"���Z�M�#%���+g�{��t�O�|�i	��k��;��oc�X�{M�i����]u�����U�0����6�Q׽o�x���F�' �$��_K}5{�Fc�9)��ZjPw�B�'�ƇYs8�jFE���u	U\��x�~�ɩ\=��\�o����,����w$g�ܳ �]���E����Lk��۽)��kK����tDu���ndF��a?	Z�r���#�#q��P1[�lc=�^��g]��H[������ ��l�����K�vØ ��K.��'��d�H�κ
�;�G���*�Ԅz���:�.��g.~6�����<�V�}�j�����[�tu�K�z�0\x�i��^�*U�ټ�M"�Bm�'��j���ҩ�NG���ƨ��-02��:w)�z����� y���<��t��hn-��eρ���h.��R�qB1y_H�q�$X��j���g淥���� 7%��u�h�wN�Cڸ�R�yԢ�O��r�7��z]����:g-�����-��u*\٭ ��qm�j������`�n9���n�
��+]Q�P���b�3��5B�BЈݸ%���b��|��L	�O'�s����I�w1�q����k�ٕ���1�$����)W.k]N�Pώ�e���lR~��B��TĖ�}rL!%��b��A�{h���Y�\����1T�m�A��J��fP���l�*i�])�d� ����W1�9m>����lJ��?G9V�W����v�#웫,���1�&.x��'������츢�n��4���1w���oO�"2�K��ϰ�����t���n�v�z�K���a�i��0���:�)�s�7W����"8��u<,���B�v+
{����_�U�S2ס�)粔P��&O�ڭaa�uq}�4�w
��Cv+��S���Ŝ}��n����8[���n���un���(ꟑǪ�[����=7Ś��������9�TO���_˘����P�o{�=��t�{[�OM�4�MƂ�����V9ϲt&���y�������)�hJ�q`�b���A��þބ��G����꯲�ù��Y����\����׿~�|Z�7�X����"��G� ��80�P��Y�	�?s��T�q��gJXؼ�z�Y���M�K�u� �C3'�{1�͊�e=9�[��|��dbg#Ϣg
��q�v��vM��>1q�'Ώ��@���)F��D�X}���>�>���5�'���.m�Z�n���jS� �{����,U<h.�z�9�@�q�"���*�XF��%J�;F����������N��[�,丶bU�jnY�W�l�D9����`Eభ�S똌������js{8ױB.�z}�����z�
�|A��⚭�X�3��T_�)��?U�^ο����.h��T����:Ws�E�b�2��C7��$NP����w��]��n�oGn*!�s�ډ1���ͼ�K�jyn��2��u	-5�m5�x����A�QÖ�:ȿ=��]�__��B�5Q�#f@K��~Z�Ƅ!��i�[�ɯ�wJ�g��j;V���KFl�/��7?wD��v����,]�YQ
G���RWj�E�����g_�)�@���$����1�,.�/X� �V��?�g���S�u��F/������=-�)����_�ei�Ru�t�uV#��Vo8b������c��.x9-[���v ܢT�k%�Y�ˢ�]ʚ��5[Hs�����}����}�����jٍ���f��N�l���;G���Hw�by�x%2�jS,���U�o�s�'�E�@�/!��;�G�ܻa2�zg���a�[vxLB�ЃNwHy�q�^�"S���uK����pb.�j�)��R/����Kc�s�}�����l���:;�y�4��sJ�|�Se��?6�*N>���Y��۔���|�7��x~��":�W�!>�zT6�W�%���W-�NЊUr{u��Df\U�:j�~�������*�r���u9>/P�/�7�"oX2�>�TZ��S,�<d^@������t� �n;�->Z�.r�9��`1�[�kyA�L蛊8[�T�m0���mewC;���l������U��5H�U�D��c^0�������ȿ��(�:N܃�ޢ�'�;�t^�ϣ�F��L�|&=��l��"L���RR�CB8�b	��od�|r����s5�z�8!���t^�����C��.����qR����p{�smR��Q��q?<�ϳ�n���/�����C��'�w<`��-}?ng�3�}D�=��(0�v�m�-`��F�g3�*����n�q�l`y1SS�$^��Cc�ͳ���u��M�=y��$�c�H{v�-/nZ���;5oa@���|��w�Ip�P����Q�"�ӆZU,	Okf�iNM��e���j-Au(pc_>�y���?7�7���_?Y�o�V�o�ٹjlefmX5`�A��X�6�ql�ڶ�ۋ�U5e+-i��_n�E�-���_��C�j�JXe(7$����k�V͟pu�v����І�4�)��7�4�{��9}�C�i��C9��/ޤ�T�2�b���Q���U[_s�W{���6��Oԟ#+��.��-�ny�3���VM��.�5E�F�G��Hݫ�s�ꋑE����$��k/fP�m���gK�FTwM,r�1bıea-�m����Ʃ�xi��e�.�oy��[zi�A�:2Q��%D*wk���n�l,���K�t��Q�N��[R��J�[e�,�������m����6��4{��^>�q�9kA��NZz��M�n<��_V�lj�Lz���/f2�#"ш��i��.�����ȑ��1�Z��&>�ιgj�J�[�\��M+�(�3��{(��ƕt���&�.�c�]���b�ݐ�C��UJ�t��φ{T���nY33���{b��C��R��$��n0dś��~`�J�XFO$u*7UJ����m�l�zxB��o�g�.A�"����4�]4�{φ�B��J��)#�3~������ h� p��Iް�5t����g���_
/t��I��N��a_f�A0],�����Imm��O��,TZ��b�"�e���Qv滜�~&��!vJ�K`�3^ƻ�%t�	|�5�ŪR���]x6>yc���9�'c�F#�03s�j�y|%���)�e&�q���tKw���T�س[7t��!��\�rXmh%\U.�ȹ]�Sn��iq�&��?u�S[�4+�%Wl�A���W$�U�/)jn�w Y��ހe�� ;&㚬�љ�f�8%�z��vq%��7��� ?!`�:��d�=��@���R;.�U�X��*�l�X�Z;�F���7��]�x�3d�ըB:i%n�C�+#B�h��C)�����ef8p�4n���HDfޮ9���M���=\ m�sp�(}��t�-ߴ����7�����H>N����G٭����M��s�Os-��&�%�8����[�h&r����w���Gٻ��l>� 83 x�
���=�m�-]���Aծ�s�����P�*�bu����mE�d���A��ѽv����2+1fY]]�u�r��*>]����\A�jv��C�9ޠC=�]C�бa%Qsp����oF�S���C0e	-�7�ѝAi�{RlDB%Ztaι����V>�M�!Ы3wv��MͰ�.�B�m�᫔Tåt��:�ch^�
��R�5����d\UBn�n-�Mκ�G�j�'0=xX�x�i�QN��Pc�����0L��\u�ۙ�������@��WQO�}}z���sL��C�]��=�]N��p�F7�ҧB�:��b� 
L�ޝz��ދ��1�.s���,�k^�P��K���,qlSQ.8���`Y�uP����J�l��[�/W`ʕ�EeXY�%䭝C��/xQ)�P.��������˕��[v�s�e\j���{M�mM1�S��-�g���`nB��i�Nхa�Mq�T<�'Ͳ^��"/kK�M�4�S[�]>��S�j��a������D��w3/��c���Yw�gM�j��0�����*���5�㲷�`W�r]d=�r��G�����5HZ}a*S�^�l��@V�}9J *�7�w�rɲ\��yc��7Cw)u�Ϭ��5�S�!g�ʈM��v�̛�OJ�#|ԙ�v[��]vT��Ԯ��KT��Qr��T%��wؤ�9b�
�̇��$��p��5��+&"�q�[TƋ v}�z]��:�GN�s�;	W3�-��3#���G7�1`�w�`[,�]̎�
y�ɒΝw�����Tic��J�ۥkz�`ړn��0�a�#����ڵ��5جJ:�h�|3�r��)�w�$NS�q�j
UD�,X�5�k��_-��Rk�S�]�0f�X�4����Q�dh��j�Jʺ.N��BUc8�X|:0r#��ƹR��V����,u.<�i�Z/�kg%F���
�Bh��=�N��Ǜ¦�����]�̱�k�5��X��o�M�܊u���ZT�Äy�F�s�2�#�^���B�+���[�s�rO����ӯ(q��@�!Z_�����M�-���-��άu
�G-��ۖ��m�M�����6նy��o�#w��x���;���Vά97Vǋ:��w`�g�rͺ�ܶܔj٩����ru7R��g&��u�1ݝLrΦo3��e	e7vr��ո�q�gV�W)��]mՔ�LVw:X���,ܶ�t�Jm���s�e+.p{��(�L���91Y�ul���s���ն9g%���oo����3��FVV��ڎ�ι��R�ulܶ�Xr��\�t��c���S7'Sn�s���ϑ�����U���W��oG��+�7�Y��r�̍o���R� ��F�L\*0`�	�� 2Q�i�}��]��u����_<�+�~���Kf3H��x{��8豨��y��/<��ا��dVU&c�:zd6LO5�k+����~��%����Ow�!��N���
�XjP��T���C}˦��	��ZhGP�U�/:6��s�C^�΋|�]�J]5�N�T�x���<��8̧k�돯�^�4:;����ţm�r��;D\+��>��+�E�>��B�Y�)�0�v(|�b2=����;�l�ne}9�/��R\WSvU�����[.=�V�G����,�TSYœ��S��W�'_-���ޞ�:m�e�'�Unl���΁*j�B!� �2q>*���Ԋ��䞯�8�S�@�����f������lnq}'	&�u�^��e�d*�j��2��R��A��ϡ)�Р��k��P����g���S{7l��izPe�*�GV�˨T�]M��FV�A�9�m?+������q��bbHs���Z��q	�B>� ś�V�}!tJUA�4��)���%�~[���V�+ל��^U|z7��z�2W�S}��B�<�"}p�m?G��3f2��.&y�+c���h�~χ��<(t \W�ִ�t��B%K_5��ۀk�V��nU�����T�7���~���̍�iaY]�}���]5B�9��v	��2��"<�X�9t�aFLbf�e�ԙ����0tY@gIw@����P���&
�v"	�.��ϯ������ןW��}�����,m���a��if1�������׿��\���9��ؽz����NC�c�����'��Z��������`��^K=B��:s�a�^[j`�W�QL��
�H�nƙ������z�>�L��ҹ��i;��/�u^��ra��ת���2;����Y}c\�i��4��\N=^�����_�lJ�ý|�ё��E�y�TP���'�U�U�-#%�cC���>�ÌW��x�n�bt�a�c4�,�LG9j&S��l]�J��Up+��Gs�"�k-]��_Z���a����h1�=)���zT
��Σy�f59�
ٶO�[�0�V0 ���FA(��Y�s΍� r9��̶��Er�ȃ�*�oHRr ,>ڹ�IӛP��,ܓhz�}4n�Z,�9z暛�D/���,.���?��Yuʀ���~?y�o^x�v)f������[�ެ�aI�����B��[�(eWt&C~�_���E*��%b���wXg�<$�e���9��)����J/cj\f9��;��r����f�X*)�_��gO���krA��-u��B�Z����jî޾�w-;%���KM���s�wkT6w8�df�(:~y�8�d�Ѷ�G�f�_0$�5���Rnhy�5gAu�y��I�� ���
�ӄ�;�m^��N��%hPV����v�Fo)(��0衵�k���;�Ϟ��e�Y��m�M��A&��f	fm-���7���3��T�L'�?DKl���@� W��Yȿn��u��2��;6K{	�m��H���6c9�v�]����$�TO��F�������
>�05�Ц�~]�x�;�SkX� ���YZ�߂���Qb]�!G�e�|h�Ut;�N ���:G�4!	н�u�>���ݰ�'*5��T�'ү���i����Y�}m�?e7�����D/I�'�X��T�i\�˖�+��般\$rc���Β�|b*e��!t�uz��0��qb�8��h[wy�s����C"x{�>G�����
�k�˒���g6�%x��?�c�.��'�/�ylMv��ډ�(�#�Df�:hK�j�>��o�������sW�q\��i�շ�;C�{FGz]����C�L��sN#�3'֮v��xcc�T7���1B+�Ur~�@�s�0+/s���=�����T9jJ�$���xLC9�S-���E��D<���[�l�+�l�=�.ݖ��⛍:�-�q�����9�ѲyY�L��0��W��F΢��5� ;��J｝j{o/�h�X����1�x��:Yl�C�{�/Шk+׸�� ����mc�>����y�\��2k�y�Y�=�n�2¥���Yi
����ݏ�C���rM{��J��
���n4t��ڪ#�_U}��1-�$lKm�[2[i`�ƓlĶim���d�Lm&f�g_>���\C-\�KC}m~H�-ˠ�Q�_RR7�p���z�:zD@�w�(0��W�LF̫����f�%�U��j~�#Z�GM��L����z��Lק��IKM����}�������B�܎�n<D������Uh�n�hl��_+�u���,'�dW�&��y9���
!�B/)A7 ��D��4%�/ |�ufPF7z���q�wu?-˦�PI�VN�s��[Qf�C�g�G����J��(7���
�oG�?wO��wd�]��B����4LF�e��+\�<e?>�&�j���P'�p(ȋ�OQ�Z6C�d�����jxX�P�n*�~��$�,���,�l��P�qE�'�~2��#�*�v��{���P�>��=��cv�*F��YWC��kX�2jYY�o}�>w6j���Pg�qW�S����ݭ�������j&�>�8�u��ρ1I�>���}�E6�S����O�	��W��M�<+k�^܇n�h��w�-�9_\h/�4�Z���sT���}3�)������x�:�A%Мl�-w�R^���i�k��H֩6�DJҷ$���	�\���Grq�ٓG��&f�B	h J��F��w���mؼ��1s��WP2��Z:�*sU���r�l�9Ý�oёN����+i�Q�٘ۙ4��a��}:��e�i6K%�H3I�)Km�3K2,ě4��,fI�$�z�����߿�����,o�9Ց����]��M��Ș�g��Z���d^�v����ާI��茻y.u.�	�5�c]�Aۺ�#�v����:��UJ�tϔa�%�D�v��.������Q���a˺�\�/��\}���l�o�C�):��A<��%F꼥.Lv�Q��+���iJ�~�R$��fwP���=Y�M�$d�����JWY�9"#j�O��\C]��ݷ��(���%�:/t��#��{�`�I��)�t��g�t	��0���":-�z����b�����+�-p.�ˁha�c}�I���hv�2�Ɵ#"���:��/rk*����QW�`��煒�Xeʇ"�H���R2�� �]�\}}7ڰ;W���� �w3�$G^m�WV{��úK�,�z�(WxB�?nEB���������yrM��4�8�5���N�6�ԭ[���K+��J��>y�Y<���j���(�~W�"aVoxv�WM�_�R�N�?�'3*�\�p��>W�i�!�R*_O�t/g�H�I|.��#��Nf_��9m�3��6�z"�}��O]�E�(&c�t�B/>M%����m���Y:\>�7�y�yu�J�vm��0��/�u9$n�"�\2����
�S*�q��6�SWu�^���˕Zj�m]fg��  �#���0����Y�m�� �W�`��$Wޜ�ǩz��/{h}ܦa��!2�
�k��k�.��y�_����#S���ǟ}�i{�?}@D{e��V"-\�*:�j�m����\/qMg;�7�2�f�O�[�H��?��?o��7�{e���~'��ҩ9�u8w�1,��t2�T
�Sr31��Z��'�B�r�m��k�Փ*�6�G�ѝ�6jSa	��c<��१��Su�BK��uc �d��	O�l{y��g�ed+8��b�܉l´8�+�x�/�3���2Tc!!��a����I�y�S-~���"��f-�3��n�f��Kss��n"�v�vM�~5��`�U�Ȩ[m@W��Ȯ�y�N��ױ:v�˴(1�$���f�B鼝W�w؂��/ܘQv��z��)S� v'�TpїiO0䌖G��u��yL���D(��6�<�x�/�-E@N1�<�5�LF�5L�Non}��D�%R��ͨkh��yJi��7��v�n6�ÉB�ݓ��gJ�C�z~P0G�i���2�[���P}˟��ލ�z����M]܉�2�z���� Em\�!^�a�fy�}<���){}q��5�K|��,&��azM�u�fa���l{8��Y�@k{�����(�B]�>S:�VK��������B�K^��w��`��jN��t�8*��+^��ю��ߏ�=^^=|�|����ж6%�2@xy�{�ev*�Vﻨ_��E��z�OU5�tx�Uȃ� (�!O�!�r���59]�ްG�Cx��;�-�;;�?1����U��;:¸�5=x\�/@���!��	�S‟H�Ys�N۰x���W�׵�����"|�O�n��C���P/���ɖ�L��)=PU�m]K5�Ƭ=����/�ױΑ��m���t��8-4�r9��BL���9�}{�g0�(�R}��rU��r�DKh�L,C�P/���NE�����T����,e���A�0<v'b���1iㇻk/���w�b1����J#a#��@��앋�e<U��U�c�}�뱠
�Bf�GC˪*�[�����4-�	���d���~��L�"E��dر�"Tm����~U�����V�G$�����V}���v����O�bYg���U勼yQ��z�+�!*.�[���y�.��������A+6(w3�L�e��S"�M�P�u�{����h�����1�zP���mV����oxX��z�����!X��/tD��na�������ih�[N��B��zx�1�EU�C��e���L��d�O:�Ў�;��_�,��|�.٧H���Jˢ� �ޅ)J��31vL������3X%p�Si.�����+��eccHq�9s\�ǳ6�9��X�Rfb��ށu#���n�d���7������S����˨���XE�12#���S�u{ &���E�>
�g�ܔ��(�7��֋4b��p�T����e�SZ�3����P�nq;~׉�O�^���V�J�[�{��v��W����L��U�{�>�[��&y<��
��<c�I(�dS�:��D�C9���N	!��'^��Ǚ�K� �N���s�4д�5Ɲy����#�:9���vB���^�V6L�F��7Ӱp'��\�,�ϱ�͍��k-ƕ��|MH�U����z����H����t���ى/�^���)���|Z�u���O�	�v3�9�#jL׉�grӳ�m�)���D�����W�W�+䇊<��}���_�;c��T:�\ΰE�DcJ�o�`~9�^q�MFێ襥9�ӊ!��wW�G2�8��P�<�.׏��d��p�ݓ���U֛��fcCX�~���>h*:�5��a$1�|Pt���#���g�Ħ��n:�s�ˍ�;���F^��8�o�Z��uJjF�Jި��yk_�p�[*ɫ����M�B��IVr/�w#BP*�<t-�זJ3i]��8&�X�+��5�v���neѢs��U-୩[�ʎr�uu���=.�i�D����[�oH/t���Щa���l�}]r[Öī�י�}ɨ�/;�l�[m�m�}|���������ξ��W�.�`h3^�qK�JK6�%�M�m@��>V�u\a7��>쿾ӡ��yyy���q�-ֽR	y�t�蕯b�,Ӹ��{����a��9�PR�O�H��f��9˴c}\�4��MH����!@Mmub:$��1I�>`���O�ж���N��×���ж��{s����W�>�T��/�9F���gؠ��?)E�<)X��X�P�m�(�5̯��g�9���� dWO�հƯi��z쏪�(�$E�9��r-mo�8��PQ3��Qv�oc̍������ �g(m���s��h�phK��.CsV٭�&���cҢ�42���oL�P�$��Q��Dn�`I�v�Xyf�`�#	y�'뿝��b<ĕ�7�q�������ζ�D���"���z����]>�.�D��JWC"�GI�x!���@�7P)�L���}=(�A�	�t.z��位��z�2*�i�f�6�Y���i]�&�F���2��a]1LT�Sk�	Co���jG�;�7ܺq��41�J5��ȶ�
�/�C�~8���v�"W.!����d7K���ٝ�L98�N%X�ŕz;ޜ#\'-%#�}f��n;�cj��25���(u2�黻��i�XS#�9�7�*d��R���ks:v�^ �8�`례�,�a.{�_!R�gM���x|���9�aɊR�㐋�����c����L$M�Y�V�HN�P�g���w,ț.�"'�������=�k�o��s�et�r�|%r��R�(E���G�T��7�z�����nx�3���d��;]}<��:9W%�zQ�<���<SZa,�
�}"0f�B�)�Vk ��Ͷ��o��B&b|�-̉���|P֙8�>1����E>�I�q(�Cv�u����2��9~Ŷ���\t.X%U�F��(7}�)O\0zUq���H�����w�H-�F�9V��Dq�~G����Gǚ_ET;��iOEYg�9NM��ĩc�.�y��QG$9���5�^�Op�BqX����uC��e�(z��d�_���2=��� ���3S��ů5���E����~ہ7�X\]����{e��m��m8��r�ċr�Z��1��tf5���|w��ίNE��[}�5yD�N���.+hV>ڼ��}����BI��\s�i��{j�yR��2���d �<o:�7a�o�L$��l�c�p>��n���>3������8��X��t3�&����G����}ï9�A�lp�h�A_vv����*�H��˴�+���OA��8�Հ�#�ƙ�2��E:5��Қ�:�Y}���l�QZ�1�ĭ�f�R�]t��ӈ\�L�h:�4gt瓜���V6e��x�tQ�X.�d��;5<�vG�-\�YK�y��I��4��fNֱP+:�����4�ɍyK�wV|s�}q٦7r(��Ts0��[Z�cm�P�3@J��H��ƕ���sdM<��L;y���=��be ������N�AV�=���V�[�H�&��-�%qc{%x�R�v�,���+��mX��r	��qj���ȸ�aᠮl��KZqu>8r5�^�;kU�^HT7�.e5F�Ja'4f��(�b!���}+�c�����l�o.�Z�,���ɤI�����.�u�T|!�h%o!1����hpȮ���3:�����gee�_)AH�`�X��+�㎻W��u6!��`�����	L���ə)R�2�)��G�Q�6��VT�CF��k�2�2;{� ��QWYn��1�[�����$�YR��w]�b�A����<�ړ�lNb�uZ��+]��tti>w;P���q��8v� �fKZ�3�c�[�4m9��-v|�`�ŀq����srh�Π����m�khH�,�G�����w�]yr�W�rv�L���zĎ�Ұ��-un��V���Yz�I�=���d|4&iXû�3Q��^,0�'�Ƃ����󜜐6��GfF�K��b��YQ�u+��D���}�R�+ 9hl�z�����-M�f�Z����� �M����5f���Mp���~�E�f�^�{̞D�4�=�����v�Xþ8u9��v*am�i����%�CY[��X�Ŗ���;`�bO���ͧ���g��6s��^��jN�1|2N�Dݔp�R�p>��n1Ѭw�޷0�#8�����r��&�q�o���ѹJ�q���mH�����^�Z���z������AJ������	э�W��5u��z�X��Y�!�e�C����6��!\�Sf��(Q.3��I���AL�f�_REXVB$��خ��uǟXQI[s�K-�qA7L�^��yB�A�[�%oP�wJ�#����C+D��p]p��1�-�����l<fka^����=��R��k{h�	/������f0�,̄ka���pe`�������K�aXp��ʜnNL���6M��p^H�z�7/c�q�a͇8k�R��yػ4��f&ջd�H ��o1�h��k�;YЀ�'�`l��FUn�{����6"�����{rROd��tM�`��嫰�3
yE��m�nv�IqD�7��wVMlf�}ݶ�:uG�&�a�X>���R���s|��3��r�c:��V�SgV��l|�3�2�����c�lV�M�M�͙�o���wm݇�m��w�ڛ>fܳ�8z�ܶ�[n[b���mɷSձ���X�m�cř��͝^�x��m��۵����'m�Kj�FA��,��ޓr��wء���m*�h�1�0\�R|黅�ʃu֬M�G��\���V
J�;[����fo�����<��:��mED�{�����^��s�<����z��aЙ�'R�m��:u�~@�V�I����;�{�)�I?�Ej���L폦�f5^�R*��WJNt�ogN��z.���#Ø�wwv�U��rC�♠�
�IC�a��,ZdL�5ި� m�v*��ў9�]�����[�!��K�lo�n/�߱��@r �0QZA1�q���ƻ¢���o�۔}5��:沰t�ٟ3Z���%���F����^�꣆�tx�\H;�HI@�z�0/�b��v�.{��)۟fT��s�������sP0g5��krg�-��/
L_�"��N�"Ė6�a��Bڪ�sU�����*�,"G����u��؁�V�r�|Wr&�k�S<zJL*vߣ�t����l��o~���GG� ��./����y�b8�����M����bG��[ܵ�^[���5v�s�n����j�酋j"NI�dH�|�+�����ym_�o��c�P�u��MW׋9��hl@mȜޛ���;U���1�=��G�)���Vܕ�ǋ�*��|��[}�u<2w3l糫LC��{��д�yZ�\U��%ʽB����%�br/T��<_k�ݝ̔p��*d��c2����K�&9�y^�����/G�(��&E�ķ)Wv�1f�;5��mH�X�=��W^�
��L%K[[��p��Im�~W!ٕ�`u3�i�NM��P_�k�>w�#��3n
�W5{��5p�̯����W�,_�l�-����,]�ڈy�g��NQ7j���2�*�2���\k��;�x��O�OR�#����؞#�!�m̞լ`d	����Y�]���5�f�k1���p1���~��Oq���j���p3}��t�i���Y��%Vݻ8�T��K\L���}Zj)o?�>��5&#�~�r��������!��H��4����ƹbE(�9���/{:<�ߙ{��1��[�R���7�G_�Q�LD5����긒�1ԟ����+uW>�ztm���s݇��@�I?�qܞ�q<TcZ���@� ��tep�O�zz���W����*��׽;c�hG�k[-*e���]E Tsv(iqvf� ���@�an�O7��㠮�8��q�f�2��ߓ��1jO4�5gr����-W��x�kQ"��ц�{`���V��9�w�Oi�C?�B����J<���k#`Yѱ�Me������t��f���mꦰ� ^��t����:5�/',v(m��qo��/l	���_M�0~��儧��B�N������(�v�
覾۶�V�V=;��C�^=d,���6��X�]��.0��N�����q}/� k�șP� �u�r�Zl\vg3g=���۞M������c�?�"	���_@�!��-]�����05�{�`#��櫺6n��k���]���w�`�'@��H��@��Pc��ҲKT�¢���kݴ1��f�3��z.!�؀�kF�7����s您��R�	A�}�5�l�Y��{=�SU=��Q�&l��/K T�6�F����Qe!��5@j����S�0��}�.�8+����j���/e���=�f�B�1}�2Y��,�ǰ�Z�~xҖe��:��ӪV�vT�.x�����L_�B/5�t����>�UĲl�N�6ߒ�ֵ8I�ZD5�M�����V����wb~	x�o�]�ԑ�8���<��k�_)k�[�Vo�*N7ƭs�ݞ��N?I��.�cO�nn׏�:�XN*=82~C�%�?O9G*�A��:A���1��0{{6]�<D�3<r�~���Ǖ�7�l;Ý�GB�_z���'��g��Z�-'�x\��{\�N��f�_l�pP����-��E'�¨�Ŕ:�]b7�\dF8�!=^�&^2�̚�t�T�T�*���q\z�v�ۭ�x�gS�7�*����}���MQ�c�kst�}��-X����%�@����e����(�H_o&l�G�+D��u]qt%N,�c��<�o4��+9�:1�1������}�eȻ�v1���ks;c|6���|;	�j&�XG��:c[h$r�����@+Ýh��7O�v�z���ŹQ���y����.�S�(��d�гr��H�e�b}X�.�!wj��nbˊ�.��x�ä���±C���8��4-�,T�c�:z6}�C��Ѱ��>��^yG� �_O����-��<#5|]�[��eq�#�1P�Q��xe\��l��u��!l9�^ǂ\Y 鰑7 �Ԍ�x�v�>���^�Y��-J]=�5�v���:��,�v��{>���ȅ��)K9�U+��Q
��ǟg~���{��@F(v2;kw O���?]w�.1C2~�qif}��JF���ds��K��5Z�,�
���on�ϥ�3�x�˝�Ѻ�)�,'�1��xX_l}w����
}N*��<�H��I;���)19qLf��7N/10���$]9)=	ؽq�u�h:��^��/\5��W�a�6�f�w��X�g��"}�"���=)/֩��Uf�e�u�\�0�JV�A�?���K�o"�S���Q[z�{�����*A]�An��Z<<��1<�����Ҟݿ�M��H����ս.I������[��ҫ���.��wr^-I_K���)f��g�]��ӻ������d��)�v+�jq�;Ya�؄����c,#��З�{!�fU�j1gVϿ��Ǯ�&f8�T����=b�<�KM���}����c���esw���̍�-�Q̩�Fs��8M�8_diz�;b����M��5mC	�"t���Ѧ�q��gE��Z��,��	؋΃Lę-���Qb��p*|����j�F��V�ZĄ�Wr dR�s���y�We�G���0{�2��>����p�i��E2��۔��i�T�DC�����7}�fs�U�-��G��ZwUJ`����/!��	�LS�T�GD�u��\��т�5"�`��K�A��))Yj�Qz��㰃;���#oP����Q�<��;�X�"թ������Z�?J"@y�a��b*>HY!�;	bӃ*��ՁQ�����Wp�k<��vB��_���֎�O�e�gl�tGs��T�q^�=+UDj�� `���`'����k��K�Uy6k*�^Yòg�]a����4��P��渃0�Ľ3�%�7⭌�Ob�T럻�K�|� ��7c�B�]W4�ʇV�v��(q�ksӦ<������V�W/�m-^O��$�rl�Mp'��r�����6��O&�"�9L�����ث�QR�4�!X)��cNS7PCg����c����<��\�S��g8�pǸR��s���͝��CV��ݗ+Z�"h�7�������ת�U�7��ի��=\���E���Ϭ$X{o�n�?���~��/��f�%t���,d�0g����uR⡔����� �H���
j���q_�],��ʂp��������u�k�d��[�0-�#T�|{m$}��an/
"{�V��)��t���/�g]��9�7�ԏ�����������O�Qf���I�y�-b���p�}�f�fGަn��s���+�z�EU6��!4��jW"m���E����9آ(1���O����z65cdK֞Ci�הSY5�cЦ�}�K'�[4�ml�{h��~ŵ��9ߏs�����7����[���2�������n|�-Q�gt�/�/V�{>3�i�^��7D��KQ�#�.��W�|������?���?
f�8�W���_uB5�����#���sw�E��q�.M�ϣ-�^�oF���|����Ɉ��4'D3��66�HR3z�!�8�?is"�;,���fo�Y���+���F���K�5�l
�*>��45[e
�������������d�G�a�/V3����O=Y��:����j�=B�f�&c~u��t�>��½�lٙ��U),Ou�����]e�,��%�Fi[\��ۖ����W\�(�0M����3y�\Tj��D|���zΝ�{���k��Λ���u�ٽpx�/�7�sb�W�n��'��顺��TV��(7D����%F��~��h���Q�zxf�S�#�[��=W���{L���5�]� �8��R�W� ��(	��Ȭ�+�sϷ=�}�0v/�	R��T�22w�����~]�ͪ�5O�j��c,'�3�%��j�����L��af�A9/��υ��|"���&�ksodǍ3��t��������6A]����fk��y�T������'(��H���(Hq|�ѵӸ�m]#���wfb���̨��j˹I����9�TE�đ���k��xԡ|��#��q3>7���%�����[�}��Gm񁃛�4GU&��R�	A�+ڠ̸�.��a�ي�8�������2wj���ޤf�nX9O�� =�>�&��T�:P'cW��`Xt��SR�6���S�>챑8è�*�_(d�Tb�z$������{1_,�SB�A���h�p��?�+�?-r=Qr(���sSW^�۪�r`�n�K9���&���8E��?�tDε��ܸ�L�륈��Lm4B����(�;���f���pr�ڽ�z�U7��ڞb�z��pChi��Ȁb䕚cP}:���;���EQ��<����]��Y+W��Y�h�9g=����:(�.;����'^����/Y�re�_W���IS��][��GZ�覞��q8�K�J~��Y{W��ݛ��?�ȣmǼ��qp��'B#��tR^4>�䜷��j5�?>�R^yG+{��j*�ns�W�u�'�k�Qi���B��V0֮79Gc�t�L��.����i����F�,�sfZUC;I��r�\"��E'�¨�,��];^�/�4F8(��-�ן����˓�q�Y���(`���S��0�M��R�=ˠ�}l�%�c��i$�xNw�PϮ��ʽ��Z����Tv<4�0#�{�/�P��0a��nSA{D�e���Uԫ�smM�Y<K��m�[���I���t���Sɵ�J�N��x]�rȿSY~�.=7������K;��Mǳ�lN����kC;��\qiRW�\jP��T���PܛV���)d\��&��]�v��Q��l-4#�]V�n<
j��A�$M�Y�V�}!�9�㛨�{쨙�b��uƆ렧rW]x����?
�K�x�>�ό�ڢ+�2D�!��l��5�2!��b>�ƒ#<3��s#ǧ�7���a�<�N���.�y5]�a�!Һ	�e���_��&tV��n��1AL.1��R�}ͬ�q���Sh�p�nB6��u�C�5o�-R�1�Õ�bv�tz�(�h���z���!l篽��������Y��ּ�����1�.�v�3���|�<SU�R�89s�)!5n���Y����o C��B��ܬX_NȻ�G1o07N*|c��s�"�=�Em�*yJ�w����NR��GŸ��b�x4+���(���@n��]i���ბ�xC�5�yy��/�ӡh��;�3p�Ϣ8~'��|�D�֫�\j
�������N��]sJ"h?^U�)�9	��������
�V}�"�">����\�*��Q>;K��j9x^�������1:��9Bd^�ؤ�iwX��)�qX�P�����aA���7~�}M�'��MC�W�_��C�i5qg��.��lK�r�z����b�~��ed*��Qck\�[������-n���z\�[W!���	�p�j�|�_EŬ8�e�P��\0cXͳ�Ț��}��[Q�ƭ7�ADY�	������0Ս�蠨a��|MJn/�9�\�y���w�f��~+�/�y��hq ixl���+�Ҝw�S�F�R*���P��v����}`j"x^�r�.-o�c:����wXȪ6����+�h&3:���Jq��]�
�u��vѩf���$�VS�9i���w�Z�C2�[\���E�š���=n�6*�S޸����,�1]� %Z/E�����Qa�gު����'� <g���Idp3�8Z���q�
�D� �|�tii�)��s��B"��\���苒1�Z��zy=���/�N����._��]�q��
����Ln��;�o�7�CHȿU���܀�4��	:�n%&2-k�D����<E�*����F:	&Y��Uou� �ͱl&����bƺ�Yk��q����\яF�KS��_�
.i`y�Y����X&��:��zDL��U(��'�x�[�9�����|^����p��}Z��vGo2�~g���Ԕ��$�M/��ۑ%��5s�x�,B~��
wry��z.���oI�W�n�ּ0�#���ͳ������c�]#��*[S�Mբr���Z��W�mN�U��|Qc�0���+X�7_=���G�a�
$܂�������N�ێn{D,��>?�t�ѻll(Ah�r	e
ǿZ�*��*!�sӽ�o;�63h�kUf�`>ɿV��(�%S��w5�9�����!�e�6u��
�t��+na����@�8
@� �ogcn�P�"5�$� �(��K�����X��NNˬ�R��ⴾ=�H���f=̂,�i���v�mk��:�#t���⧌̰1�@�̓�j�Hs#���.KS��Y��'%`PyY\}�M�;��JVR�DY���f[�=�%o(�ھ���N�b�Hc�;k� �_3{��]�������̃�!�[eVo���FZ�*�����Gv�jV[W�cD(��{hp�a=8�QNf;u��!��c���2���:��fF�NP��g@17��(2@��	2�Tw�b,�F��*��:Y�H5%��5;X�����BƜ��uY��K��7H��,�m茧٥��·i^�7b�8r�[���e�X�񉡍�؂W;�5���y�_V@z��!��p�)����1�C�V����d��Y��yg{L����b��ƶ]G瓝^�u�ԥ��;� :r�A`���u�9em4{V]��m�뎅�Nu.�z��V����9wi���4�f�6�+)������2�v��]vdSJ0mm�Sv4�*Q���WeGc:&��K�,-�V��ֻ;d�2"�4��^����֌���{�͏h�R�ܲ�H�[�O`�;��0���*Ӈ�I&� ��ͫ����E���v���8�-Dͽn��n�j���=Bge+�rV��pG�J�b�� 02#��n�W5U�­�;ǝd�;=���s#Qvw����j�A��Ti�`nai܃w@��xL�U��Ȉ�^`,H�#@�꾻�5��}�� ]�'���=�L�=�P����N+[��P���]h�gk��A�KNgtM3j�űr�H�Y�e鎓�q��'7h��v�2������V��$\[؆�,)��m��ěVW|+����u@\w�u%��]<�g=�QbmJ\-�C'k�0]9S���ޗ�ۀ�G��l�/��@��\٦DnkU�$����t����S�I,��}�fT2T�YЋtq�3�d|Pcn�O��C�m�Y0mmr�7V��gs�\�'��륚$�xַS�^��^���U�{=��o;h�6��#�Ҧ�gn�伋�ɼ��cfd���2,{�tмݸ� �����r╦�6�:����]����"��.v[�����{-Hƍ�:ށv���sQJ�k���z��v6K�8��ɧ�R��4S��c�[F�K�nX�%9w
j����-����Yɣ�7��b�Ԡ�N]$�Y1vH�94�l�Vf}��.�G��۹�u�ʆ���{I!_�7I�h���ɼ(��^`����&[Ss��b�jw8-�m[7Ґ��7�VX��Û}�n�h����P{w�)!�<�A���)%Գ#�@��h��'fk��Q7thˊH�S���t�͈��د�J h�ͧO)֚�m�̎�� ��=����.+&��mr�3T�e����Q�)�z���j�v��vYn�39�'yl����+�(fg]uw]x���[rj�=X���wm�նܝ��j�%�)��:��nY��c�+c���ݛ���lr=ޭ��oV��6z�u5aX+:�uc����_�^�� S�9罄�M�Pw\mX����0�=�3l5Y�ZJ�UD��w�N�ظ6�=ޮ�o�%5����{�.�EP���}g��O����^C�7��/ş(�CG���pC�#�e���uE��G/���C-ټgy�����
�_���1���oK"�L^��Z�c}}��-��䡦FN�����<ڟ����Y��?X�}ޖ:�=�}�곐� |�%F#��f��v�;|�.uq�U���.o9p��y�5=-�'���v��kO��r(駷@��i/���=�+x�سn���*�)� ��oL�m���k1^�R7U����H�ג��\�C��"��k�h61���Lgk���Dk��8=zh���J��8�1�*9�lb�,���ssKX*~��M^�,~�	����j�*Z�R�᜜����k^��9��\j���l��Qk�M�~�M"ӵ� �� �9@`��A�Wʅ�jGѻ#Z�GM��&}��o9FΊ�<��5�Ƭ��،b<����}RR�Z��NAqƍ`k�Zk�/�Cƣ��Q�?d��8�_	�{�#	xwy@�렠z4��H��B����@�$dB7��PM�5��-"\YQ�v�<.�
&ko:A���k��|�:��fu_
���G�^?R�g�Ҹs���\j��kx�:��7})
�nfn\i��I���ߘc�9�6���/����btm<�Ձ]�ұ׀��CkU�U��|�>��s9��G��jϼJ��)a�n�0m�?}�-Ϛ
���T5JXe(7%{TЋS6�皰����wz�uݨi��&��`�oJ3����#�~{�!OϽI��Ic��Y��������oԅӯ>@���MG�nD�W<���Y)������Շ�PGnW{2j�D����e�y�a9��j��Hݫ�-s'��"��T�eH�ˡ�S��t0xӸ��jסl�]������v�g�T���ֵ����P��Q<��������\��~T�=6���q�E[Έ��1���=�g�����=覶�	>���x���\"�@��oE%�By�9yo�\upJoVUDFr��G;�*`��U����Z��Jq9;ʅ�ɶ���!ο�����P���&`�{�E������viN�g����gu���@|��8��3�Q����F���ȶ�m�s%[�N;�۵�������P�*2�	\3��F�tS�g)֠M�.�2�r1}1��9`�Z�^��I����of'mwu�{a�>s�	x\�%�"y�_)���&^�C1�[�u�@�\�_+��{x}A+tU�����F���kƻ<��^V_�T^�j� GE7O�.T�1fM���vc�i�j�
����AmL۽	Iӣ�T4�^���ͺ��&��ܲ2t��N[��]G#��-d<D6���}QT�Hk�&��wY�Lv_g/�#'q�3g�&��%���#������c	�qz���{ۋ�dU�Za������5��Wt9�E��=>��T�5}}��t#�f"ɏ�F�%s\hJ}e9����s1�1fHR纅m y�g8��{�:�l9�V�x�}ȃ��nAY�V�_N������G�v��q*�#��8Xohu���rc�f��.+�hJ�CT��J��r��Q�R�u}����YF��o�*�y?�&^��#g�nO���M���sR�F�����.���$'ǧa�z��}�_���n�K墵5c�n��f�'ƀ���{��'��4���X+�c�o�u��5ȿ~���9���[H�y�H��S�N8��{Kl��q�c�5t���F��^5�<�流�z̉k��x����q.�K(�}%~��(��,����0��ލ~�+�U/pE��z�:����5��+5ψ_	X-��)ڄ^f��Wy}!lJU��;�u.�'�̩�k��}��+�ښ�f���j�q\�ݙB��U���T����S[8����/6�&Xa��	�i�++��.��S�j����(>�5怡+.�^�z�s��H
E�cݗ���r>"ϵV�2�^`�^����\JW�a�81��$)Rhٌa(Mu�,wM��R+k�엧g]����X1�I-���:�v	\��j��'��k���C}.��[c1���d��9�4Z�be'�	O�.���7Q��t��FZ��WRk��{$�L�p�oJ��[�\�H&F��âe����Ŷ9��S�3��<+�IɅ����x����c�ǽ0�ʨ
�$�C��Ta�������S��,n��%�]�Y���3]G׊8���v�9�))Yf$�t�WãU���v|]Hgs�5�gr��q�Ǉ|[.WI`�2Y��$���V�V"�!d�b0��-3�LA�z1��zNTNv�!x�n.�vWS�3�6���uY���cVD�i+^�8��Qա��^��I�t&aR��:z�z�:�n�L�[ZUL�Q�ڨ�\H9��a���~������HR9�$B����~�i�8�1�o�y��@5RZ`�*=�[�Q�������=�~�qB}"$��4������W7���53+����E���ó�����X{!fKn��mIK��+P��a7�"D��B&������ʁ��4�#��U����\�{7_�/�3\	7F(��z��5���6(��ϋ���uN�Lz��vl���Zs�K��"�g>f�=Jg*�h:Νyrv��u�Ό�EZ���rܫ�-<��jY�Ά��퍝�|9�ع��&�.��0�m�G���|A��|SU�Jx�"D>�����j�v��Q�:x���J���F�v��Ŕ?2��H��Ր���Ԉ����FD������g�r'����Lol��NP�[�=x����݌K2�7�6��دr�U[��Ze+*;.rL�=̟���mnd���E�q<��Fk6�ů�N5qR����2�[Z��^X�<�x��ΆuO;y�)�TC��0�L���5�/������]��w7������/��{�T������>a�U�������l�T#����p9}��t�vF�ݻڱ�>�םf{Is�͘�����h[��U��>7��!*+�#f4&s���6�"9{N��5emڶ�ޖ�!�ԫK�R�� ;����N�9v����GAT��*>ƒ��f_��Wc���쯘�i�raO�w�[���⧓��	uآGOC�����J�@�*�蹘�t�M8�9~�=�Ĩ�L��S'=�x����K#Fq�;"�Lq���p�Fv	[�sO��.wՃ���uҭ��|�i���6��b�F�Y�ñ�Pc���_|$��t4U��j�H���-f��2Q�0Q�ٺG;fJy����;KpD�=b��b��Hmڑ��i�s�5Yٱl��Թm|gМ0.���6=�π.N�l���3t|�44�!�7���K�:j����ƶ�O���rW�tt7�1_��X�k�nW�54�s��_C�X�	(�������?��	�|�xY�O����3�O�0	[;��\��~�=�uC���##�~���%.47�Tq���Hq|�Ѵ��H�0f�N�G���n�l�:6��	��UH��)���DHȄoiA7�3���7���$d���W�\�vaUG�8~��3�y��4�����SA_��I�܊�mIU����*5��u��S��V��^*j,��e}�s2�n��-�l҈�(��|���v��&V�21���n��XON�?t(�W@�1�mP����욳GP���}@u�<��q6���7S�խ�j��zL��Y�-p���ߔI]}��Y�Wx*Ǌ��%G^����z�ܾ�k�2g�@�$!�:c8�}��	bܷ� ��	��<Ef����u�����I�A��r2�����I�'�����1��{���M=V�5��Q���^�s�!U�"�@�� OBK�~� d�9����-n� �q�x:>�ѿP.�پsC�����i涆YT�{=�^r�N˾��.�m*�u]+w}��C�I��"bt�Iw�9)va��s�N�;jr�/*��܆?��?h�yx&t�s2�7��ħ��w���&Cƿ��G;��ga�B�C%pm��A./�%Q������������ñ�ό'm-�9���U�}�Q��⠴�z4��ꂚGrTZ��EE�!��O��P%�+�ܮE���fs�xu�:�OB�����]:�pJ��(F�7J9�P���u'��G̣܌Z5<�c�N�\DLZti�����ϒ��( �#L��H�+uA������^�[����f�4'p�KJq){�pj"��挅Mx���K��ƻ�kKh*>\)��x���㿡�_>����Ί�P����=���c�)��)��~�wD�ϯ��_N�ql�d�ZU|z�R�a��S��[��Q���Yz�*�C�-�p1��2��P�V���U<�Qa�=>rAd�w�sH�Bo1��X�0���#�����O�>P���^�=Ϫ/|��]=���=�G��@~�wѲe��qE¾��ͭ+���נ#E�5BBgz�̢s˼G�m�U�����;�y�YwoI���D�~�^#�i:*�Nu\H�zz2"D��L[r{��@�ɨj��qg�&m��>�_,�ˉ���|�S0*u��E#r�x��%k��{'�ݒ-��=���>F�KkdK��ɵk�42�O����JM�o+��w���9U9��>u�!YY��M,��[���Q�/xV�t��XE (��pR�M3�;uU�(i�s;��=��L?U���3���'�;Ԋ�3��u��8�
qJ�H������1�Y ���w�t��B�|��Q'8B!�gB��#"Z�u�'��h�9���/��t��OEY)�[��:��Z��u�:dk�i�v�\C�sڽ{	ږ�9�
�s�$�r��H��,�����{ϣ5���]d�&����jEfz��f��2�y�SY�eg�:�C��`��Fߒ�uB��PΥn�v'�~���1e�)�Cǉ���k��4Z�12��%>\o�l^�W���_SW�L9��(�}�q�5 ˀ����+�{W#����ۗ��ӶQL���ih�s�Xg��K�uC���:�1O��lo�=��
?F��R��\^���-O�u�APޖE���c`����'jv�]�-1P�Z_b�9�;�t8%%��Ԁ�,��ؘ�*�Z�V�m�!m�渒�9���ca¥j���%��|�S�Q�tN:ATM`
��GJii�vY춰J���h۫��y�Ϫ5�
���b�(R��[.�@W�2�)����ڐ+�&isf��Ma�UQ�������"]��J��K���	NuK3�,�ȳ�3_S�*��`�`,ץ/%Gg]ӳ�N]ܲq�ѱ���0�V����*��EF���n(]�bʟ	Å�\To&�<��31.x`���L�U��U*h���h�p�i��}·�����������n�:&�{��`��x�/@L��6*)����uX�	I������r^����}��'p��Gq���Rd��F�qa�й�K����W5;ZË�K�:�.�\��۸�=�s���+R���~��@E5��(��&~ȾR%���^;��l@�+n�u�X
L�}�s�}�X�)�p,���f�꒓��%b�d o�D˛�(M\�^�qQ�<i��C�ԋ����۟^���tn��ˣ��ď�> �E��´�"L+�a�p3���[��4��B��^[�ʻ�����8��ე5�t��O�Q0�� �M�Έ�{���p���Ol[\�X���(q��=U��ɳ�v1,�	wA��	e
ǾZ�*��*"b���T���lx���]�%e����CS�Dm���s���l�V5�*Y?Z٦[kk[�:5t�U؈�����-V�j�0��C��D<��[���iQ�U+�WBԎ|�GTlOz!2��-�;�405�M�ڸ��p-�b\�b��Q�,(%���E'��;ҍ��X�8���A}\:K�Z����'�Uz�����ՓrRf���u�������]5�rD��*������R�݆���q_aJ�,ܺu�(|�-�;#U�&,��M�8���\.靠��͊���ղHV�s=���Y�U������$�Rc���ba'�]Wܧ@�Nk�$��Ԣ%9a`%�I��n�rq��T�d9aM>��x�s�pНΣ�u��D�^_�"�H�����w!�u:֭tSZ|1Ɲ�r�i��:��*>肽q���M-ny�1�)�d�^Ȗ]�a���&(Gs�k������^ǌj��R_/W���q��Q7}�����
�AԨdLD3�~��m�0�jcڕSc��Tsr�P�[�蛮T��f��5�}lO|��#"��R,#���O&jT�3��^>�y?`]%� 8��:̪��6򫎮�L=��Y�ҋ�������zB���T���U�j~;�4�7�z�xI��{O��V�w�q����j�����h�_�	���Jq�H��� 5|����d����`˓X�,�-/]fF�'3�|Q�龡��Ϛ��(D���҂n>.8�WV<U꼨���QXظfV��B\�+۰N:����GA}ø��-Ϛ
�t��8�tE�X0A�go������l����Jq`����8���{��C���٨˰����ǂ�H
���X��/�0t��	͕�K}S���j�β�R���5�l�@-,F��m ��Um9�m���fc׺Dɘ����۲�C�1���_�Zn	 �-P�o쾹r�Z�*��	d�X��q7�A��V�>癆I�E1�+o��� Wc��VMл471�r��;�s�k;i#�j\ي_'3N�[B����k��C6u�j�T;�AiU�J����ݏ��J��|b�� [��P�;m��<}��!ty+V'V�D��{��K�n�7waʐu�ynh��,sy�iT�Uh��9;�Ѩ�P�a!�k
{���֗7�ky�t���W5�vk*�ɫG�@+OP�{/v�Q-��� �k�x$�}��zB��ȓ���u�ͻ��������^ZK��7��־ ՗C�S��`�*��͹OC�ʐ���j�V�k.".;&�q�*�ss�8��{]�/ʋ��&ҽnS}>�5�ܷh�Z#qS��.Q��/��w�
��Xr%���C,�Y��J�]rN���O�������1���o�v� N9R<�����	�`V�Ҕ�{vխ�M�+uq��ƣ�R��1�;�1	���%�l:�*Љb�8FᗁGf:HNt�;�+K�۸���͂�na�5<z�-���ceJ�,/Z&������҇�p�C�G'vg)*X�3�kht��p���l�������.�v�7�=�
�Y�{C��}2�VS��^����*^��̭�~��u3{
f%��{כ]��=81�΀t�����(�a��������ӠP�d�N��5+#���n"fŜ᮶�s���a aȀ7cf�)iv��#��ҽȶ^�Ǆ�}����(�dy2C0)�6�;��d[�n������U�hx�iQ�4!ph��[AX�;�P��}`���'�=��&�4T�0�U�P��0U�����X�jGE�M����ڋ6�5��)���m�s3n�m^��b� �K]jKFos�%.9����aZc"�5
����r�#���c��G�8.phr�v�/�jH�fA|��Kk�wu�٧� ��?�gT�)�U���Ǹ��݇n����t��ȯ�ŅY@w�S'iF�.�s�K���t���ͱ��v�$q��׃�[��ƚ�.����O�E��O����z4i��jih�aX
��8�U��!6(�kpXˋR�z(v�c�$���iQ�ʔeb�	N/�ݸ�"���K�52l�`Œb�=鳕I�,V�e�e�����˙k����j)(4fyW-�c���\�^٫C6��RL�s����&�`�{�fK��LaaL���uݩ+�A��U��f8���)J�� �������Ҏ�XTW(�\S4Iѳwx�)����Z��a�ےD��_��{uwUUv�r�$�un�ճ�g&��r�$�ܲ��V��YO���Χ*�ܗ8�%#|NL�8=��:��2�\�nY��ss�6��Z���YT��T���ZmB����VQY�TjQ�嶵T��[y�-LQ��
��7|�īR���4�����V��)�MU�R����*�TR���-Z�*U�j�ʓT�U-R>N�;���j*#��$si��Wx&n^��\�Hw��ٗe�_K�q��v�g��ދ�k��q�����Mo�ӗ�>zw=Ou��4�����j=��^��u�Ԫ�S�x�T�b�S�d��̩��l�{�W�7<eɶʂ$_G�"F�K�P�ԇ*E�d�e� ��̼�ps��UWm�
�n&�Ve_�����glɓt��d9��9��$%��=�B#i#�>���eÓ�k���ywۦ���
2��)�ս�km�����1]��p�z��1���m��`]{wt��ng�:%����do:��a�\�)=���yu��ۧnO-x:�|�[���T��1�iג�xC��?O�>��IjdC&��چv�e�V[�EBiOkJ�K�Ŕ;w�9�7u]EM���z�Opb�/!�T=Px7��fF^�FEm����g�Y[(�錺E���*��aܻl��i��z����)��F>c t��Tʖ��)��꯾ug�������쯁wܦ=�
����7<^_˧�eJW�i#�!m~\)Ӧ?|���|~�������L�d�^,��ƍ�x��(b�J��S�5_;��=]�Zo��_^�qm�"kiPa���mC��jSX�ۼ����E����!��qJ�e΍j��V���nBK�Λ�x�(C���P���`8?�������lKs�:*5::o;2���o/Kw���t��ԣ�jq�-� ���ƞ:���[����A3�\ߟd�ۻuK��V�;)�!G9�}�Z��_d��1���_�T��\Χ���'��F����n<
j�"�	ux*픢ͺ�[�U�ƨ�ґ.�����G�Nr��\���c%܀L���.(6%��5�"�/�;�s�ý[
�p��>��!q�B�=#�+��{3u��aw�2�����Mݝ�K'bTwq�yjR�Zq�W)KqO�܈'�wG�9�?T>��H�^���(
u}j�=�T�g=:u�6�ˏ!����|�����)�}�+�n[U*�
5��U�G��Q��١S`�?(�E����UnX;���}	N��(3��k�Dz�1R)��@��uu�C9��+�u˗[n��V0�wA��rc.��>�'�XE�s��E�Vn�f42���\}��=��[��D��t"�YS��:bI���e�x��wr*�s~�B�nJ#7�z��nym�{o��]�m�c�����T�&q>���j5�o�z��_L$��y7��нv�v�	���g&������kd+�#zU�<�#�����$��r�xtL�� �_������:�>��S�毎��LJ��:od	(w1�����10�ǒ�Z�j
��ϯՏs��À���O��@7t��ҩN�pg������Sk��Z�L	bw�m��Wx� >�)r�.;��m��&�72�wL����FB7����p�c6]?������}0L��^u���^4a�;�����"1�C�\�+��UjZ����kƚ9�bz'�ݸ�,~!۩�ܬ.�e���Ӽ��sI,�e�t�WãU��8ǽ�&6LNY�e��'�ݗK�YO"���K�m֑��x뿏N� <���ڎ!d�����|�x�y*qG��)/�^,LƧ66�ݜdN*�8����dw8£��<gMr �u�v*���s����8���q9�1��VA0��K�Bf7Wz����-��V5#1oI����[A�۴���w����cD���9
NC!��`zh��6����]�V�i�s_g)�,�.����z��u�Sf��%[ ���_'�"g&�T��v±�~zϽZQP���r$�����H�!&uL�꒓��J��">�}(K��*j�7�^��Y1b�[�n��^�H=qv�wg�-ZL���'���!����f'QpZ�=s��O�Y��(�x��p����yq��N{�-ml[��P�mr'+˫!�ϑ�v��c�:�!� e�B4��7�Ǧ�zT�n�=�xzLԟ���������S�k�ܺ�NFQE���`o�#�*b���ոMN�s�.�J��6/U��w��ܛH`�mDM��h���V�*�	���.��(̼Ղ���ڮ��nv��]�Iϭ��־�z:�Z&�۪�'<9���5��H-�R��9�vk_y���s�S�n����0��x��Ο�Q^hs9�]}�}�O�Jv/��&��^�Ƿ熗�mtgE�Ɂ��?0���멅�����..��+��G|�{�؞";v��|��\��g"k�-�9�ʱ���0��{b�'Q�+1�w���/U����o�G6X��M彣~a+�L8�i���YͶ��hc��]
MB��b`G��&֣a�cZڈ�WD=����@MY�!g9|����sV���i����ﾊ�Ag�m�޳_G�3�D���jޖ��~>���=��Ȗ3ت݄Ĉ�*���=j�ױ��'��Q�Up���=h��'���:G�g6�L��z���ԦXځ�b��n���c�&���vs՜S��f�	�(`4�d)=�����{���|������z�M}��Y!�tm"�Hl��a*�dEB;ȃ�� a��!O،>U�Wʅ�kEW%Fi�Y~����*&���%7t�ᜂ�÷)�s�O�OAtE��K헰�]��������*��D/�eO+y�ݑGZ���G�J��ܲ�Ɵ7��Ej<��򀀈ʓ���{��X&=jqI�t�M�d�B�]�<n���8��S�2�Jg��_�R�j��k$�S�}�f���}��y���L����QJ�qrD�D��t	��}��f�wﴽ��ǀ�.p��m�l�� {S�y#CEz�e�~�6����4F�ѮϏDy��_}�G���bs'�o�>�M���df�R;��8��#�[�4�Ӣ7׺_Q�l�?g��Z������Vڃ2㚯W��e��� �ݻ��&Y�@JHeH˰��Z�=�+2�1�����z�J��,�P'^C�
i��/SQ�؛e�ǣ�ר�*z�&�{
<;=�[x�׺E<-dc���3�F���0��w��H�w���K��0[~�<���{�6^f�d���v-��<|9Ag����a�8�(8<����M�c��"G�"��|r��}�E��uٷO<�c۲1GD�{b��|�覷�[�F����{��%��!T}�YP���(�5���
�����cY���i�8C�.^&�5��Ecw�Y|������p�JFϺ4��-�z�g0ٟ�GA���i1���玎��M)�4�� ��n9��3ف�%����aem�Րsza�eH��x[���d2���آc)�ź�`�g@k-:Z�U��pgfV��
��9y��=i�.��5�]��wG�U�b;�����Arm�5#�J��>F>x�4�\��9��u���A���/}[�n�B��1�^��Qp=���	P�T�E-,��ģ������:�);��5;c.�-�6��h^��^3���'R@�h'�:
�V%K[ީ�}�E{����dBL��ivb�nqy�͊�[.��-	�#%���ycE;��t�%�����o*�S�w2�1��=~��S��8U�vE=E���ͩ��6}g�[��c�([�+��y_K
���=!t(��n��.���A�MN����Χi�kM�U�A(�z!���&���>�Sy�g�R$&}{F����ϗ��>��SW3����U�اr����d4��~�_�����	n��BFG�P���pM�ڻ���k�Pc]�-r֞I�ڳ��'
c�/���P~<�>/���^u�L�Y�V�W�J�Z��U�~��f[BXy����Tp0�|w�B��3\�c�rh�i�WH��>�$�폎8�S�B�H�}7<��)��X&S�[���}��#;�g�&f��C�0g\>���R5ϡA���>����T�U�M'�&��p�LuL%�����.}R��W���r��=x�Q��nԨn��(<�eN(w��ٺ+�
V�a��Ӂʤm�8�_J�lth��.+�*������f�4��ݚa#w	�D5�Y彌�g����9�V�+WJo�(���~�yzp�9�oG�Ƕ��<��0�q�Z���r��j�s����I�n�!N�,N!�{8�JϰEF\�wY햏�OW�t�X�ZϪ�p�ىfϷ�����SX�$ViU���ln�j�c<ڴF�_e��S�BpG�#��M�����-�"��u�Z���k12��x����ꥷ̦�1G��lm�C��J�_��}z�>��iA�2�C�V�W��G��	�p�S��o�y���aM���a��fߘ������u�j�,�<2�)`u�D}�~��X����J�E��Y�OS����!.U�Sږy�N�����=���	��iH�8�\����Wí��c�V�0��772��,#t��\��ۑ[}=(WS�!���q}�4�iIV}�Ũ�HY*������㛪z�;=���k���)������b�U)q�za9Y�0��ㆡ�Z��1�6[��=�,�!BC� �/���1�����gOQoi+he�=�1�p��|�}e�2E=�Y��q�acS/�ˉ{>
�-�
~9����k�Mz��i���x�Ό{�mOD@�'|��^��V�	��N��	��|9�{�o��o/*ș�A����rR�<��K���|IZÝ�o�:���}�Oש���τ�b���7��"���8�1�+�B)?��������dר�����q��q>�R�����.�m<Y{�Z���N���VW~�d�^��JD{+��-�Q�Γ��猩vO�3�#@�nc��U��ݕ��o1�y�#t�･f�L�ߩ��JN�$�]B#��"��7�r1Hb1ƿ�mG>�7]��D9�ţ�G޻��Cv��P(C_K5�qD�������P�y�3ry���s�b��i�Ln��,>�@ɨő�l�gv�\���T ]k&�ϡa��Q����Azj}Z��<�;�cX>�/��\�ܖ;J�ln��%4זHM��P�z���Z�B���4֢�W��}�"�x�pbş��Hq��i�[�ͫ�k�S�\T�~��d�Ɍ�4��_N	Q��/��[�@P<����w1�V�5Bڔ��P[G�H!��kha�&�z27Z�w4֞`����p%Tȹ��m�j�RQ�=i:�J�gzQ����oU����9Y����("hUz;z�9hN�%0[s�h��l E%�|����x��i�ܣ�0l���Zq;�X�2hv₭�|��s�h
�}�M��y�y��?HH��OR�Ch����7^1
͹X��L���	�r�^�B�`�i�N�
d�K���Ͷ���n�"m�2=�X(E�m_ir�:��kέ���kr���l�z+-�w$q_H�cynTx��}���k�<+9L"���\����Ҳd�q�ێ�V��0"#V�h��\�����{����Z���	uآGs�������<E�ڤd�N�ُ,8���AOP�BI��2s�.���]a����1Tڃޓ��\�֋��p������z�i�3��HEl�
݀���T%N&hJ��~�Ϋf�oyN��VC�K,�՝ėĢ|9G�Π�j>ͪìT#܈8{�@�w�*!�u_&;�� S��~�t�.���b�e�Ld��c�1�s{&9���)q��`��2$�G.��l?BSpc1N�]UHPy�c�>��C�25�W��#T9�i��.�9�閯�J��kÜzNnO����~�r�.0��vl�]���x�;p.9�|KH�#��H*{�D�H�ѳ�uCV�ؤ���L+#����.�,����V�Ȇ��Q�nX9�޳���'��B�̮�����e��oz�-2�<
�p(�-o�MG��^�c\�|v��9�V��[_w��Z�)b�YT���=ʂ-���}���*��M@�\
.�5��Gf��^�+���ޑ=�F��m! ���k���Ⴜ�<���=V��2X�Z���E��z��c�N�р0�H��T�uy'3\+�;}(��Ho>��q��ۖ5�뼡���_Y��u����<�6̬f� ,�@άs(�o�	u���e�5�T��vRl��B���JjB�&���|;�Q=�xaMAdK&�V�6��ӆ���(> ��h՞�٪u������3al��[N�̠�����V��������2��n��ۋ7֔��}����H�[>��S�����Ж䜫�m��(-r�P����m�{q��;773�����㢃��~��#��D�3?O�:Y_z4��ڂ��sƁ��X/I�h�܇�L^h���,ۗ���y={t7�^�GW�`{h�C�T=U+��>PY���(��8Ϋ
*���G�c�tvL4.���=�Ŏ���H�~yI@���]zS+��_Ǽ����Nn�R��s��tVխT����O�g���yk��vb���91'(!G���rP���L�s�G&uЧ���v	T�m�S���,��]x��<����������;n��ٱ���E2�ˍ}(;ثT�����x-=п|�в�t��s8���)���P�E4TO���э/
>$T�!�])�C�sC#�{U��;�:��S�%�h�P��4$�FF�E�C����m^`s&Z�bx��2�'����ԯB��7P�W��W�%��܃�;{�>8�]Y����̵��K����]�<���8͍Cw9䬻��v��K�`أWQt��9W˶f<�6&��S�Z�o��y�G�t��Ÿ2��g+~Э��'�����[�@#+U>�OO�)}p��/L��v+�i��������]HQm�}��uӽ9
.P��gf%�dr�ܬ�w��'�8���2�����U�{�2����0��C�sDW�'-Cy�m9M-Jw=:���k@y����^ŷY]M�CxnX����Μe7,v-S�Mm�v��2F�Ƭ��eSg�!�q��vQ@�V`�b�	��` !�\��[}%on�:��sY�o(]�Զ#��m�ۃ�SɆ�ϐN�zl���5��ܥ8����o_\w1�C�"҃Fgd��4OE�wd�&�ݶ#�5�-T�5��A5,���Qਜ਼|:t���yqP�;SC����.���ܜ���T��v���˹�u۝�Z��
.�5/�J�A��Q�C���Cb�JJlWq��&M����G2���g_�J*Lb��`�|4od5�n����wc��ڝ.�i��3۫1�0����J��i=�����Dȡ�vs=�\�p�H���լG+!�SX��Jx�Yt�}�3cP-��eݸ�_2�FTĠI9���4������p�7���X%���XVҿK惠4���c��ႳWغ�i�v��MB`��铅����pv���J��j��`Jt*Su�?M�rP~��w/'ɟ6��B�f��35�W�����
���{�Z���E�M�U�Xv�/6uu�6%]���Vg{��.E+n�ͷ��U��n�4��IlkiWL��/�����L�sF�@�}W�g|�p'�Su�X�2]�W� #�wa�m�If>9� �����v���o������ѻ9��&P��Wcz0������ʏ�����1V�ejԒ�@�����,=�m�v����Lɨ#�b��5�Vc�1DoML�|{���!nF�f�j��\hɭ>ΕnL)�ڽԭd��Գ�)L־'R��N�f�A�wئn(��S�������ͼ��n�-��|�Sz ���hq�K/V��75�x�:���͡�0nv�̾T�o�����{J_�C?XG��)nS�:�X�,��s��O`��E۴{��RС���Qj_d�ŐbW�YE�����kX���T�ʕg�6�s�q�|��%�.����J ��C�"X� ���i��d�\6�%����ށ$kv(9%��;���e.Zj�l�$�kN�ڨm�{Kd��+�������W;��#��x��̠��*:ٟD����Y-aظ�f��$r�nU����5��^s��+���r����:^<vĈg�
8m�"�6r���<f���xI�ĪH�RI$�<��
�� ιλ�J��i��Ȑ�(��I5j�E|qȥ�=]J�V�K%�*��V��U��T�Z��QU���ZV�<⪩J�T�R�+H�jkN��T�R�VU��*��R�����]ۚ�J�E�ID�ے����,R��������*UZ��4J�J��-�뚊��V�qZ�JZ�j|ܑZV�&���i$�m*��i^9ʴ�V��ZV����7%j��jV��Q,�+U&�GS���Jҕ%��*�JV��]�*֪KVKKV��k,��RS�r��U-Z���5�t�롓�lڱ��v;����ԅK�M��z�#+�eg)i�w*�O{n�6{z��¤�.CV"�E"h�F��3�J3�W~������g���٠�P�1�d{P�g�fQ8z�d�{Չk��7F����v=C�)?��I`��},���MP͊K{�@�Rd��-��5c�7�(�}�v+��k��{�j�(f�&��x��s�"���'Ccͪ&u��fE�AN�Y��m�Ƈ΋}�xסB�q�ϫ��K' �Wp��z���\�>���R��Pgj��Dz�-�\�r��OQ���P7��B#v�e�Q��(��0��= re/CN͗�$L�U�)�[Q����S554���ca��[���K�P0Z�]N�Pώ��-���SY�C���Vr�BJ�ؽ]���c��C��0�&";��������jG�'��6g���9g��|�ٝ��[����w���ځ��B���5������1��G9V��\ڹ��	Zg����zv�;�5N���[μ����)���T����I[+��qᐲ�?�P���k,�E�9P�LPS�^�םi���g��u/_ڣN�r�
���H����0� xc�* 4}�/�N=��2!E*��G|�
ôI�+?]����'{�)ڦ����K���u�v�3Yڦ��!�EEN0pY����]I�wIl��^���X���v�o:���Ϋ��ϛ�ڃs-��gRx�vDm��R���_��r�v���x�ܞ�y���߷�n۞5���c�ǔ�؞EWa�.(Y�\��2Ysu�('kg֑Ϯ�saIE��.�['Z��x�}l^���a2���l]��K��-�������.H�y)Z{�t�[�U��@��?�D�P��W��GC�>�2���N�oP$걸���&͇��(�q�����Y�|c#fN��Eb�A�j�oHRC"~���k�Mz��p�R�����:X�t�B/��K�gg޴n0�S������|��Q�`��B8�8="0+�`�VG�'�c%c���g=`��eACWY�d@���,丶6�3_.�)=PV.��G��Dv�q�MO*��"�i����`���8�8^�S�{�=w*�a��x-r�ި,s���|SU��c7��:����]{6]�3q�#�`\�{���n�ڒ���zUnX;�t��Y��f)UY������G"�{@(�r
ּk��(#L�e������]lN�w��������n��wU��c;(N?��iY�TC��IY�������m��9૚���U���'����w0��ѵ��A}��2n�{)�C�q������4'^�3)�*bu�}���.��-#���y�S�h�n�b@i;�����N��X����յ�7
\FV�]F,ɄeJ�bu�V�[��{GhȾKΖ�*��ˬS��o�Nw�~��BL���-gV�٢�ò��8G7yb��yg���W�]�	Qv�@��s*�JQ��e7��f��k�7�����a}YbS,���۪��0I��^C��w����F��f���?Vv��� �&�wPz��4��1�0��Sog�+�6;d��|\N�\�}*.s��Y��z����]�<hK�j�q��蠫z_ z\�ZE5��i�����#g`N�E�e���˿D1��hNqQ�Ն5]�ȖRb�oOa1B(*�=��_QL�׮��4	��Q�]����C>=�v	Q�H��s|*�U��F�q�Qǝ�2�9�?D��:9q�8{���3p��n;�8�xjQ�����-�5��T�f��8S�^�}7���mȏK�ss��q^�?;�6wG�t8�(=Q�-�
NC����|.��խoL�Ji"�^}��C��DQ{�>8�p���3C�ByF	��F�:Hu{�Mrv�3a��Viv1��[�#��T�]C\��]"�՝��Xg��>h�Qt1��U{�=I����X�w�a���2��1p��%��Lû�\��e��XΔd��E����;{/P˓�D�O�R���*U���g�<�׾9�P����$*�N��79�
g��F��R��=s����5���"�q�J�:�"�qf����U��zb�Ƈ�/{����9pA���O�g�W�b#}?U{e`���=e7 w2�R�٧�k�zg��G����œ���P�-�{�X=�Y'�fIb���������J48�Z����a��Z[.��r���a����+�� G��@�{&���Fh����	��0n-�{��P㳼�\�|���n=���*�Wh�^��L�����3��5��K�z8Ϋ}"�nl��b`����{*�x���d��Pk�C�"ix�K��y���[zn�ձD:H�'�:s���؞�������5����y�ڪnl�+Ӄc#�s�sw,ǞV4kY���R^5��r���v��q�%R�Ģ��]"������F��2$|�6O=.a�z�����k�"��J��"�MF�{'J3��q�b*4�0q!Y�0��9�,��@��|���PG�����-�*�<�(�u���s�G�����&o�1�����rS��ܺLkm�X6[� p�4��B�[�0�Ja�c�A�0�8Ѓ9ǒfe�r�����&y;i���6�W_�bH�h�R��jw��\���,���g�v�-x�%>�j�����ѻ���\`��m�"tE�d����vo<�=�Ȫt�&�wV����[bZ�u��PǇ�P�|7�s^��v[�8�:x���೤�гr��	�����;1I]dD��`1�q�g���ӪO�uB4�PZ[�/%ν�S�~�2+	T�m�gOAfϢ虮j����N-˨�7]�;C�=�������_[1"ޓ�i�Ōbq��H����ȗU��{P;vߦAǹ�!�<yq �ip
z��}<hHN�P̟��i0N��_)��~<�6hj���������`lϭ
]�)��,����"�{W�&y�g�7�_w��3}�|
J��^��	(|����P}$���!�~3�'}(�z]~9�I��覚���F�FN89� ��l�-y����zj��!?7KT�&G?R*_O�t6>8�@�>�S��H�D��b��,՗���uF����h8v��Q0��2��p���I�=�����(;)Z��ds�ט�52�v`�x0wnf����2�B#�`e��S��u�/�,z92�*{*Z��w�ՑG,N۲^��2m���s:!d�{�7%o��D�\����p��ѱ����Z�d���Q�43��+J��2`t�
��g�[J��"�ټ��w��f�oSȻ��[�z�7Sf���=iN�`��O/Q�L�����:�o�
�er��֩9����Oo�q\�x�WwL�Pz�-\���\�9
Y�V�i�aj���n���9���t�뻶6����7t�Z�4�2<-*�q_iօ\�G��������_�������nZ������(�?Y:�#�Q3䍅�/^�j򆣒|6c]ķy�d,p�_Ҹ5�p8�2^D��C0+#��j����ԭ�^y�5��e��^-��Ϻ}Hݍ�S���t�����sí�@ŞF�r[j9q�[w�!0-�"{�Y�V���ڣNo�������/˞<���^����۱&��ǿ`����cα�{Ȫ�a�.,Ҟa�$d�6N�/!x�=9cN\����c�}�ˤΝ�f��G:h�	���tOg�<U�q�7���~��]�GM{���Y9u�����>�r�����!@�i���bf59�TS)9�[��uP��Q���1�F�oC�]�B3"ayd{�*�����\�gAr!��'!�0,��4e�۾����O'B����Q�~Z�`oEb3bϕk�1j���z�#ځ7�ȍ*��t�מ2d1g����u`��o&��C)A��ӗ}�t��n��*��Y2�3_.�):�U�Q+�2>>�U�׽+��s~�`�3nL�t�W$qfl��b�r�{�����t5o�^���亱h��6��rl�Bnv>��x�|����n�̰,&�Y���5�]I>�m����9ج�*�+4�:cv��y[�z����=�K��rm�1��l�OTw��]���ۉ�;�
�rIqSY(��v�y�e�wAN��Ρ��!"����(ͳ��%͢W�C�w�g��Ƨ��b"N�;D�|*zj,�_�c[��e��vAc/A(A���$O�ǹ%M����,wq]0�{��)��d.����lX�=L�	���)��>:�����z�~��ڣ�\�`�6�wW�w��_g��n��p���'��@*�'Ųn�����z3.���o	��̵)d��%������W�.��j!��V����%ړ�+.�X�c�9s��Q�/��H.�=#�GD��&9���Ev8������@�=p�E ������v�JO�g�^�����J�!�V;\��h�"C��}%�3��&���ü�Ѭw�8��(8'&����,Q�b<g�R����q� ����C��H��4��d�[��9��[�G)&�B�sC#2�rz%ޭ,:�ҟ�`VP���O�Bz_�6i�Sm�����W'���B51�dԯ��lf#Ox��\�<��ǒW��$'�tʍ"b!��
�9#����2%��}�1$���
,�y E=@ӱ����\��+�������;Q�����5z�DRJGm�7,�wav�����T�{e���C��*y�P���AO����Y��:^[�sy�Cd��,�f���l�1MŻ����	:a���[�Z�݄�UFg��`QC�T�+�a�C�R���'�T��A�咧S.}�y�x�c�N
�����2=H�6T�m�g�k��>&gZ�H�v40nb�4�[��pN��x��d�كt��-�(�ګT���466|��t��Uu���_OuIK����c*����>�"U�n�����Nȷ�"�O��
�хf#��#b�:�������N%�p��ai8�"�{O�$C�(�؄{iA7Õ%	�5(_8�D�H�����R;��m9J�����5�E����z3�8�t2P�T�A�/|e8�{.��ỻ"��V���J�X�^k���GhCzPm�9K���.����n��q��Ҋ����P?ԭw�S��]������/w�j�"�xl^ꎕ�)rS^�qI�<�kw4o��PD�n=��Kܪڐ����\�����m�����9�T�/5�yc��N53(2k�m�����ֻ�;"�6���ipzz����������D�Yp[=6���GD��oE4�X{�ہ'�Ǽ��D�묣���T󙓳��85�H�,�� X!�eL�6���h�U��nygL���~�`���M�1��`���927u0�3g��m*Ėv����@��J���azLSWZ	h!�6q�s:���}���gޓ�m��$6�8�m��1s(<��;lM߮���������{����p��^}QN���J]��-g�7j�4ʓ�eE�&Z���vvm�ު��,o�׈�A��j�#�E�� ��HBپ&��R�V�-}gc_i��|c(�;:��fw5 ��*���z��mm�����:ǡǅ����Y�O[X0�z�b	ǁƎ�˗tn�k��3G�gd2�0��W̕�[�˜�꧞�w��3��=�LH2�J'ùn9����F��}V.uN���w�Ϳ�o��(�.����5^��V�\�b���&{���^C�2*l��ɵ�mY�&}Z��zav�P:8��`�Vmi觙Ad�l�VQOtEA��kQ���؍@VdY�=�����fjZ%��u;����ȷ�'X瞲X�Օ�6�4��l3�w�쀊�%�<�M�Iz�їS��s�������<���y[��Ci��x�aa���;
����W�B6![��ǧ�s��)Ф2��w�|	����Jbj���-q8	|v
B�2&�GPc�qS>h��J�v�>�ޭ����q$��t�u���Z{F��Wq��f8[v�ice�<��W��eL����L�O�)<�N���!D�́wr�ũ�2~|hG:%���o̭7VF���ӣ\y�|��ݿ�׋U�p��R�ց��#J����C��7�ClO<C"���ĺ��7<ls���㦦���%�u�s���� m�ְU�	&�ނ����	U��>��el��_?+Ӊ��sz��r��!���V��tòj�'�ǌ�^�Um��{�6ٞ��Y6֛��b.�^6��\^�cU#�3�Ix��:R+6v=*��|�hf1Mz��6ގD�-�3j{,������iM�IgG����;'��k�v��g�x�h�M{U�ͨn�k�£BSpc�;G��*&�V�R��ݞF�<�2'_�4c9p�^���5^�9�f#ڟo^F�j�}}���V��]�[��+���35��f�G���$O�آ�d[r"4$�vq��Af�  �,
��0�,�M㛷o[ȇ1�mA�q�Mo[�d3��2�r z�O0ڮ���hz�C#0N:*�%�������尦X���g����v��-��,�	8����]�kFv��̏�E%T,�nX�
��Ξ��u�w*�*��N��9Gw����݆fꆌ�P���MZ�6lek�q=�N�%��s��[ 10��V0GJ8��N�8ze�(=�,�����˻[#ξ�oj<S�r���yy��ݜ�W���E�u*aM̭�������Xr��x28
V"g#��-8So����	�W��r��uoK�qU��q��.�S5�K(L��i�C���&͚0r�[�=۲�pq:���=�UfAս�a�l����$ˣB0v��l|��j��R�k��ː���,N}��$䩷[F�ʈF��jV�M܏�)�V:u���:Й��6M�G�A@H��"7)����߻���~�G��a��L³�W;+��ݼ#�9�H�qi3/Kv�n��r]�Z)gTl�G���F�9�˗N�b�ES�S�7�#�����]2Q#��״��ș��X�����!��k��ĕJ��Lr��ދ�����Gt���T;f]�]��f�`B����jax%=�Mot�(d�t}x�T�{6c$��ft?�[5��Զ*J�q��������ν�Uz�g;'jo���%�I`�,��j����3%D屪�
J�ع����mJ4k*�P`A�k>�:ٻ�ӷ���ɭ���:��t����r���zƙ��`P{�^�=�O/����
B�i�V��sy+xnE9��.��� ��u�~�Q�����F�ǋB�$+����k���}W\��i�S}M4�+�*Z@���ݓ�t��7T��T۳��\U^'ʺ>�pMaɏ1*+%���z��`�՜e�����l̮�jmgJb����s�d��SD�B�denV�;�R� G�0`Mn�:��.W�١�\��̤ͬ��}����}ăD_n3S$�|#���o+�CS�750����d YSl��d��4O:g���2C�R�U �Ψ^�uÝ�|fD�^g�!i���ʣ��ިI.�.%	E�ڷ껃kUr��͔:N��)��ѼM�c"gwi���,���:�͹c=.4^��y���@>������Qa��ٽJ&닕��S�;&�*�D'	(��Ђ�1:5q �ڗ����)�y�����
�hziV��"�����Ko��e�)c����ɝC{$z2;IIر"�o�@2���].�����+�B��I4�q�X2^e:���O���w�h�z��T�R�ͻ�����^����n�0��ҍ�c��fk���<2�"�@f,���ͺ���o��_�n�[@h+], ������e�²�u�gD����b3�.e�8��F���0_k��L����7�ww!L�yLl8�+��P�Ԭ��/<�iUU�j�Ig��j�E*�k�Ū�E�nR�K�yYʪZZ���	*IS*EUJ�*ʓw�l�IU%54KZ�)�H�G.,ґT��R�MZ�K%j�e�sQʢ�JԖ�㮜�jj����%�)T��ZX��YY]\�VV��-*�Ԓ��J�Jk�6咢ҍJ��

�Ul�M[QT�+KZʬ��ZB�Ѫ�m�Z�Yշ�S��+k��V(���j̥jՕ���5�+b�F��nN,�V���=�׿�O_����U��ϖ��]��A/yS������Y���yڷ��M�Z\�Ƶ�(E��+E��c���t;��Y��}UX�������Ο"�����8m,��mx#2�2t�q��������w�7ߣV�>��8�֩���ܭ� }�\m7���o�6�WO���C��~ܭ�r6��&�
,Ɲ������I=q �-���[L���J�{Gl[�+�i\��eW�ȼ��[��[����t�J�0X�l4��{-�_wOs�9kk�Ԧ&ɬ= ^'�)��\2u�bAWM=4V�����V����p6$#��V!=��aR"l�ngH�ݧ��LJH"�b�w;����h����|;<��b��6��y��o��]���3��+�[���q�b�y�߅�գ��od�*h����-wmʚ�Z�PcT���o���eL�l�����\��'Ƞ��v�b�`
��Ŏ��^/$zӵ0>��Z�G���4���k><EVf�9]�	�R�X�[>�v����>S�on)����i5w]腢ESHd�ǆ��ج���w}����k�ix^kD��1�9ᢦ�ú��g�=�`��ܬ'�;Y��:�O��ñ��|]���.�Z����D����%���bM�f�i#X�#p�{:��=x�a"�q>M�j�:�oZ�ZG�e��W������oG���_���<��ipbW%KM�[*�66�f�>^#���ms�T�j���p�َo���\Q��c'X��"6C>ۈ�U9&��y���L�Fq�ȗ!mz8o[��9��L;ϒ.�'ZD���ǌZzrC��bt횝ҥ�O3;g�����ͣ���ϫk8#S��ް^� ���Ǣh�sEw,�cKg&�Ѱ��s!�7'2�4�M_p�"��OpֵˣWqոy���$��"�����Ó�;OZw۩�ɞ$۶C�F} ��}յ�ֲ�Ov5��0gI��9�" e,~���r<^������9[��ٟX��l�~��J8$�V'�r�]�2:^l���A�� 8�n.�́
�`vcgm�M�A��6�jH�h�����8�_�=�OIx�� �T}�������$�S¾;X���;W3sf����S�H���l>�:���p؛�����2�Vw)��~-��<N�b�S�!r�x�ǻX)�*�
S��է#u����Q��eőV���;Y��b�w!���-=N�خnΪ9V:y�ѷ��'��9�v)��G"�$���߯:_�*fO�nV�.-��hX�=ᣬ7d�Dp&��^��h�č�����v�#L�t�)x�k5>��m�f���5�e�9���p煸�ua�L�6%1*��-�S���t��{��ō7wM�t>W>���F^�YyGϊ�X�`M�.�W\�$�V�Y9@��w��Al�^�ۓw��	��^Cm[l4Ժ�C|�9ca,9��X��ib�r�B�u��f�l��3/:���uO�>�k�AM�����ן�%�+1���%�F����m�6�|0�녻�˝ټw�S\�[7��{��nsy�24]̴Fw'�/j�.�c+6��Vkt�曞��>e�F�른.�`�[U�7wW�R�E9��x~��;��v�ϻ>H�Q����e��g�%����x��|DF�NI��2;p��KUZ����;4o,���G�Oz"3�[�S����QR#�H�Dצ{_L��En.dG麣���U�����U���װ<��k!isi�݁�17�0�@[�,Һ����*J4uk�_�����!�4��ã���)v��s0U�B�\��U%ٻhM��Z�2U�U|�bC�M�Hf.���;U�E�M�){5��q��f�S:S�h��f�&h[��Ws��G��7���>e��.{������tN�Q�x'KgS�e�cv�\�=�ٍ���׻ژl���i�mF@��H�Oi��qA��ot5ᑵo�aݞ��^�1:�A�2�n�a�Ϝc�O�� "�5k?��]u��M�Eo$p�e�#�r�>nV띴���k/X���U��7�����WB@D�U�ز�/QmD�G��U�OS(m;��SGdb�·���]Aj̘�j�qjV�k@�ǆN�7K��e�q?Π�{+�F�hnz��w���S�X�5[+5-�@��+��q��ZrOeT�٭�$Lő��V��y٣*��7CM�TL��u~��e��ʿɰ ����T�;�܇[@���
�fͺ��FZ�=��$AM�dhO8�pfi�CNw6=��.����k����R�~[[Jk0#���c/��n���F�P��P�8�ŋ�+k�yz"�u�h�f�߰�NKUqO����w}1���M;<�V�w��p�\Nk��;�
��sf]@���e	�&�Wt�u����pcܡwH�Ɍ����D��%�s��]x����T"��{H����N�3��(�zXq�mO��-}{2F����+���,7~����� �F�xI[9���g6����ٲ5�\��ѽޛ��� :��!v����F�%@�E[)K�ln�#k���5��U�V�k[�3 �;>wl2��#��o�<�=ұ$��S*��˥�;�b��R�2��%�<��~�zg�R�(�}3u{�x�>gtcN��ë��j�}���8m-	�z_Q�J���ƶOT�X:o:Dܥ�om����֘���v�~�}�k��1�6��'��S[�r���=�Nzs����[�-�ė�o���Kia�F^�X�0/�p���޳�uqZ�<�r�b�Ų9��u���O`J�2�NÇN�#G6��{����$Z7^�,R"l�����9 g̸�(EKmxO22Y�ʱr�F�����gZ4a���!�Ҧ';�e��r7v_o���;o��~�]�,y�rt��xi؛O�+jc�
�^�~����X>�|�N�(�΢P�9)�:�Eu���1��m�R4�d�e��\SC���R�p�C8J;��!��|3C��l#�\u��j?�Ϫ��z��]uΏ���ͧn�o����x��R�&c�g׹Y�x��MI��VN�X�&�^X����̕ru[FZ�x�k2��nU/}Mw�צ"��Zx{�ޑ]��`�SՓ������:r�iW�C;��e�����R0�W
̞6��B-�o���5k�I�t�����*٣v�%��Ѳu�ޫ��E�6�;g[4Vl�!#Մ?��4����x%ZT�Ú�U�Q7)tlSÎ�k����F�ot�f�� U�k�����Q��.��Ҵ��[1�~6ݜz���uN%���W�	v��w�>�Z�7���-��ʞgfj��͈ẇ@�A�q��1�uTv�fv����DBގ�Ǣ��n��em�i�o�w�е�h�j��+2oY�Ł|wN��g�>�����d�K�jBd�ؽ7|�e�j��J3��c��ު��������1(����#�6\�-���w��%��M�"V쫋t�.h���R����^���<6���dҸŦ��G�]u0�2�2_=�y@&�@��&��z�.*K"��76��Qꔖc<�{\2R���*L�,�̚A�� i��`��^w9��`�,-�����d��i<On5x��1�,�y�|^������Ö�dv��c�|#p��@��l=�����'��®�I�[��W�&���tP��[��C��Y=�:�Vg�p�����1�L+�G�9�z�J�9����O����h_:d���2���>��ȉ�y�����!A����y�I�r��%����\��de��S��d��7��U���6�P��s�݄F-�ӊ���8��)��n��)�+w�t�������ywD�K@��]ryzrh�텇���Y+h���U�S/=����}8A:'e�<;�M�"�� �k�-Q��N`8��kL.Ñ��`�aϓ�t�g^�>�|�.��eQX�x��4�0Sl�kM?$A1P���u�C��~�6�N��|�W��[�[C�c�۬��5ψ[� 0��,�Z=��l1P|��-���=ֱ9�qۢS����u#*T���$m�ҏqπŗ�lK���ST�O���'Ɲ�����؇��Ǌ�A�%tz7#W�eX�P�:.�޺��ٷ����5`N�+N����Ш�:�7���Ț�͚���6VY��rp�6�/f4�V�Vo.ޮ���.��\ϼφ}�e�n|V��R��G-�+>�<���[~�Hݧ������lq;����aV	��I?Ve�"��d|��F�C��l��v(�uI_q�[�m-|�IaS�]q�9������?��:�/��u���v9���?^���ɂ����m���3ٹ-x[)��|��Q���,���-�s�7�7ڑ'El쉬�$|���?H�=)Pc=�Pc��Cb3Y�^J}\OA�G��"��&����3�i�M5�8��,h1���.0$������;�Bs$��y�H�m���p�����G��yjXz�y��^�=k{c�^�Ѻ�7������ݧ�-��R�P��
��1���*It;Ҟ��{����%<h욋Jbo���:hw)y�Ax))��]6�a֪5[j�����ŶB��q� K8�3ǭ.�&ejs;Quޛ��=��㘫�~�/U�8W�B�W��^�#��������j��㝾%��Q�0�k���������Y���!Ψ��9�"���_.���.}s��y�[�9U}[�^�.�6=`�P�[-{/��R�j�	�7uz��!;��ŉmj�ݼ������Ÿ�'~�_��ڥ��1��8R+=79�Y+1gyɋ��C�c����'R]`-��eex���{몘?u�o����68잢9Xg����'^�wn�|���z�2�����ҫ�G$^1��fPv�c�\�ѱW�K�'Z^Gq����j�$d������ߦW휧��:l���K�%/��,��v����0Ӽ��i�������R�	��"����~���c��m����ϣ��GG\��ǞGJ�Uov^z�c��3��� ��4v9��G$nW޲j9�����=���T���jl��2�����v���kq��'1e��>�Sux�z紴���F�k>-ϛ]w(��n�ˈ����lT�]�E�im<��������g��R�:���t�Ig�������Kr�<�z�Ñ�k�/�/��N�c"�ck*�U�7N*�H<5�%/2�Bx�{������R�{���Mm�㵇q\�$�j͝��*w$�*lٗ���Q1&��1)M��vѼyW[���s���{{�9�n|�k%���7=�l��a��m��rfL�7Pn�-�ce,%9�Kn�wX�0�/���œ#�y��v���<{����D��5�)k�nT�k�Pny�n^C�^��U�:�(��SdFt�x4��q�ogNX�[)���t6�d��6n��v�Þ�e�u��8uƉ�x���M��
z��m�o�(�-��u@�ڊ��ɣ���Wu{.k��◤���mvbM��[[c��|-[��Y����U��e�F���,a����ؙi�q����ù�5m���R�v7�U�'�h�!v��V���l>e���\2lx��XkϱƉ���*D��Ě�V��g�5����T�^�Cײj�����=�v�����>���N T&�6�5�]��;ll�w4�ʢ�=ǜ���l��|Y����� � 0��8������;�׫�WonT<uT��m��L�W�j�Yb�k{ ���Q��+R�����Ą���_��^��9��60��ͮO��N];�S� ^GD*j�p�/y^��k�v�I�ܬTr�f�F�!@�����R�'����ݗ
�&��T�ޕz�*&rh���a�8I
��Q|�k�1Mf1X�r����vn�
���up� ����W������q�*��u�
ې�Q�!u�]gZ[(sZ/����>s-�KR�֜�zjYs)o�d5ڲ�Kf_�T���Dɗ�r�m�N�bj�;�j���;�l�m�ή�]�;�e3V(��)�h��;k�����E�U}v��d�Z]`5��smV�'u�Qr�dƻ�)��ܢW�G�T4���-��ݏ{���!��0p[u����5�P���<��uy�̣ݙ@�9}:��pAJwmr�1��N�00���0V�U��íx����m��m�*��w�d��Gb�㕎�5�6�^�D�l�]�v"[�3Oh4��ʗ�a�x1b��%:<��v��C�ުnN��@-c���N��r�}����R��Rw͢8ث�O[9�]�\�lHi��Ήhʎ���53(��F��d.�L�Zġ�8�\���y��;��Fh�B*v>�WRwLכI�2��,�Y]�sV�2��ǡ�3����Lk���e��ۮ�Eg�e������Y�2�v!�"��ͺ�ot�LrU�nu��,��t�5�`:&R��l����:���P�UA��� �$c�B�.�6ԭ�B���_kLy��Ws�>4���ښ���7`�֔ M�FM������"�)�NF"�M���ڹk"Ǻ��1��_,��7�k�]���試�E{�b������*��t/Ao��j�d���)�m��Ie��5ud�hk�:�|�O�8�Yd�4���ʸ��	�X[���M�B�����%���T��׍�9y��h�s("W����Mp�EuPtv�V���6��{yu����۠
Z��Ul�V�1�t���ٲ�4�ŧhN>&֘FLV�yz��wY��͂r���ٮЮ:���X�ӡ�9ͺ��VԵm%���Ed櫮eU��I�os�\I���J�⡶��7�`�ݝ��p��m��ѱ���i�֌�'W�#j�m⹪r
�ЗB��i�os�=u�+|�z�X��i4)U�xVv�A�����ڀ�Zj�T�r���Sw�ǅ���Q��#y���N�"ü~:=/w�;=DD�bڳti�dQz�� �6���W���[]�6�ǈ���-�6�C�R.t��@�b���&%g2N��A�:π�ky�t����T�{d`�Tq�*dD�;����mdewuL���9�
XD��G���A�x����ڙ�x��V{v��)γ�_l���J���8���r�+�%B�\vQ*�,��V
*��R����rV�5l�Z��R�YJ�V��>#��JLKS�nYZ�&V��*��J)U�Ƣ�jڛV�����R�j�BJ�x�:���j�F�����ElVڙ[+����EkZ���E�����6rڊK)��U��Sef��U[V��[R���+j�eeQ���QEHk����j�[R�
�j�TQ*jԭ[�o3���[ų��Vۗ�V�[VkEb����6qa"�h��|O� H ����B\��G)���TVL!Z#�x�q�1��p]���u�+�r��5�bN���g%�c��(BB;5�Q�unJ��S��i�3q������|��7��a��2�߯ڻ��}^RK����g��_���, #�Vnb�4���ơ�o^ ޹�������q�3?�w�M�O�}an4��@����t��j��/�r������+\׊�Yj:Ɩ��z|�;P��O����w���6�H�%P�ؽ���U�k�+�T�;$�bvj]��"��gI�K�=�sL�07�w,�u���{�u�E�AU�����L��t�"EoPn��L2@bH���@Xs�ű|�����l����2�ęv�w�����.d�������2�"�!Y�8U`���O~���wyq���vfcWe"�#�R�� �)a�Hx�k�tU���m�UUSMh鈍6� �ݧ����\�̮E��iF�I�͐񕽨[�Y};P/k";��Zۓf��V��M�c���J�u8��@���ݛ��e�Z�[������y��L���G����k�b��ƧVt��F�8���l2K�P�r�)���k?t�������7�:+�|�G��Vr�l�4���vE�֒��
��%�p�Ϻl�ɅL'"�OJUr��I����T^N�f ����=�G$���՞es·.~��/�V���[�j��S����_9n�Rn���[t4ׂ�V����a/=ѻ�sZ�Ϳ\V�";��U�	̪d�废��k�	�ᶴ�.z�c3,�X¨�<�{ݡ�h�]����[\n��ٗ�p��./�+U3~L��m�c�&C�;��un�X�$UR�Y]��i٦Q�n\a2�.ʥ+����t�%�1��������h���wR�lW"�nl�~�oD�������Q��ۼ�'����?)�ȸݴ�a14i*	w�� ��6L�ɿ�=Q������,^�oht��޼3c��.eBWc��)�w��F���?��ϳ�����|����ډ*:8�t�4˽>>0OQ�m�� q�֗��)��T�}���'\�|�n�	�Df�ӢTY�"�D]P�cre��.7$�Y*E����I`��闥qD�7�$&jmW��E�Ŏ�^#�i�}��.��\ޚ���v�Ԟ0g,w�Y�rK�ew=�169��.�a��[���yiDkisU!�\ ,��M��`�W�:4f=U��공;3�Mj�ԝ:t(��|���s'M9o�>�����2�䴎�9FlϘ�=?h�"��ڱ5�QĴ\��DW3W��{D`
�첻����A����T�F���i�4�B�C7g��anz����r^=T��u0.�G�x�W$���~*��zW���'�eWwi�e���k/
��{J|"k�n�wr��]�H͈�s�̶Y5q1/&�뫣��*Ҏ;q��jX�R�e�4eMm�n޻�=E��l�Kn�0LN�{
4��7�n���b�~��3�ˤ�h>c|yFab��W1gFm�o4׻����Y%,��
����u ^2�w�Y��G8��#�c^��⍖G�[w��g����	u���k^j�MM��vi�����ž�����j9�u�}�KrD���zVm��Y�V�m�Q��y�f���ژ�]�0
����F���O�]�ۼ�2�
hWY��S�3�%iK��ך&tgm�9wg���9�x\���k�!��ߐ�s�m`ߚ�2<�7(>ެ�%�w��{Kq̴.�p���ܫO�q�Z��@lD��Й�ܩ&<�v�%)M�7CYs���>�l�gk�G�*�W����ɲ�^�������5+-�~�2�����ϤZ��=���鮶�ё[�	�ѱ�������7e�,��	@݈�ȅ��'��?Y�ěo�������E���鳎���c���^�;#�l|�#�`�9F�F��
�S+n��p�}>�p�6��K�舰7��$ws^>��Y�&kh=F��y�M@m�-��@W�.Si��H���/s���o�	�^��G�������M�� +3r��5lvGa�l�t�h;|��S;�T{7\�I�o0?2��H09t�p� C�^�V��[�☍���_A������Þ͑B8��2ˮ�>�j��BJbl�nOH��� �f��cݬ�^���3u�����FO��@)�/�$�HQp�Z��m~�}�dut�u��k��&���%�����[�^��H� �䇎Kk�[Ҵ�N�~�ȼ7O�
�<}yO���\�N� ����EҎ��h}��ձ�(����4e���u[X�9fʔ��i�B�gk�:���I�z����d�og	ׁ��+���ks�9*s��	�$�v;��젘�1j�.�BU����-:���T�?7~
����m �I4=7��_rps�ż�ȵn꽄����l���H�!�����}i���q�e-����jso8�Y���n��l����ј5^���n��mK��	]1eze/��8M�[:�e~�܋���Ǎ���AhwX�{4��
�����ݯV�����ã� Wt����|�[.�g�l9�dY�]����C�z�>�.�;>W*��6^{���pp���������W]=�b|�	ӵ�Έ���ο��M1cmtW�]�-B�v�M{�F�@w��We.����@k0��ܳ�;��=��,�:��B&r!F��vu/�$$�\�{گ(�,xE(�B
��O �fDu���!��~՗�z���(cJە��=��R�^H���!�w��u�1�;�HoP{�ӹ�������&\N]� ���t�%�E����@����o7`��*��j�v���\���*�n�[�]�M�#��4�]/�l���%�X76	9܉Vg
�<���TQn�b��g2����a�͗�/Ғ�}�ޟ�}棼v�s�oH����U�#�\vvw�v�Ly�u���wiXz;�du���/Ț��#�R�4�v���5�-���xh���h�;���ձ�7�^��2��E�$FO��W!%���p�2/�:efw/t�ۛ�컒֪cV�\<�Sq�@�2
��-�\)&��ͮ��z��eo�g��P�T��T�9�!�RˮM747��C��X��zj�Ҧ�hYݧ������o�{�M���CMwcP�2˷�V.-��Eƽswn̰��n�{���ӽ'�s�^�+v�v<z��Ϙ��k�)�¸5�boeG4������u�/d�uRxC�/��9Y4imn��e�.g�G�I�K�O��ٽ��q��H{9�x���"m���j���s��wbS��^fm{E�v�W.��)�~��W G�����m�X;�q%�tn�H��mL<=�yn��;�p��H�В��x�]����J��VWdbպ?:u�\du���tl�Һ��������C��D��sU6���،����5�i>�[�ٺ,*K[�~��6�u�������'�Lk�n`��u�w��e���+��n�l���ٙ�'��aQ5�C��\g��cm*��dܥ!-�Hy�i7:���~��3v�_����0;Xv9�oH�S���v9�^s�''�47\S��u��H��t
Μ"�d��$6����F�J�N�@�zv�V3#��oS���g�u������>�=)S��0o4��==��95�Q��\Eu���}ȓ�[@&�t�7v��6A����f02�&1�pP����~{�uj��"�le�=�[��l��ho*�T��=Ȥ�C=伩�H�zv��͉��Cp�^����2��ݗ��bErHd�Z��c��.�����;rV�#��N[KpA��s���U��I��߽��`��n��{�ř=�����}eM��;-C����b�^�Ⱥ��^RӬQ��V�-���)�r������|o�G��6��c�?Kl�zx�GH�����8��Cx���V�,�ח�e 5V�ӎ��>IH�'��m�*wu���M���b�w��:�$��������,�.�y� �w�n���z�L�e� �݅=o����.�=x�8�^J��n��Zq(CK����9�/_e�m�ݎ���[8,̒�­��:�x˅��1"'_�`-�WÅ��ʇ�d�C��ڛ��ބr�K����}J�Q�}�u���+!������{��?_O2#-����D>����xJ�2st��k��[ssli�U�.�t��y50�P蝯GӸ�Y�����(����a�ϻ��K���{ӿo�����3,�(K{V����¸��V��ݻz��}��i(矺G�Fw3`k�-�GU﹛/��^'�������ܶ���wmX+�sSt���Hm$)�u��ibl���^��Km^��jԋ�z������nhq �=�wU��Ƿ����h���7��������p��҆3�V"�Zߙ�6S�hF_l���}�� ��<Z�{ |L.9ؚܹ®e��xOm5�o-��|�SC��&�͛���؍N�Λ׭B9��z�>%���{r��=��
Ao��i�}��N<�]G��N�p�0��`n�Z��n �=fcM�k�[o���ݦĥ���,f����C;J��.����Kg*���]��7\s�w�}���]{!�CF�_H�b^!a�E�6/��<~�����>Y޽:��{$v�e5�l����+�!16nꋃ0md�u�	,�F��":��NS��9���I�b�<�`v�y��
.��kp���#�f�ڶ�k���u����XF:���|�:}��,Ӽ)j3�/qt������&(Gl�Uu4�ǪC�7\�	��C�P%���*�\g+-Yb:���l����3j^>g��!&ɴ�M�26x߼a�����t�5���A���'{�en�%��x�d6j��\g�]��>̐m��a�~0I���Է��y)�Sy�V���* g����ɭY�0���D�60@�{387ه�3�t���ίٵ�sG}@�c-ճ�{2!��ӥ�&�	�'��wQ�P�Ր2*���.򳡺ʭ��*��4�4{5�ѧw����\ye�(��˽q��M9��ꓣ�b̖�����CG�C}W�^�#թ]�~��e��N��3�pD���R�q6�z6n�_���ʁ�:��7�d⥰f�3�Րo ���K�p�o�ֲH�+W�^-�jN��w�_��Ix��B���2~����׵�C�s!-Ӗ8V���Ow����D�5Y]�Y��a�Ye�F�%S;�ު��Y�2T����h��ީWfl^O�i�Wn�� �2�+�,�T;X����և�mg�������VB	O����}� ��4��k��e�1���n��"��6Z�GT=^�׽i�b~rW��U7�k���n�p
$i��k�ΕP��:0����.���;r3V6�&��Z�x�S�4�F�	}�|<":F�����tz���&���=��)$Cs��>#��K~F�/j}��$"k8ם�2���;K�@�eV�E�H�9�4�4 bJC%(��/��da'��z���4ۣ�����_5P��t�ƮR.'q+��
t�e3��ufe�+^��G"������Vx=�1��"W(mo{��,��,8L����h{f#ְ*U2O�Ǘ�;��<Xd)W��[�&�4�6+/9&19�hח��]�L9
�y���Y�{V� N,���e�Ը��4�$w�n����6�9�Qx��RCA�C
�[k��CuHp��m����-�z��3`rԷ�<�q���4�e�ԻLeN�8��/�Dت=_,��0�tm�n��@e�h��Ǌ����:;3���Y������_s��"m�%$czB�:U�������z����8���1Ku�b��H��:�Ibm�v��am��F��+��<ib��N��n�M�YY}Z�E1�G:�!��r��}��{��6^෰���]�w�������KL4h�BT��t�>7I)�&�ރ�&����;�fL9]�p,�a'[+0;dt�%�h��tM_$Ǫ��GoB��[1V�[�麌��*Ӏa�F�*\<�Ek:\�Tz�o,I^XU3����Y��W[�h��֔3f�r�\��Y%p;6��SD�5���Iz�ݫ�+�+jֵ��]�:��<t!�V��#]w���e��n��ɛ�X)]�U�ޫ���&۬RAz-#+�w��f�h��5�,�L4�Q����̳�'��b`�c���*��c�{p�7��~�H�en+�=-'z�¹yEqrY��렞N{]�ݶ�V�I)���uݹ�.���T��*ѻ����L� �V*���!���������\Q�F�N�KUz�b}A�0���ؠ�4`�F� ��j�nI$��u���a�Qr�Ӫo�1!q��qw��jv�ooq*�z)���e�ʈl%<\
�`�v���ܴ�-�e�#��r��2��@f�*�6����4eK�iD{�s]�ۉD��׊�#1�ʲ�y�D��!O�K������ɐ]KvK�A�WC��'i�X�m�l���WՆ	;��/��[�� �wG���V�"�憉��r���n�	�)8�޻z�N�����0�q�.���K:H󹤋��w*�,�N)/ �
lk\z)U�${�y�����$�Or��p��2��v���r�3:0� K�����+�)]�[3�ǚ��QpHe�[��Z�e
�V�&�e�VС���ї����n�rQlڱ�up]X D�lO����3�C�;�-�{��bk�t��R�5�A�����y�N�n��5Yc��9؎��F��J�!�*n�0!��0��7r��dm<:!8�11Q룔��o�sv�=\h��P��䜜��D%n=�`����W{'l��ݱtj����J���Ll�]q6���@�Q�7�)����r`���X QLe�w�΋�f�e���fq��p����ѣ@NS��9\��s��2���%�t���7����;���V���:N��y���6�1�T+�<���u��ޟ�S�������gn�&����]:�ϯ;�)�+H�Y�Y��P�Vg�g-��&ܩ�7�ܫ+emF��V(ն�5ef�mB����J���ʦ��B�1i����nY��Ǹ�g�m�|Fr���1��sI6;��b�X=\��r��+j�c(�՛�r��&�6��:�Ul)��Vάrګ2�j2�Q�f<Xά�)�f���=s��4>�o6�f+�F��X�7�1�x���j�O
��ʓyb�5s������xK
���aPm�Sռ&[㶇u�gu����p<և���Gh�����*���z�[�_M5Ϡ��Kv����<sgb3��Χ���J7`��@�d�4��Y��P�ړ���{K�C�]���,�w��d�A2/��m���i$+�+`*��4���di/�vs2�-.m�4��=��#TfJ��h��Uи��G�uQ�j�Gn(�Gec��
�f����ȇ=0�ȸ��J����4�L`{�n�|�/(���+kڴ�,q�h܌�Q�A�l�Bޘ��u�f��Co�E�������[��yv����7��"�g�������tu�ιC��������� ���w	�\B����Ҧ=�L,o3�B�҅>����/7��7zwpz�������-�I� �c��e�e����9O119��n;�`��F>E
'p����l��B9Q@I��r%K�{����yYjGI���M9�gM<ayj�����vj.d�8{֩����A�W����}ذb���+�r�u+P�v�����=Dy����,U�Y�e^t��@���ۉ��yO�ڟ\�w�B����FV/���=;��H�g)Ʊd�C5(#�?�_�/�!���3���5�|�y�_x��A=�T�;^7f��Ub�Ff�{B/h쁌����
ʘ�ˬ�[��-���v�����~�9zF�**W[�i��Yc����O�"$�|i��~��\;gw;zk�vI�@���z�ڬV�-��Pܻu�Zbk3!�xnKm�VKZ�Ή���{9$�ym����z����2�R�*���uO+�z'5����F_mik�:9Ѻ������*�֒:+#{a��jqd�o�/Ot�Pl��d�[.-�D�-=���t�9�C�͎7��si��1X��6�G�D��+$G�i͗h���Z#`s,�/��ȪY�F�y�7p����׽�C��~�ZL��IwF<�]�K��h��YJ�n��Ӑ���U$J�Q�/)f�>�#�3`��nD�GN�qV�r*"9��q��H�wnsî�KT���S;1�[��;�$Wf��~�xϽKq�ܩ�s}q6�ac+�=@��U6���Q|��٢'���6��{٬�� Wbtr�(��<���P���5*C���h�$��:�b���ٛ~��.L�/<k�ᱺ���r���s q�Y~+��M�og�3�-���r�Ge�nw���2u���:����Z�"�Ԅ�ޖ���T��9��ĕ�R���d�tdTz�8�mhj���P��F��7�v�I��F��pl��V���Y�T�l��5�r� {���E��v����<6�E1�77Q9�]�E�"�G�R�7Hh��_�"�!a�Tع��X��]���P��M�{m1'huP�)��]���|�]�!�Q�Z���A�DEk�C��D�"�Ϲ
���;E�I�*�ň	y�b���nT(}��>�:�ڊ����c}���NW�cZ�qp�oN��(��]����i��l���1*��A*~88��|����.�ks�5�%YҦ�y�P̀j����g'֞)a�>�&R�mX�`Zݷ�;��z�k���g�+�u�!�x:��&�='����=��F����KM��8�t�hi5���%�ZW�X�KZ1ժ�n�a�)�]k���T�ڏB�GMr��ۏ.������0�5M���z�]ogRm<r����t�V>����v�'���W>^4�}�i�����R�F�?U�@��rm�x�˕/��L��*�u�7��}��Y����Ⱥ��Iź�;ǘ��uHN�Jf=���Ev�)_W��2�[,�k.�n]Z_s]����Z��0�W)�e�k�2|	V��3m��lǫ�����jE=������}V�5�߀��8��;�ˢ@�)�y.喡CM��ۖ���&9���L^���M�9�������9z��}�}cG^��(6b����k�#�j��)����7����5C�[[������3WC��Q�Wֹ��e M��b��"�f-��h+$���)N�GM�0�|:��ԒkM%>Q(t�V6:|�2m���[�����n�.Y�m�������4/���\�I�����X*���>N��'@F5~e�2<.�i{S�uل\d�9D2�qu��wm���^�
9x��W6ݥpӨ�,{w�Q��ߝ:�eJ�y��\���P�>΂H�#N9][�NKY�4�3y0�b���QI���v��$v��]I�"`ʸ��JV���b��U|�b�U<V��zk2ZF�hKE�Y\��vw�'+��S���J���U�ƝH�o(��Mm��Ԩ��;�$2S,����N���F."�6�M;�];�
���x+�M�H�ĥ����A�����4�Mi����̗����-�Ic/���`̽|���;z��R������o^��ˠx���v�*ª�
ǁ���FY����/bA����t��HڽM���Ѵ�ޯ��F��v�wi�ӵ�c���J���/v�@����=�WW:I
�J��ճ4疵�E���mf{�?Jz��? �̇v���N�u�_,�t�6�ʓ#1D0C�Wo�9we�&���W�eʁ�'�v]ޅ�E��8;	�[e����O*��c���4=oq<z���cQ��%||�~y��^u�;���o���2{czN�ݬ��j'fi��AU�y�E�>�P�4>�/z�W^����;�s*E@��
���xi3��	��Ѳn�����c��K ~�-77���e�z���k%���g��z���٨��ENM��������P��y&x�����	�(no�K��\�B�ۡ�8�W���s�<����=U5p��x&�+ƶ��MUm��;�VY<��/��Sҕ1�j��1���WQ�o��-����2\�8����;WH.o+NSOv�1G�cv��bU���m�4;4���ㆧ�
�`r�]b���GKa4/9f�R�w�LX��y�ʞ׌6���ȅf�"_�`�v^Fo���vv�ԭ�ɾ����jЀz���ڧ����O�y��ܘ���S6�,�x��p�=�G_f�o�iRh.�hG|-���^��k3��V��:�ⶻs*���%��1��[ܯ|u
���x��w�����ʽ�ps>+��_�I}w�y̶x]�2.V윱�-Y+�<����q-�+qyU�:����̴��kNأ���l�!�֚~�#z�R�?�ٰ>���Ro4j������F�:�^Xw�gv�.�r�w�È�Y����ƻ��Ҳr���Z�^��_�p��Q������������]`Ş������q�W��tr�K����fM�+��Ƶ%��F�g^�sb�s6�v�,ΪS��tp���������y�D%�,�s8�$K:&X]h����BZ���Hv)xu4��}��{�)b�*���Z��r!�	]e���p�
�Ć�I4bݟF�)�h^0y�5�o
�#�_x�L+�ϯ�qo��}{�a�q�!.�'�#��y�z�]I����F���,�ss	�)<V�}�;�
�����'txo��{c��{n`�e���*"u�c�wp�(%�w�V�G�N�Ѯ��yV�����J��w@X�|c�m���Vm4��F�N[vU!�=�^�C2X���̈�!č_�5�ya���gpgv-���9�k���A�ͽðڶ9[3���;= �>�|��jn�!a����lnJ�|כS���㹽#�r��(drF�B8�iF�vý��zړ_�$�gܩo��?�;Ih$7�8�T�.��7XY�¦�!\}��j�ɢ��|��J�5��}rZ�6��!�ul�mu��FPLe'�:t�$�5t̫ޙ� J�s6Jw\���]�����j��M�ĳ�b�m��3����H4:����qobW�U�Oeק�N��r�݆fK����I�Z�-�h��e;-��N(�v�0��]_���<�rD%26�ɴbZ8��+%k���s[��yzS�T���Ⱦ��-J|*-�i�.U��&���W^%�4B�"���ڎ�꫻�ۭ�v�Gb�8������ez96O�8Ky�8�ns��ԥ���CX�֐��wA���w��[ݪl7v�zˡ*��o'��X'����SV�(�q4�*�T��������\���5Ӕ���D:э�[��4��ff������ ܸ�2q-�z�x�2�7u��,���^5_gk�=W7)B.}z��e'���$�V�N��ǉV���^ uLf��ݤsq�א׆a�;����ǅ^��]�+�sA.��=	+;�R�ڿMJJO���K���ֶ����W�v67��rX���y�/��iu5��r�?:���1� ���e�,�)`͸(@7�3��bp��'Ӳr4�C��c�a�{9���DU��ɴ+��	8ڧӫS<���HN�-�; ���v�#)$>yf���뮣��j�p��Y��ܣ�GK�p�odUwr�jְ���]>��T섅�w�[��o41O�fz�d���X7wh�{�xۘ��Q�\wWI�r�6ɠ�{��an˹�f�S]]�C��Y|�6��z�?|8��; s�����SH/��w�ڂ���+�B��F��S�u�_X��لQ���wN65ŬG��'���{V��f_�=Y�BI��6u�*ʬ�̗�$o�#$�+�-����D���;�T#{&�X��\N��|o¦��j�p�XJ�����opѯa�W������w9���}#6�q�{�k2�Q/O<�}\�rjo�&��9�}�g�<�n�<
��V�d�s5?BUo���H���rz�D��U����z�d����Cc����sƎ*�^U}��P��䞸�I��x<�U�^��Sf��V
5��:&K�J֣����id���?~�\+���%�T3Əu[V ���4#�niz�o���z�iGL����ԍBN|��]BP�+���q��R{��)��e^���ZHpf�gV��N���p8�w��N��?(�L��7�ZoV���9��_@*Ux�e�i�y����Egs������ϐ�5Ê�Β6�M�f�+�KDf�~Z�ssm�����y��C>@t��ӗ�$�gYR`��3��f1���z;za��d��k��d�r�3^K�Y�!�O�q�ݤ�bm��n��A��YC�vH���w��� ���}��c�����y�ϕt�!^���{}==H�1gj��������ogim�`��g�7�H�vƨ�E⎺ ���wc��0�U���9H=ذ�W�-/�!OJT�G{S��)'u�����^����R�۱�]I%��g�����8�4�u��.iqx�5.{`��yv���ee��`3��_8J�
��FGq��l�P��e�mz[�����r6�p4a���W���,8"r��]�s�;�$8nP��{Ǒ�o[9�3�G8���/�hu�;������|��>�:�����������s����ٶ���l�m�7��l��F�o����<Y��<n����cts�f��n�E�07E���fY�Ͷ�`�u�v�v[`E�M����"��3���0"�-�#������f�nLX@`0 E�G]��,&��6�D`E�E�m��,,:��@6[6�&,#m�M���9��"`"�" ��"`"�"ٶ�E�\�h��f���,�#m�CD�G]���&�&�&�&�&�-��ammY�h�����e�=Y��}����2,ٙ��ҖW�s����~��>߆����������f���/�f��g�?w���Ǧ���_w��\�=����>��[1�m�?㿆��{�ٛo����m�6��?��oݞ4ά�|��o�����|��g��cl������?�/���.�C�l���޳��Y��������<�����ηl6��`�,@m���M0e�L�	��#b�� ���h��Y�f�$`b�m��Y��rm��68���5��ٳ���������ɿ�a��P�Ce�6P�ٳ���ο�����ݳgᜳ���������|o�~�>��~lm�n��3�~�?w���������ɞ���������lm�n�����������o��6�~vcl�>��[>}�~�1�fۿ�>ïTy�l�m�[8~��������\�=7�Y���0����=�3�xgy��m�_~�����lm�o�>���~?_�w�׬���Y�&�?V^~���f���#��vg�M�`��+6�mXڱ���b�m[f��
+6b�`��)�³0�0��+m����2�5c1[c�a[l��aCfaY��aX(͵3l1Y��l�j�
���͊ff+1�+l٫6�M�j�b�`�0���m��S6��b�1�l�fSl�j
lV³[5fճSmCSQ�6՛+�j�jٕ�+aLV��g^vl�e�~]l�Vߖ?V�����~�\��>[��|g�~���m߶yo���w�z�z66ͷ�����������Λ�g�y����o�|����~fm��~c��ngy��3m������?���6u�����'��PVI��vF�� E�W��@���y�d���[Wx�>��R�BUR�D�U(�BQ"�"�ي$�IRT��AR%T*Q!�yҽ�ke�VP�KYm�Y�[6����ʹV��Z��,fț���6�[f�]�E@<v�mi�jm�&�E*�Jm$*�MV�ڍ��Ҫ�m��l[SAU[`��T5���%_v9��ip>:�m��X�X�UJ�5��SwY\�Kju��*틫�\wu��i��L��CeYD*�8C��ε�մ��^@=QE 
/9�**����Ժ�7WR�EM5�[v�jd5B��Kc�Wkw:ن��f��L�o;�(��ͅ��\����E�g`ˢf�4���Z��c�k$��R�.;mU�%e.��^7KY�+f����J�lF�s0�T�U]u5��Y�kTӵ��snk[�N�B��5�m�D��=[M���)�\kv�;����t��ێ���nq�8�nk�n�ڶ�GJ�ٴ�YV���PyӖ��dj�n�����K���:�a�r��7;�uwN�R]��ۺ����Z��5��#����+ywB�u��i��h�v�֢�IŶ��i�먻b�Xb�i��s �ͭkf��٥�Z� �G��h���� np:�	�@\� �� ;0C�`�t�Ve�Y�6���� �4P�� .��Ӵ� 8��Q������t�@N��Mݜ a����5DK��cG�� =�p +������ �n��R�� �;�� n� 9��N�
��  � �~@e)R$M22b�4� OhaJRR �A��{LM%*� 4  b  �#D�J���  &i���"&�hi�D�=�2jJBR�@@    �?�G�/�g�9��廻WQ�"?�HA�E
�uj�j���DH��z��XF�I!"C��RX�!���$H^I��"$.o�?�u�9O�����'ʐ�#� (�i�/��(��W�'CU�)��J�����_���[�}�S���=H�D���2�XQ��E�w[����3�,Yj�\ܕ��0�m�ۅ���_�V��q��֣�1R[��������9�*���+2'�LQ��3%�f��-�A<xfḟ�]ٺ��j�6bUf%��7�8k��/y>0K�.]�dH������C�1;�5��]� ӅP�)�&M���8��f�.�-a%�wt#s�%�Y���LYl��t���t�md�������F�Yr��o�i!>��e8�϶+61���R=-]����H\�IɊ�^�Lb�r�n,�W�m�$��PKd�U6�ܪ�RPK��U,aR�/7h�P8�۳a+��l�X��p�Q#A���wgfѴ�E+Ɔ����A9�-��VX�ձ�j��(�+W"�9��);�v޺iYI&���S)}x�*�z�"��L����[�i���F�;�V��v��³W��%��Ua�!�@���2 ���[l�Hnc�N�I�5(�Y(#t��·)8sRt^�M(�9��B�m��h!���\d���07y�EZGs^�,A��++7�m�oa`�b��ZV�t�=�@NQR��Jy)���3 ����s��n%h��`U�بˡ����i�� jk���\I�AR, CbԒL�m�*���pP�Ԇ�{4�P����ÛN�W�m̉��#/`��i5�7E�҅�hU�ma��Ee���,����{ �F:a���-�;B��
�Z�7׵��Ų����&B��[e�#�T�Q���p�t-ꔃWs@rO,��U�F�)z!ڔ�<�x�bbج�P�;��d�pjl�m`����\BU�V%������4F���R���!+.
��	r3���Veވ�MSGdd�v�v�&�$��t��	j��8���BɏfB��$9��Y��6�B�7�-�腤����Օ�&u�3�(�N\,
Ȼĭc`) ��d�pZ;�2U��0蠅Xj-S\�\����V�5�e���]ۘ�#��Į��ҏ�Ơ7�r��;w�H�wRF�ID��.���s�p�%�-�0ÌR���B2�ٚd���{)���%�eʺ�E�U%��e:��i��ҘZ�.Vjl�D��n���KYZtfYV�M�,[
_�Um(��*�aQ�B�C�n�;���̓w�P[3#������]G��������WN�nY7e���ͽ�$n�TJ�*cv�A���&Y��cF�J�]��X�;�tUi�֭{v5J-�ZM�
�Ui\��7q\E�D�X5}6���d�wd���X�R�����w��ӊų�6�8�;hL&�)�n^@r�	�@���EX�mm+w�W�\Y�ZB���\x�ʸ�Eɕ���E��*�����VmiZ������� ��Cx�'4D�(ٓfe��x����Am�y�6�[1k$ ���z��ϱ��clf�j��m�zW��1��߅�J�bL#���Z+�D�eћ���f#�&B,EiM!�%�g�z��r��M4�˩�o2Sb��e�sj�`F�{"�p�&[�,ޡY�%;27%7�5�t�j�3jC2�	:���+��Y�6�
<ۉb��j��0�$�F֛n��r�4݄[s*�e��&��W+]����ۭ��q�۹��&�-��8&)m��sek�^l�*��tK�~#����urj��Q����5a��Dؕ�.���-�c��p��B�M��]�@w@��Ƃ����x7�@���E��;�ky�2�Jqv&�v�����=�C�"��{P��@Z����v�Vj��j�dae�2ƜL�)�rњl;�ww��rdf�7[S>�g@��GP�*����hB�ִ��b��%��ӡ�Z������el���@j�.:5����M0��k�
[q�N��^PF�M�u>s�4�{��lhDl
��	/	���wR����d�C{���o�(B������`k Wc6-��AJ)�G1��(�[�o^e�Եr���	`��}w��	�)��a��B򠕋P��
j�B��fQÊ�ך��"N���o]$�K-K�4,?3�ڲ2�
�����r�x%8��`�hn@���SMX�"���l��I�����4�];W0��e*�f�ܰ�`4��R��=�wcK���	d�Ej���p���YZrT�c"��a�LB��LZ�c������&B�V�g�`�[F��ՍįtZ�.Ǹ�IZ82�1d���F��K`md�7�a;�D�r��[�yF�q걆^�����W	t���T[�,R�`��pV��a)[�w��TPc�m�y���s5�]F��R�D�n��	���Z�7�dU�T�PVw&,#\sV�iB�˒�;��]�7�iU��-�tn��r��]An���nkʎ+6���Ccm5FŔjU֔�6�ɱ}*`(&�
����&�*�mn �������yO@�5����u� �f���:N���*;�τCH�>�-�p���
�UkC���7>5�WE���݂���ӣt��-��+�T�i��Ḽ Tܡ�Z�jة�dˍ����nE���ې;��N�f�����V+#�X&ub�]���0����j�DIJV��M��Bj�?	V�y����f}x��w�6W��0�&fc�>!�r�P�mSTCq^JW[�e$ݡE�X ˤ,1pc�k�z��,8䀻ڗH��+a�%Ƅ�PU��b��-��CknF�ۤ�62��M���kbz�sXm+,e�w^�T�r;csr��03�*1mHviV%ac�t�(U�l!{/ �me(au7A�RVA�	!Z��,H�E`<?
liR��VU�c�1,u�<�2��*�%�u�Ua%��.��u����)c*Y͘���
�QQ��	mG�.bBb;t���9DR�)*a��
ԺR�x4�*�Z槱�%X8��k�wLQ�B�Ԙj-˼�)�M`��^`�z�.���	��1�V1��D�V����q��K��n�y,Tج�R���.��F����"3�K�/2���^���dI{-JɰT���l�-L�KV��D�&�q%u�ɔe$� `*�^�d����U�EeIO�,],?:m��>Q���9��ͥ�r�E�e�èw[V����0r=7�"��&;wJ��Wb��ё��G�aI+V������U����C(�%M�'�v��ɦ�(����5�¬��1����Kic˟'q��Ь�4����;Bb�b;�����GF;m3.���6D��g2#���V%���a2-��Fú�����V��:`V
���5�ZY.���О�t����ea��&�Z�kf��,���,`-)���`Eq]�f�UԦ��Ht�ei����2��bb&n!U�����q��J�6�@�SL���$��(re$�wNjf��$�&`��	�n����j���a#6�0�vt��勍'ayq�ʬ�x�ʬ��/�A�"n����n�o5�3J(E�[���]���VM��:��x)��(bN*QJ�94
���"�dն�Tư�q軲����J��-X��`K��7A �`���7P�Ik4t�T�f��ofmb��S���x1=��Uc�j!���Fs"���B�*��&������Iа�qڥ��rcͱk.�<;q�'�N *H2n4p;�1)��5�ARj���=4��vuݵ%��P�5AnB�'�(��c]JR婙W�nL[*M��b��.����]]�U��R��4�gA�g Y��45���vL��c�'Υ�N�FF��p|�� �&�%Jq�X3X�vD�����j�\Y�І�+�I�dѠ�T�A��L9-6��M	WJ*m�P���� ���(mM̎õ㢎����H١#ϲ�Ę�R�O7
�bKN�7l=��cv�&չ�j �b��k6����Cl���$k�W�^��jJ����\v�`�{F��ka�q�̱LD�hÂ����6ȝ�i��Y���̠1��U�g ɥ�{���
]����Q��;V�6�����,e��Lpa{zK�E!l�`Cw����2"�f���������n�6wM��O+jJ264�)��r$��r=���pCe#�n�J`�l�qm�e{3p*/nefEu�Ʃ�F&,�D���R�N��l�
���ڋD�k�1��w�F!��%�/R��f�E��ō��%WS-� ��E=�0��d̂�Pz㨀j��X�S��fV��[R��z���7#y�+L �
:���n��^Vw���fο5�OsЦx,��٦�u�+������Q��#?�5x�J�p�Sצ���C�;������J(�WZs�:��u��]4�9���/��{ٹ-�����\u$8m�<��%�������B(�9��g�YHg.�K%�؉�]j����k�&�k�G�;���+��H%�V�h�4���t�Uv] ���W��ш#/ٽ�+�Uy@�)��p�)�S�*��ԙ�Lv�.��TuH�r��&�٨��k���v�V鼷a��`��U�ɽ�g^U��z���u�@ޙ([�設�Pr��ج��t^�3���*��B��r�Թm��P�6��(��Ol:�Zs$��|Y쾩�v-�B�R�P��'�B�\w��ҝ.e��J�H:4j#�t���;�aM��ͮ��T�%n�i�����hR�Y��IP�ߴ�Ĩ��:��ƅ9B�4��Vj7�����L$�}Y��-�tSyn.��r���G6�c92��M5��^�,bΏM7��7�0�6[=��P���c
E�Eu���J��b��\���ch��#.@�=�\}�f��z/4���=�d,�xc)ŵ���B�^uu® y	��؍��܅Nu�u�i���*R��������D��]C~w�0��W�܉����8�	K՚
/F�y�ũ3V���[���-���[}���"]NFÔDK�����<U�W�:�6k0vk�J}h��<ro�}l��ky=�1b�PQ7o�*�.ڏ]���j_nzjT�
� KޜLi\oaj9��1��y3��:F'm��t��M�?���k���|��ݖ�RE$����/���Žͬ�S����ڷ�f������Q�Hu]��O\����+ۉL�[��b�d��աrک��O�BX�[4���n�^QN������[�<wU��VgU�����:���L�t�^m��4�F"�����=�甀��Wj�	C
p!���F$���b�3��u굕���@Vn��
&Ww[+.�,���n, �6��eccKZi]r �bgcps�Q�� �w�*褼�ܹ51Z��Ĵ�1e���n������V(4��{��KԨtӱtFZ�σι�z�#�r,�MM)���:�����"����i�]�<:+�Jn_By�" �9�}��]�\Е�	��7i�[7���z2D���DC�
����s[;�pd޸tԑ�i��b��#L1�Ͷ�!�5��\��t\�z��y$�&S��ŕ��`|�1�����ΛLbʮ�����2(�4�'\���٬�rP����3r��sC;f����^�88��ZW[@^_x�߄��Y!.F�un�(�������]�s��3�db΍f[�`<�L� ��+UΔ�����s���u���O4�X��v��4mr�Q��Y�E��"Ӿ�]��fZ�2��wE���U���9:���XR���r$�Y�qܼ��a"�;��)^c�H�$T��'ڪ�d�v�c:ɩ��Y���i��37�<DU��쉶ᗿ���Eh�K��=��P�:V��I,�*�ob���C
DP���N���{�j�"�H�Vm1AN��^����D��B��]���ҊN��{�UM�ΠÔ���(�ݗG�.L�[�]!�.��M�w����^�Wk��T�72p�^���ڤ��m��^ŷg�
�B�
��E�U�8��4�;�Wc��� �$��%����b%u(���֬�'j��!�{A�%���R�\���vltD��"�����[O��[gCu1db��K�M��`�2�ܫfJ3�Oq%��#�k���nj��R�S�A��f;�S�|z�g<��Y+uRƻ��F��3�C6��˵�WR�tњ��/E��PaHK��t�;��-'f��P]�!\5sx�g5�\=�kp���)�wh�L[�d����7�.0� �X���lٯ��#�%���V�k%e�Rl��d��j}��9k侂X�f�J�f`d�G7��b�gbϒ�¼�Wt��g3R�v�P��vk�;̌�֯���U�%*-�r�h�O�b� ,;�>�G�����3
ڸ^�L�Bŵ�q+�Ӻ�|��+-ʿMy�	5�Ib��͆�R󏓮n�oV����\T˜��)v��b��2������U�M�e����FX�M�c{t��E<cqR�
�i�{@ZfRm[�BxnD�:
f�f��.�����Fp�Ǽf�]t��J"��Õq7:�K�����N�,���&e��|Z%�5P.��h�öD��d���gf�Œ.7B����1�K�G/�7�
Z�Ye���ޫa��۠ѝe�R-�	n��e�� ��`�J��&e�ˡΦG9��7H�f�E��PTNJ䵧Dq*�B:��J9Ň���\�z
�Z�}�QRY��&S��\*��-E�oQz�0���5��%�ҹu<a|2[�U�E�s/v�qT��EҔЙ�ʲ���r�9��'^L�8b�>[4&��W&E�B�����*T��gP�n����K.�� ��?uF�p���p]��X��7����<��V>픎兔Ҷ��g_uHl��a(��/m5+f��%d�o�U���pHl��'��]�h&J������teL��*��$��aunQ�DI�(ۉ(����u(1Y��U�u��h��U>�4��<��^���
���xi�u��m����SͲ>�Sn+�@��d�ʊ�4ZÏ
9�Nk;(c���b6x�pX%�qm�`�F�;P������Z,�f;����ڑV�j]t�(������,�	��TM_�ϵ�	^ID�V@����D���dU�98[��Δ��:�%����CX*�ހUj�������md��-�c0t̫��C���]��J�	�7ZH,;P*p�]iA�]bu��}�=�T!�enu3sSb'�o�	ԫ5��j�ծ�v�{iȎ�ʼ���<�dt3Jw�Y�X��:����S4&����v�X.�D��g��.��ê]f����e3l���d�Ro������Sv�g�,��`>V:ZƬI>�-�*ؚʉ<���o�+� �J���v��zi�������%�� 
�s��>����g�N��5�Xr�� �1���eꅄ.�]�°��0)��CS6��sj-١�v�	�sxIK�k�*���2D�c�j��ę֯���r�N�fn��&h)�m��X�@ս�G�2�<��-��0�A$9����9VNt4����Q���Z��>HVr1�GV��������f���@��in�70q�5�5����B���}V7�w0d/R��Q��4�P�}��u7m�&�R�8k��K�w�&h' ZU������P�N�|���_Y]V&�XW�Wf��_$�e�i��٪��ۙ)S�c�F(�	�fo�s���>��<7��\��%K����-��*$E��1h�־WE³y�B�a5�]���PJyA|P�F��k̂+�OY7��˔�{L�\�1�L�ے��S-=6����ѕ3��83�l3%b�P[�����t4V�;`k��.�R�[F��ad9(��H�:�����X$ǗS��[B��� ��)C�ޤ@�݂.�ڷ� �h=՝��e�<�cG��wC��5кw9o�;�]3���6�V%�Yb�S�x��͜m�.K9�$7��0o/�C�p�|�V�9^
6���̬��pd7����N�3��릭��R�\l*���YO��ԇ�zM��%�5f�����'SW��-�FnB�m���c���G��H��st/5�2�M���֞Ҙ���B��C�M��Le������N��� ��vb�ʱ]�!ͥ�\s>nn]2�[�1S��n!�&.3E\p�<�A�m���tn���}��VM���Z~�J�'��U�O�@U:L��t��.A���S+��v�h�~3�@�رfB�=�D�#l��UC�U�#�k1|�U��Ae�WbZ��#4�	'��8�Y�J]����&�<����x��Z*�����ҩ���k"*B�-mQ�Q9�-��8=�m�B8���/��-�Ņ׈^M[�����t�:�A���(�k�����KBhp`P�S ޶���sQ]Vi}m���'����a�c"8��A$i�H��U��t�{�$,�UA����ܮEc�s�z�ǲ��<��l�*�uҭ�ѝ*��
rI$�I$�I$�I$�I$�I&�M�"��cq��NI$�I$�I#��i��0�IKad��S݆��`�h�}�jD�|�����i�FG�:���@���8�rN^-Kb�O�l��G�S�[-9n��iͫ��Z�o�	$Bx����Wsi�8�rI���Gl���K���M�e-���߳,���m��ef[����5��5}�B����tgZ��I2
�!K�®�k����v��v��u�f�fR�[Ԫ�SP�W{�eۂ�K-�{Ge�0]00�ٖ%���9
}g�=���0Ҽzdy.�J�K��6�F����;��\�����,Ö��ݻ���P�r�S�W�� ��5+�*�R&�p�w,��b��リ,ud=y�fZ��k�V���q�i�k+:�
N��`�cwa[V��8GS��V+U��Ts�;h�W�+�Ϋ��lK���;��t*f��as�s%���s�_|ˎ��c5˴g,�.dyCb�/,��:�B�H+�32-Yq�atV��-����剂���B�+��5b��P�E�y�H����E���������+�f���A!��=���n��B8�(����֨�Aen����kr�Q����r� ��K?\<"���f'�ԭ�QGod[I�	0@���Wh�F1�Yo�땆��KЖ�n�i�iS����ͱ�,�[n�A�κ�Nq
ր�k0v�	�VSw�q�����װ0��һt���r�ں%�7�{p5Gc�TҟI�8Dد��e��9N!�@�2���q�d�
��b0��Cd�Ae��>7ck�@1]��93r7�I�Uj�ۺ�
�9��t�P���V���jK�N�������uC_9��Y}�|�э*�	���z�җ��T�U2��x����KS)[T(aw()up7%UA�ڟ=��WKo��tF�57�]lu�:*
F�&B��b��sn�{���u�Mf>�i.fd�yT,�W6Q�26n�Z_h�g��bm�Q�^��%���-�B�u�٦H�9�����KFS�|]֮W��cb8�Fe�k벦+�]���S�͗2��6��J�c0��ҫ�l�H*^�f"�Գ9��w�+Yq��w�QF���5��������[`��9�̧B�GoG�j�9#Ob	��ޖ��xե��Ku�@w.���5P�1B���f��l]��i����Q�I�V_pi3g%�6F�ӖɈ=C���)R���F�w-�wf�A��\�s�\!��K�CY�E�c	�>�o�&f�:n�����hrW�]
����Bnb\�iA��2gI��VY�J�.��*� ���z�8�`�:O]�"����i�v;jj�շβe^�\]r�����>�Xp�F�څob�k��N���Zy�r�ћ-g1��d	zw��!
�]n�c�5��K�b2_AGX��tY�H���@��`��|��#F���f<
�F�I�'l�A�DA��e�Y@`��($��f�S�����dm
��\���ݥ�o1�V�q�Z���-vWP���d���j��!�0�@��G׀�&9g�"�<4[��s�1.9q�^g}wLu���A<��j��g ��§-��t��,�vT����%�
-��4���30��yA5"�U�R��1��T�
��EX�z9Q�ds��@��7:�O���	����3T�[̶����+�G5�co{����I�S-�l����%2��@��?�k�oPU7x���b�QS50����3/�waK�B�R�`;�W6m��W��G�
��z5�6xpcV��[�.Ѭ<9�p0/x�9�mw;γz֧F�KØլH��9B�Fأ���
W+:�[��3�a���r͓b^,�e�]Z�*�'$P��hf��7�C���Mҩ��� �)VVl6P_e��*�r��j�
}S-�PW�Y���U��.�²�T���JW6��w�`t��
^p��M5tN`/0�9ODY��k��gD�m�eڦ]C��[�fq\���$��J������� ��/B�Zi�w��wq�PK������F�J ��h�M�ð��5��$�9p��@F]rG�
�Gn� ��w���+������������%GC�Ùd$��h��y�"��_+�e�VP�H�S�{e���T�Q*\s�_�}�Gë��;�+j�Z�*�Jє�/4dv�'B����I����E!G��N�yui��B<Lj�.���[��m�nr�;���_bX,N4���N�O�31�5��DyWVY�(�r,�ZwQT�\�ҫY�5W�o�h������Z���u����cpUoO�`�Th��wYr&�N��]]��	fՍ_^B�:��Ɗ5H��F���#VMaJ%��d
\L-��-�׳�10Y�(;Oy�L�%���ʞ���F΁�v���h�0]��]�w"����bʒ5�1\>A��<�!v)`:���@��\M��I��Ps�;�����qGo�����v��w���ӛа���0j<ͯ�.n�"������H-�6ɻl'�.�ZV.Т�b�Ei6��5��ol�8��X1�1�0�ϰ�s�A���n]c�ЭI���)Z�)�	ܞiB���!]ƴ��ھ]���W�wb� �\��o/�%]���K�J_9�ЇgD(]�j����ѕ���bs�{\d�1V��7�[#���U`�st�#6�meroU�Ovqټ��gѩ��q�۱��;0k[��Ӎ���w:6�T5���b�K���B��Bo�o���B��ӷ)�ќ~�y�[�1m�@�x�M��Z�� �=x���3� `[���}P=�]jb�w �ZlK�	��u���4���[����5�T��br͌W�)��=����lj�uy�ujY�gY"�`�q�SZI�R۫����9's*�g[�T�� �48(\?(���wa[n��D�+�
�P��cU��C��ger� �ą�(.�I*��4_r�5�L1f�q���BJ����R;CI��W{�񻺔Jʓ���@�}�*qJ��]�C#t�u��AЧx���Gs��)fl�#��郯TER����Y[�� 4,U���2�ɮ7  %HjsIwa��+L}�f�w�]��?Y�!�����G�p�.�\_T�ji4��n�m�,3�ʭ�S��g�	�)�:R�(Ô-R����z�8:<�	�f����#��H�3jl��a.���y�B�%��sYW-`��
4�5����8`h����9}{�>���6�ނu]�
*��<�9��m:)��/_,�Q�ab��{qJ�#�F��n��T@K�w:Z�V#��u�$z�a5�v�T]�0VG8-C�f;@1��ʔ���۰ ��s5d��J�Ѥ�Nk�e�A*�{�`e۠�g+1q���H�M���u(�i��v�h���p#��j�<�{�%N�,�;�z��ޫ�RM��oz9ʯl,b� 2\N��5����i k�)l�V�GAl��tP�AaJX�N��H�o�yc.%'q[ί�������l�bG&9���]�g�޺���!��S�m�I+9>�:�#y;+ ��$a�ƅT�m'd�V��&�G&�"n|n��eZ�mm�wD�oU�k(v�j�E��5�c�ނ�h�n���&1��]օoX���0��̶���\�k (>��aV�IIg:O��`7��@acU��F�b�RU��I�ġ	��=�hT�Wɋ�%wb���A]�ͷ{2J��5�t�KU��F#��ʽf,��s��b��u�f�:%Gb�,F:�oY������+F�v�m�n
�#7`qH �͍[�������@G(9�+]J�s��D�Ea`�`J4�$�oHo��èÛrQlb��/k3+����* L2�ηO
���^�`�PILrU�Ҷ���&7 �A⾎ʻ"U�j`���9�[�M�\�OV-֒�+z�����fӚ�xqvH�\��LFu���e��0"4��*�B��ʸ����mtZw��]O2�:݈��9�D����P�-�D+�Lg;�$�W�0�1T��0��ҡ2�.n�G���8��Y/��@vdzu�bl̼{R�,"���.�UЛ��C?J�{^f��M>��+�@�e8�%��M) ̡l"ik����
��!�	��7�H�أÔ��U�o�q�Q�(l��u���;T/o6D1��d��C=g�G��@[.Z��WY��RNfV��9����������zV��u�r��㡑n*�N��ʕ����
*Ľ���Zr���	*aíK�y$�K[wg��%�/17�t\�JBGD�v�orʽ�y����Kx|V	��3z��$۬�V�����9��m�D@�;԰���'�ri6u�w���9�
�Eg8��2���"m�WQq�;����ħ�Y6�	���5n%/i�����Z�,SB��n�nʾ�VF��.�_Ͼ����QB����\���	O���@�?՛�{6ڽ�v�t��;]�>���4��,}.��c�۫��G�Y���}-m�u+I�i���'>����B�L�"��'��dS�����[\u�[��n�>ƕ�1�h�(�()����v)�Fæ��}�,jUj�sAֳl�n��%Y�_ݒ���^6��a3�f�����]e*V�{]�jYq��Sʖ'f�F�8��o�t&	��i��>�Ip�:��[��J_px��#��R��S��X�C�f���h�m%q{�6�mBB
��Ϥy��(G�7v�PX����XYB�)��aP{���I�c���������ֆ����_���u*
����k��c�) E�7��\�C7�#�,)O�um]���G�.���<���kqh^]z^Ū�A�����8���Q� ##")�_;�~���Nढ���iB��)R�"JB��)� 8Iʔ)B��(JC�i
iZh
��=�����(i���`N�'rbV��)iH�J��Q����
�"R4��)�.�%)hJi����J����j����J�4�CB�QICuuuu��+��Z�z�Dd�� OP��zx���mU�zp�&�U��zo�K7BQ�^���䓙U�Ep,hf���j��!P#D*1�t#�w]������6H~��/H��"aF0D��u@$��u�ڑ��q���B 0�}t�Z���0�&���?^�/뙺+*~H��E󘔦# !:{M��3����q�������}��2�OR�bш0�E5#cP����F�}Z]��\Xzc��GC��Z��?��j��~`�\���v�w�fe->#�6+]�a� _�:�Yk�i�	`��+`��0�8�"U��~$A��1W��
�E5U|�ŲgW+��Z���-���,h�8h=�Mr��yTn���D��;�<Q.�p`Zr��eKUz~v�
,We% Mk$A�w(�����J"AH�F�}������7F{iӼE����X�d��,K�
F�r�U�Kr�[����6v`է*:�DaQ"�vE&5�e���7��J���Z�C-9��-V��D�9 c]ݩ��1��/;1@�U�)i�|�\.����@�[�O3J��#3;~8@��$(n���ׇY��V���<�ڹd�-�+KS� ����_�[���L���B�Z�iUd�_��s��v�1�=J|(�F��rb�� �B��j�����R|����#>n@چ����8O��>@�����"w}:Dnz�P�O!x}��IB[�4q1q�0cp�	����ڼ�jl�����d��ATSs��?*�Wn�Y7Q����vv1�>Y0�iY�S`�O�<,!��4�	>`X����lϽ[֨����MSǼKŠ
>5��~H�3��۔	\�vߡ�5A!_@�#w�r�b0t�Ֆ�+7F��t蜎���+pu�$Cp(�W&	7��:tY�
[��|�i��4�D�ڰ�y����Y �� E��YQ�zN#l�%4ۆ^移��Wg��ꢫc��ób&	����m}7���s\o�ꗮ���C����V�>5W]7[�\m>nR5��u1�E��^[2'��0s:8/��U9�'F��_�'%���޿��	�X��J������1�8Z8,B<�.�igqV�sy�1N�Q5W���
�狳�����Y/_�����G�������KV�l����!������R<�d����Z�Қ
\�r�A\F�AT)�0K0u�h����-j�C��T�q!�=<��@OO#!9��:og�-�H�j|�ﮩ��μ�9
߂��������a��vm��f,
t,�]mm�4�����J�'ͩg��:�D�j�j�uH��&��b���p���OgI
|y��C�!�[W��QJ��/3�H��q��Β���˺#�5x]�1U��'��8������ ��{��2��	��1B(h���#�DS�j�n���h��\H��@�g:��n_:�V(�U�jJn�7-�6d���ꨚ���?*� GphH�><5dP��f�n5��SQ�_ܠ��T'.8���Z��}�����w�l&`�r�i��W.
�r� �� �B�%��i��������r-���� O�xV�'���N�3%���5!Yԕo�ɿ�?E�
n�Ҫ�_k�U��_�O�W�G�w����%�c�e=�R��1��,�g�X������05��~� .����F"Fi�	�.��aڮ赧��WX�h�N�g��R��*9�ݺ\�h��tٴ.�.m��c� ��) ���u9�N]Ι"U���y]J�V�7��E!�������=��J�囯Y�{7M�@���Tt��o����;�JB���h�,T��t��ǅG���t`�>�83u��m[�t2n�s?v�^S#��6��6�D�dJ)ɻ��7�G����N�B�4a�/�Z�&���Qn�����:�n�sR��Y{��U�����j	��0gr��Bs�c�K*��f{��Q[�kvr�u���s��o"?]��Q ���x��LvvfV��{�qs�%�6�ƀ9��� Q�lA��*��-���=�7:{�R&�W� 3�����c~� !:{HI���t,S�\ڎ#���,�pÁ��hc����0��I���m�"Â��D�%!��c���ۙv�H>��ʘn,��U��G�P%(�(�y�R��f�ɲ<:��V�7��b�Տ ]����m 1��1�CQ{� ź�w���D��V��.l䕷���-�ܭ���!w���k�l: �:�Tr &�+^��U[�m��*8!���1Xb��N��t�î���+1�j��ޝ�ת
w��X��ؠn]T+�P��-��.Zy;Q��2'��b3Lel�"�M �"�v% ڵ�_�Ξ����iѡ�iWq�eZ�C���Zs��㖫E^�#�WT �h��M��
N�$F�4k,`��E���vX4�Π<�{�2��+V�l�������̈�-�aY��m;P>�J���k�j���41������h?U�V���$2������Aħ����nx���e	�y҂;1 ���
-��:+{+��:U7s �#9HP�D�#@n4U֐�ڕm�1U�*ռv�yxuۈli�j��ݪ�_B��М �ŵ����:��û��
qG:��̖P%΁������y�F������}��ܕ��*#�á��k)TX��|~�H��|@���B��J�;����S^[SD�e�\��4��:~��q��T�����/Ȥ�:�pD]�S{>,u�K5���%��@Q2"p-���?8�$:���,�3���+�S'  �������Z�TP`Qq �0gC�B�s5��BxU/6��a�~�J��Rã�Sʊ�uҪ�ób� m�{4��^V�������jD�쨇���Uz�/�p��8W�������`�Ur�4pE���)h�n�
|��;�f���8�s�u�Y���l���'�?ec�)�$���vjMg���+E�<"x�W��8{&Z�Z�V�B)� D[?h:@أ�j��4c�7�H�c�nU�Z��j��Z�,)�w2IF���z!����(�k�y���p��G��[E��9,�Y��\��1o�׏ ��T��́��N�!�Q�oS�Z����z�����s�e���ui^;�n�N���P��������m�MŽ���T~�E����Q1˕d�\�	�PH�&&1�=]M����𘫘��"�!ÑQu("yB4t1��	F+�w��|#x����B*Hȁzbrv����L+���_(�Z���Z\�ʐ �ʊ�r���2���V��(	�s�K�K����?���?t��Θ�Ć�g��b�6a���!�Zru�\�R������l��8[���1�(A���"sUf�w+Gp���3P:b|���4a1�	kML
�o���K�&�dQ-���� kM5K9hxt�CD�L���X����y.���	��K�7�"*4�4\'6`� (��J���~�e	۹�!d=�Vn;��y^��t Z3�1�tEJ�y�Ӏ�"{;%:�e�6��+��m:;��I����uיX��w�Zj=q�C����e�x)a�C�R��ٍ:�!�bcDH����`�S6�����DME�C��V5Ɋ�0ԩ�ٵ�"���Ł�xi�Ŝ�EhϪf1��?�5��˼[��/���b��ܻ�he7�TD�"�-�*�i�����m��Z���]X�^��`xV��
�@O%^��;�=,�,ׅ!��փ�r�N�:uf������ۻEƅ*󷴖���Ȓ{LTj��^S#��6�
�G*�+�J9�v�+_��#�O�% �48.s�����P�nf�Kc�ƻ�"4,4HOA�ܘb��c�O̡����fsV2���1�`nb�IO��Q��!F�G4�c	��6�x�׶�n.��Y���	cU���v�g�[붑������;���$�"��Cȭ ��u�%��p�s��V3�n�2D�>lެ�U5|�+.N��m���� �ڐ�w��h�hp �L���|~�Z�ɳ8�.��\���t���]3���e��c�)��0���e]b�]���z�}�1~�LX�^(��9T�B#��ȟ�Jzr�
�_$X0�h�S+h�KC��i�am��a8�S8�7���:m�}'�q�Z�h����" S���q��zoXL���\|)Wj�Th���$A���S���1׼��sf�ة�o���9V��.��_o,��F����B�u	H:�{9�f!�E.��k!��=?4@0�lW�S�˦��1}S�ܕ�OYvPbɅ�������BqUƮ�h�����۾��].@YqUL0G,艆P�����p~�G�?A �����%�=���r0�a];9�����CX��cI㫬u�h��t�jZ;υD���#�v֛�W�<=m��7K����N�b�޹W��¬#0���j�#�;�r�Qw�dѴ�gMچ�$�5ܢZ� ����?�mQrx,�+��y����
�U���x�U�~
����V��5:�����_+->W$��^Cxu`��IC �.��So�pYs�'^
���$؁�3�(_Ͳj!����2S��DZ���/�hNț/Vճ\�rtԐop�n��*EB��fVh>��ߕ��r�)�u3����6C�1f'����*��ܶ��Ǻ��m��ʠ�c4>laV�m�9�9Ϥ�1�6
F)=U��(�:�Vv�9y��'W%�г{y�C�}ݵ��Rpd�Qz��벹����>!_e!�o=Z�яB����mM��+����E��`�D�E�e�d���	C)��j��M\��ނ$z?ű|f��Ǿ���
RJ�F�
���hӗp��mݙ�g�����Zj�,)���V�{N��&��Ӥ���3�lӡN"Y��X���Dc�l3{JV���A;�es�:��nu�A=��qTu[U�|��o��'%���u�kOC.{!n�����-
��+��zS������o^W�M����k����	*�r�x.5�ՓMZf�Y\�YDYh�P�Ep��Ŷ��1)�W�X}�\�y�]]�����7/H3�u�N*�֠F`��7fւ�)#�Ou��93��f�Ԕk0�s^5�R��;�sF�M,�
�	2���s�	�ܴ�e�X>���y��OC�SB��s���A
D�H��
�PUj�WF�)7����-��|�n�5j���̻ݝ�b�W2	�e)N}��h�6Իz�٪e�u��Cf��'���	%d)�)7 ���9Ljn&swL��yG(�̤�¿T�=�Uz���(hD�Or���
hR���){�R�)M	H�%4R�"U"�hZ��R��@LACHPJ�T4�CB�w!�B�Q�B���M�h��ЁE �������yz��翱|�t{��q�;�j��r[1%�z�,13>}����%?$�����%Q���!�{�C���������PF�����? ���:��&��8B_2{����%�4{����>��y�7�����w�ן���>A�:��·�{�sy!�J}����w	O���rB�lU!C�>G.�d9u!���?GP#C���s�O���C�HLn�ޟZ�w�����C�
1"D@���~ߣ�|�G/���w	O�u]w��u�4��'/�r������f�B_���B�^��xB8}�4�}��:�_>�z4}���B�s!���'�޸�BU/��������䜓@}�.�>�g���)z>�:��!+�z��䘈�A�z��;�f�/o��>#�_�4u�B�������<6^BWp{�9	O�<=c��{�BWݐ�}�g��u�CC��@h�G�����DD�� �5����^{��"$�4�����A�}��(q�0~�O%��`(;�Tɡ��K�9��!/^�t�����JK�� ��9��� G�#%dz�gVy{ʽ	ZC^KF��4�Xy? �<��`�%P���!�	_o0u	A�X>GP��]A�Y�)>ɿm~����G�䜹�!�<���_�}�{�w�������F����u=K�/�x'*B�S�s	��{�����!)�ۗ�	T�������'�9' �������g�箺�]u��~����J�����߬�	\����@w9����=I�@j���rpkԆ��BWQ�O#�J}Ͽ0u�/s��z�搜�S���ް�}���=��}`�`��/�4�?�䇻BU�4{����A��N�)}]G �:z�|�r!�s/!�� ����O_p+�B�
#�dn�NJ}Α[ѻ�"�!�fX8�����w�����!���=I/�jr;�1��78]��g:ov�.̜�Q]����Yܼs�W';%��.���9̴�}��"#�bt�G(G�c�O��J����w	Z����>F�!Op{�A��BR��pi
���P�B>y���^�˯�?{��?�!׸�u�<��������|���̯���+�|�=ry�O�� �/��N����~�x~�D�wڑ?du�N��9�,hʙ�^U�Z<4C�1x�Z��M�X�j�H\5r� |���s��^ܫqk��}t������㢛��(��o��@h���CA�r�ҬR�Od�nQ�B�����
t�(( .(�4�@8jMf��}H}bſ�X���*bѰ�Dq�j�P�3��>V"�`#խ��{��WNU��:�p!Pj򰨛��<O�Z�Edt�ڦ��R�q g�&�W��_r�i��?���d��Br�is|�p�A���p2���rS �[�++��a۴� �G6��!.��+�z�	��婽�j����sDL�
��ע�ua!lf���������.>��]�!yc_'&�t��*V|�}x�ḱ>
�e/M�yb�󎂝^�2�sd����m��?z\W��A��]IX��,�]lV���)�}��V��~>�P9H䨥�gvX��u��)�)��{���{;>�f�G�K��#�3�'��rLG�s���;C:X�G�S��jb�'[�ŗ��L��Ń�5l��(V?B����̕���.+��+"�R���ʭ��~�1�۔�"xՄ����zu�W��x�����,5�����K�ag�����{�R���1?εNs�ݛ������.`��X����yp�<7VȓíF��K�hKv���W���	�z����3���uƟk(v���2띮��X�r�X��*q�҉�O�_}��ȯOeoE֏���U����w��������G<z����� ��k5�uc	�ܻU˶w�Zm�V2�]&��{>u�v�,���y�A�:�����.J>��������x9bˇ��7���v�\#�3	ƺ��Pc4^� �K�?�{w_��m��)���Ӥ&ޢR�R&�n�g�]�dgc!ɶ�uMMZ�f-�-�r�		G�)�L�m]R;b��i�������yG�/ڜ�G���s�ǷڪR5J<���(����*�-�{�n�U�ן��ݸ�x��u\�3~��yb�	^�	��%3��r�i}�U+,YW���˥*:�u\u��8A���zLoٓٓ�)�Sb����&��2�eӶ�u�.�{aoo�r�����}�ԒS�O0���y����>�;�j����{��d���q/��(��vj*��Ayns֘1H��f/gP�K5<�1��޵7اw%M��6��v��~� 5^^5��z�Z�7kվ\���71�[t�w�fG��k�5�{�ע���k�˗(Dwp���bY��y�˕l�q�a:��RQ1˖�eD�5�'��Yϗj�2a>w]���;��g<5�{s7�~��x+{�*F�M�����&4Sٺ���@T�e�r�u�c�AOͿ��an?E%�ww��*����\�si(��pͅZ�2���ى9���,*���T�Ϧb��Q{j:��:����5s�[��ѹ7gVƩ�k���<3Kɝ���_W�QǤ�=3��i��ʛ3x�3`��K����i	��p����6r����KLe�h:E�E?{�+�1L5Ҽ"��`�k�ԅ|�DKv��~�癮�'Zr�A�nQ�~0������'3�����p���>�<K���b�T���5VqU�`���f���҂���~K=�m!Y:�/����F�5��g���'Y��M2w�j��t�Ŋ����뢻4�ST�9=�/���7*ۻϭ*��J�p=S�L/�E���>�&+j\�\�|!)	
�A�_L5�$�v�.[������o�[�#z�U��P��U����P�7�qJWf�����c/�y��8Ō��e	�9��.�!6VE�h��X*^�1��(�Ii�>��������/:���U����қ�IjsawM>תc�]�!�«�g�Tt��͔�2�uh2{=Z�058��1:�Q�����=���.H��^��t���h��ܱBz��)=��C�!�c�]A��1{�z�WOԠ�����5��#8��J��ʶ)��N���;4T���W2��}�Ѫ�%])�&��޿G�}Lz�<���!���9HJ*
R���^WK8�2���X�5��a�Ɯ���5��~�E���w�orZlS�쥓^)�`x�څ�\�����u�Ce����r�]�H*Gr�mކe�FXf�.�c���U���J��?W�,�5ƣ��8�6
�JM���D�겸��n�=�i9���>�����1�������n��G��ۭ���i���)��<W?ux�j.��������:��i�R�Fl�|�Jj9�(�ax�躏cT���X�-:xv�)�J��V���G"v�+�=H�~2D�1��U���)�z)��5p���sv������ ����vy��R�
�����sR�p ��1A��?f:Aۗʥts��'��^n��n�;�_�(�l�!u�;{V��5�bo4>Y7����Ӎz�+�w(��[1tI��9ޚ��v��x�i
[hu��
z.1�"�m�FVV�)hc��0�h��r���n���f�,lT�Æ-ˣ��3�涺Kw�%s�����u�Kh�&�%���Md�u���U_U}T��W�����.<���ܮ^���x��W*;�-s	gV#�?|�,�;���!M>��moڽ��K�n�dl���)��^T9���e{�����̸�v�{�u)��[���Q��VPO�mi�':����o�qR��x��`�������P�����^>��3�19.(Co�����D�r�;N��}R��ߏnWT���jg�ޗ7/���|�����s�=������g��GЭ�\Λ^��w��^�Q�IK?_ZX �ϲ?M�J֔+��o�c��W�D㓮�����S2�*��1�%o�N����*�߲.�F�R�[&X�p�F�xq���t�i����e��:�K��)�%evG�R�S�7�[����IBy铥B�ﾯ����^\ק���{���q8��Jq®�g��d���~�r�P��K/�r��b�)Um�+z�6ԭcn~P �֪����x�4�z�����������ΐm**]b��ں������r�=4���f>,%���ۋ�Y��xT	�s���n�����x2�/^��!�%�N8ؒ��]-tGm���e(���DQ�.4`N����,SDXә^� N�(������G�k��)Y][軰�r�~��.!�;�4���P�W��|�;��>��3�WJ9e�7���iO$��ݨ��.�i��+�Mc�(���>�?t����2�Q�H̗w9`�bK����Jɒ�Ӆ���2m,���ZF�DJ �$�= ���H�����6�M�/��O&*���S] t�kބлU�K+�6D�Yktݾ�=�ri���Ć5s[[*Ct�[�������{��W�$�]�Ԭ���Zb� ���N=)��r9�Si�(�]ۚr֗�G�Q�N��%$j��8�/y����ג����� @ݎ�����滭\��Q�8^��̜K��h�]V��MF΋h,̚y��N<�Z�X��d���|�q��]r�gQ�r��nWw	��Y���ث��Y:����)��v!����]��2'c���O5�9��dp�
V���f*�(3���%t�s�.���S����{����X�w�D^��_ҵ12�����`�u��`A�mˣL���w��51�\�HkV�id�h�s��D�Q����9���^ٹ�od����ٮ\��"�y*�Fhs��{�����;9�U�f�S�3�b���iX��`�5�F�@ޑV�͜�����:�)K��,�@��ug):s�^2
0|d��D5{7���y;b���o��f
|�\܅�^�ژ�jbf���np��qb�U�C�I#w1]�ڸh���O1G>w!�?�2�:f�[���ƚi�|n�b[73�5\�ή]��ݗM�m�\Y{���WY-Ȅܚ�_k�]�զ҆h�$|Ԗ�ü�P�uCKz�ʏ�=T���KFL�
�G&�SM�z�
꒧VZ����-&p�YK�jhY�������fѺ���E��+sq�IC�mamIaȯ�b	���iݲm,՗��Xŕ�d�r��c�SLY�Ѥ���,<�I����5I8�(�����I���W�S���������zi��j��B����)�?]@��	I@��1P4�(S�	��h�)�
��F�����{�(�� �]!AI@ST4,B'p�(� �;�-4�4s|��^n����]�|=t%b�f=��&*y�ٽ�g�X�{��X�H�'0�n�_}_}�UP���	�u�t��`TeT�U�G??ف��y����Nm��t�GN��r���L�oO����	�����Ⲏ5I�rc-%(W�u���TmۊyV�bs��ԷoR���y�ռ�sd�8��ɭ��%��������R������5VF)�o�V��;�޾��S;ˑ����e@g��|�|��pV]����ڋ,5�T����V�	�r�ɑ��i� ��u9ʐTtV]�'f:�����u�!�n�e�~�}�o��ǝ1~��}������vX����}�Ա��6+�f�LF�&^�
W�EX)���a��U3|�Q���Bu�Ka�x@�������42������͞s�/�������3�s?-U?E�E�Rި��RT��'�"z*q�����I[΍keD�v�B�Ւx��m�x:�}o2��a��)K����K�b�B�;�'��H��9�����.����b4}&��^lLs������c��|}��Mmz�ꓑI�˃��A_w��W���fw7�ѧ��Og�L�ۋLT���zr���՜[���s
Ԉ-��3�/�+�RH����Mf��l�]��b|�^Θ��uѩw�8|�3{O`�F�L�t<�	��?h�o{_���E��uN�I�sɦ�Ld�\hU�cd� �)@�P�f����e��n��۩[����rT�Uܕ��*;�q�t��G85ۻ���u���]��<��}���W���<��$�o���JB?od�}�ۊ��%�y�s�I���%�6a�B*6������g��{HZ�k)�RR���*�=�]�҇2���9z�K�X��J�-��xf���]U����{udk�F&�P7I�����ѧcDڻm�[e-�a����SM�w�iBg��
OM�7�o-�^��m`Z����+��<��`�3�OL�}���<�/t�,$w�|�G-s�'X�:ה����5v�s�쑽S_!{�J֒�S�9�M��A��
Z��n$ǽ�Ӯ��i�W������T�+u�"�u����(
e=��nu�Z��B������w��`��L�f��#��ں�*P��BRƞ�����湴���V�W��8�h;s����WR���:�����U �X�+�Nj��7+�l�n:vt置.�/1RYe`d����KY�Nњx�=�=!޿��m	1���o��b2��֝)^s�dﺖ�W�\��)F������y
^��n%�O!����\���7S�e�:Mm;S�s���.6b:�ccL_L�֨M8�`*��kP�R��xX=�
��=�Tb�Y�n%�߰^{��,T�4��*c��b�GM+o�'�`MK��K����Y٢HKΣ�``�o=I4����B�,��"w����B������L���fj��,�v>�ס�|�!�t�*9+0hӈ���I��u99qƤ��>������$��H.+�HB�S:�-��EvD��?ts���Ol����bt�d�)a�|�ظ���E����jg\~9vӕ�d|�
}3�y׈��+ӽ�}��
��=0���
.ǽ�VP{�KR�ӎ��r���o��Fq�i�n�es{�5��8޾�n�co�U
��b��){��ZZ�N��+�MyЎX�%F��+m��"\s�Kv��5��U�5g{#������u�h�=����=��l�T�.奈��\R�����.��G%�0Ωv`V���������:x��9&�)^꿰U��Yx�Nix�7�����9o!��l	�'�v���Pn��Z��}��>�ı�4�<�yH�p�������D@���MґU�ˣ����|�L�;q�^ѵ�x��Ŵ�q0��,��H|xgL�����ٙ��K�*�r^��~B�(�֞�Ř������<�=}H�4�V	kV#���g����^�mM��z��N��olw9VQ��W�sr6ѿS�ʽ��1����t�����<,2�)^f�/*�0�A1>Ɂ���=��w�<�i�]A�+Ӽ�[�~y�N"e�wk^4�M����O����/ސ�a��e�}���Z�ĸ�M_�<�+Ag���r4�]�>�V�(� �s�o-�1q�8M��v�~�*h�bGv 勬�OE-k"i�/;I��5Ժ��f(���2K6�eFi�ZD��ٟn�0��C��y���}U�S�ӓ}��P�?p�{����*<�7Azw��⣦�a*�J��	W��m�*��2!�0�q��on�p#�F�fy�q_���)�[�k/_�Zi����\�rxuֶ7�����x�
0�ĶJ�uI����ԃ�6��*��Q"���;�O
k!��վ�u�z��F7۫�V�����k8�a��E(�z]OrU���@QK �Cr�}�՜�b
[{.�7����kf��1��o93��L�6����і�nL��:Lw,�q�B��)4�ށq�e0��9���5lvbJ��&#cp�JR���u�F=1S�|]J�0�5ј!�����q���$x5]�28�֪|��g/��N��T��,*^���F~����ɑ&ۓS�9�D�t�dI���}r�MZ�����3]4�TC�:��Yy؁9�)�����H��]�o7��-YU�
/OA��/t�%�c���.+]6��f�%�!�~Էˆ�X6Z����E��̈́�F'�j7�cI���Z�`EŢ.5c���T�����4�����ʇ���>T�YWt}q����3����yb��a}�8ay���m��p֧;q'���5u�Q�	ⰱ)FuZ�ަڞ�"��{P:c[�]����,ثhT�^s�A|�幙�0R��&+,tT������vK[[�[V�q��gP����ޥŤ�$-eܾ��]�(�n���s�3�l�*�T�KF���_}_W�e^$�eFUxs���ccO��po]X�hZʏٓ�T��W��Vz#X�£Z�t�ֹ>Gjj1�Lv�{.�F�.5n�1@>9�O��s�ČB���ȮV'���W���?1�Dэ���M����&C�L|跴k�������'y\'��5d���N�-���N^D�����R�̨j{�Tc�+��R�Kˣ�˗g�x��t�6�^����_^n^m�i�S�����������1�0{ ة�1Z�������j��N��3g'ʯ~���)CEߒ��;��}��	���h�%����'zE��tO�f4�����������I���%JV0�n3���ب `�H�ܳ��{��5��>������ܔ�c�(������l��hm�.�]��IBpOlV75�1B"��j�ژr��6m��L�}X�.�0��u}jkB�t�4k�g{�O9=Tp�^4Ы��wTy�ˉ�.��=]�[����1\̆�ʴ�_�eP]�2x�z�ĚE�!㢣�P����] ��3���Z���<��d��i���s��D�
�2���>I�WӮ��q��.T�+�;#��`\v\����ߝ/oB��h�MW��>�}-֨�V/.���Y���v�X8�`T��2w�t�W�͊���f_�e:�y�+{��s��/�k�U{�ɤﯥ�� f����vN��PU�<�����Ү��1��c�+���0Vl�[��3kRRlUȈ����+/��j�&ʛ����ݐ�gjT�u32Դ,����� ��mv�^�O�/W��>�i�Њ�x�U��tTQpj�U�P#�(9�F!�	{
�M�)]]���Y�s"�c7따��/�:<إ;�@�x���RVMwe[af�#��
�Z��u���e�������aP���:f�+u5|aX����5��1]Ǫ$�4�i\7h���v���F�N]�P)y�:�5ٽy�[l><	a�r�A� >�VgAY�]Đc�.�Ց,\��f�ѣ�Rt�p;���R�h����l��'"�.��RG��T�ͫ��ǥ!i"�`���ؾ�qtR�EǬ_-}{I��0%[po*˥�(M�Z�;��w sEC |u�U����4ػ5�9IZt~�*�۴Q3�P��y�qSC��o4i͍b�ţ���-��ęh�{t��rّ>&�Pa3��&�' �Cj�E����b��c{�.-pV9�Vv`'L�/I*�[��F�TA`r]��`Θ�ӛM��o(�����,�^�ș�SV�0!@G��������[o���N�Y1}���bt�'��NK�e�2���u��a镽�r�m�"ʃ8��8x.�@Qj\�������u+YJ���2�t�=�z�:
#\�2�r�ض���Ns�(��,�!�M�;^2�2�y����T5�ǂ��u-�^b�D���܍�*���J��IW;l��/�3�'(�x�$�2�V�����K��2�+������p�M��N�x\�)v��V%G�O�7;��׿����ݜ�j��(
*��";��-Q�4�K���_R�Zn��i4�.���iM�-���A�n�
@��G{'	��#B1-U��@�MQE�G6
u��Z*���  
�>��-���=m�O��[{$H��F��ν�xO$١bI�=�ǰE7^_UW�\����۴��~���ԩ��b3Δ��a�LN>�ϫϋ3�>�[`�sCTBū�s�Jo����Ǵ��;i���Tw2�SIzv��Ը�vz/=q��Ǳj�9�.��ߏ��^+"g��.]=R������o���SV��^�:�k=1ʞ�.o�$���|��/���}�踋��uy��^n��߻�<����o��|�Ӱ����R��Wc�)� �i�J`#�`C�b���������RF�I^\��9F�|�_MJ���*9Yy ��#i9���71�*�Ss��kN��
݊�Z�)��0���t�9n'�kʗ�:���0v�u/~teDqD��]o��>�U[���g�����5�t�t㞩zgN`��m�7@�JS������ko>�.p
~,�*�e�L�45J�W�M{��;yUֿ��A��ע�
k�i4����y�����>L�7M����x#����5�<xz����D3��1������q{=jf�]ar�U��5�vι3�VW.f��臽WZ���}��R���)m�,mJuU�S��Vm�K�-v��W�������y�J;�������$���G���Q<�1��s]څ���^ʺ\���`�
��$ݽ\a�������qR�����GR����ݙ�7*��ĸ��N�b[�uh�Y\�,-��8�3�7��6�����i?y��ZEy�Դz'��*J�p/F����
\�Oy��d�$]˳�0�O.K���''e�,�oSK�xR5	�=�(A��\ߜ�v�,$�x��njŃ��̍R�\C��nki�֚��JF+�w��Sp$���͹So[�7ی���,�{j!�;j�{��kМ���Z���\�Ok��bc9xN<����W�~]��4��!�(\&7��m���%�U[�q��r�<K��aՖ��Y�'�yxױe2�x�K���Ө�N�W�ͤ6$���-�����꡵�
4
�}<H}>U��ω�VV7^1%�L��x�ӯ�Nj�j�9�{ә�,J�b�Y�����b�����og���b��E���c�r��H_������5z�Ŗ�/w >�ם'�c��)�O���N�N�kA�������<����tu�<�d�j�T(��B�0��r���e���ڞ�=^#�5ó���{:�{�*�e/�ڜ����y�0	P������	����#~��Y�3V	�j�jr��m!��ԹG�v���<�1:��ݍj��m��z1�itR�Q�>;q<���wm;z�}����^ʅ�b
�����9s#�j2\s��'j���'�gn�t�1ir��0�/A%����6��))��O0>K�{2��I[�}P�v��nue$K�p�#u,�m�\ �;ACޜm��u�t�?Ȉ��\�i�#ݝ1n���ҟ��h��,��jm;�\�6�Mt��=�o��.W ���߯-�k[�q�����D�{X�^-�j��ڞ�K+�qA���j�o�7jC����ԅI\WH_�gMC������
ڱ�.nb���nMvY~�7V�ب�:?R|���X�^�6�1�P�ms��x�����um?z�h�9�9N����`ph�k��Q�Q��׹$��X�^�H��%<2U����D��w�[1zk�"�4I��osU+��]�~TE�0hJ��ey��vE�x1���)�<9fC!M�@x�'riwu&�E��XT��S)��w�U�rm���w�^|���/���/�UU]�F���y�n9�\ǷM堅y��'�-��z��|[����O՝1S��t��EQr�y�jG���~}YϐU�i(Y��o���[�E8����gF�)�Y�[q������+����sru�m��ut��M�OR4��C�!���_�v�U�]�o{�/\�]��&T�E9��V)YԒ��h�y�u=���v�2�>�A�$�a{�o����mJ��Shf�U�e�a����=�:���l�U
8�5^�$��eg�^aWD��r��ޥ�=��q�V/w��/U缕	z�*���H����V��	QK=t�=�z��{{�БR钗;��َE��T��Z�o1S/L<�4���B���}TD�d�Ջ�~Ǚ;����#{���˻���+ 1o��S�aF�����C�\��<v��ދa�V��,47rv㘬��fg�9YX����K�1��Y�]21�9ۂ����ݯ���den/n��E��**u�p��Iwir{��wZ��E���T��8�lm�0���Vk�1�]J0�7%ꭒ�Vr*�Sv�>��r��$�����̵2�#�Ż�	��w��5[=)��g׽(�:q5x%g6�t,��y�zP�L�4��xˁ�����;���s�Fժ�ˀr��rh��bƃ�A&�Kα#��I����2��3��H��5��8�M�̘\N���ݎds&�����}��󯹧���\��ӆ�@Q��S�i��ipQ?OH��l{�;ܾ���(\7��-zƝ�r�e�M��2�{�Κ�at0�x�/E�{�c�7Nua���;Y��)5۩�I���j��m�csj�Aݬ�.��w<�e��I?Ep��˸B7�$^����~�n(kh�d�7�o��q?4a^uF�K"b�u��u���������l`P��H�#���F�xdMN����ݭ��Q�9q�"��d����Qx���T5�]�޿�f��|L��ls1zקe��T�Ԯ����.�7�52��}5=��P��ٯ$��Yu�2%����خT���!0-"w���*�,�/�Mi3�.k&�{3s�}UU٩I��L���Uɕ{=\��n�=q?9��z�˘GR܁��d��dO9չ�y�qN)PlLod����A��T�t41[�qs��9z��A5�1�<\[�^k��b���FU���YK{q���Wi7��T(ϥ��ۛv��++��3�r��������T��y�*$�G�����jji�h�[�i��4#a���c;nL�រjܡ+��c��~��F�MY^��
�J%LT1g�d���g>�����U�t��#���O=+�%V[ȽGt�<��
�hꪹ,ԛd��0 ��0�s~�OF�H}���t���A�<r�mn��]G�P�[S�Wt���4F1�S6��6&OA' O�W9"��פw�7��k���!��m�W�pt��ɥ1-l�;�>y}�[�"��A�L�LY㮄
�)J?-4�*gʽ�\�܁�w�6tQI��w�Z��\,тҩ營]{�_<�s]}+T��y�����X�j&Y��r��﫴g}\��ٽ�L�<�į��=֓}�jb�J�W�r�ql��Hhfm�\o�׮�J�:~ޙ��Z9s��Q�G\nȞ	�W��z]z�
�έߜ}���`����$B����(c�F�o�v��TG����l6�N2Vu�TG3r�D�q"Ob)�kxR�7�u�l��ۜ�TS�gݛ��%bC���SF^�c�(V�c��9w�j��	-tu�r��`�J��c���j�8�T��˸;oJv�V:�#��s'�nvb�Q��f�1�zˇGS`��q3g�fk�.Nnc/H��ݺ���Xb�����ʚ����U.,�sD�e���Sf��([cy���Y�m��J�w�&I�-9�\��p��^����Tcˆ���[�j-kMv�)S��-Z�XE�H�
�¾���|EpZ�(�5S`ʹ�Eai�AHKʗA�dwv ݆	��N��q����R/iݍ��=���˺���^��0U��¯Y�� ������rq���nn��RqLMT[$��9D���ۻ�ۉb(��1}c�%FmY����/B^X�)���q�̏GLܷ��Vn�s����m#���{%3ʶ,|iv�
�YV�cRV��bp�[W��x�Ռ�W��P3��q�P��k�8욓5MȐ]�W)"���&�&�3@%昞F�W��X���\�A,x�
=Ֆ���'n��%]�G�k�3D��f�t��G��1ԬI�{��ʛ�e
��E��Ȗ���Z�ə��9U��N��Z���cC��������fV�zN����Է���=2p�˭�P�`]G{;v齸���Ύ4/�^�0��[@��X�Im˸��K�U�ܬ"!�L�u�h��dj���P����n.<���k�����4nn�.����5qDcڀ�����y"�a�Q�Wn����jEY׽B�X����w{ݢ�����U�F�ؕ��h�"�j+�\��T�]���@�7[xr�qZۭ���+b��)�4F)�y��̜���r�$�¤R]+M*�޺A"%�k�Ѭ�r��)ql��3MfΊF[�P���(�w?�U��N���6�Bi
f����M)4�htև�))�{�T�_v��l�6$�"��[cX4��bS�4�Ս�1�[��ryy��b5CE�ƍh���-m��Xƌ���:��<�'1���9rh�cTTE��������*���!k��]g<u�\�%;�]�u�7��<QCwnX��w6�R%ݸ�:��p�ק�?��痥���O���;��f�;���\d�s���Q1�Np܂�����X�qo��f�Ώ��Y2������쌉}�ЂZ�wR�y�.ܽ���~mm���(I�_o��^�^ei8����ތ�mt1�~�r s+�b��^w�:/��:.+��_���3S�e�{�>��|�l,��^T6�?�-�i�k5c��]a�s	��)�1{װ,\c�<Di����3dp�Jfy�E��!\�i�E���� [8}�D�Z�馱̯gO�����V�5��9��*�ri5#Q&G�H�w��p�(v8/P֗[���3l�j�h#f.LoU���m�)��q)����9�[��(JX����e%e���[�1Q�'X�����a �r"�Z�h�q*��i��f!�=}_3���'5��ZY�C��1��FmX�=�6W*F	���Wm�kĸ|��e�k����k�5%x�b�)�ß�0du^��A��533om�֠}�|WX̓��_�+���̣��qs�����f�]�pg���3��e��ѱ��M=�Ҩ��-䊙W���%~�ʛPY:���ۓ������XK����M�v:��b^�F��r�RM���P�vol�L�ZoN@}=P]����e'�&��h�«{}�a��*Z�U�+;Sʮ���ųmu@���تShmm:���xx�%J�ɍn����/,��Y�� �dud��NV�rcJJ�~���⦧?9���ɏv�9�����<�}��9��Ӈ��ln�?>�f\��[=ӟl�n
5��s����b�����1��ڤ�������C+ȃ%*��9���v�bY;�9����eI�7M�?_��}����5�o�1>yE�g��.s�J�yWi�c�?L�h1c�K�\��MY��*ӼL�CR�5�5��=��앺�^���\�ݮ;�ʂ��Ӭ�O%s��q�9H1�kW�}te#�1���h�F�V�kR���[]���P�O�nB�7{W��K�t�(PىT��IL'�i7Zߢ�L�鉻�59�vvD��n
rŃ����QU�g�5p��i9����>��-̤�p��Y��s7y袡W��ݱ�$��������K��M�^��YC��&b�YW�ǾǛ��fqՎ&ϫ����.�ވz�@�����L{����;7���|��Q����OE�����=��������J��7n�е���k���ٷ�g��������Co͞�K�uoe�V�Gg�~��W�N��R���������Y=��
�pG�O���j�F��J�y��
�1B��gըx>�P}����6bˤ��B�g���a��?5=�Io�t��S��Iլ�&�zQ���9]�� �9lux�Ŝ(L����T�Ysz������k�-"���}]nR���;�M��M�pU�����\�L���}��j���kS��N����_���ի��sY���w�?S�r� $�#��3W=\�IGbm�������r���t��J.q�ʄ�Qڍ��.�a���.�Zc�\�y�����Z[4��Ln�H��;$~%N��Ա�ߍJ��I��1�TJ�Gs�oz���NtG�Z.�ڻ��>�����ӵyU�QpjR����&S3��;$�*�������r��re[�]�iK���ow��=�ei"�5k]�����}:�滱٫��^%���j�W5���=p!
�m�#��	�Z�T�b�hl^�sW��o;哒�NP��0e�*��s��˸h����F�o-�]8�=?�;�y�{:%������m}:����F����*N����������ڞ�*h��_c�)Ԟ��R�Tϴž9
��G��j�3<�Y&��T���
���u�Kr��1B��s{�8���L[j�:\�����=����=�<E/z��q�=끽?ol��Y�뀦F�0��觗v�.|�5An6a��͹���]�B�]y4�5��O�&#{<��zh5�j�ˏ+�v�����]Q��2�;�p�L=p����u��ih��kk���b�NLS8�v���wo^��u�1���$f"�Ĺ�����~�J�1n��B-S��7f�c�k�B-z�<#�.ء�.[��zS5��]��,��@}���=cp_o��Y�-nӿ�ŝ^��s���TӼ�.��e�7�sT�!����[������ȚܑR�'�T�؝�f��p�M%q��"f���nz��Ƶۋ�^{�VWA^�lŖ^��U�N�a(H߽�C�C������I�v�82��#mV(n��79�L8���)c��gطl���x����a�\�ب�sL���OW���<�7�y�l��ꤲ�T���z��(p-{Q����>�%�f���C/���;�U˺ԓ�+J��Rz˗m��z���r/W\"��/�PۙA:۰�Y��e�s}��U��6�X�ӥDt���ȓH�V�v��m���᫡4��v4s�N�jp�Vfָ�ƚrT�����森~}Z��;L�ܒ�#}��x�ܛ�_Î�ڼ�*�c����2r���s C��`�px��x����m-ء��ޤ�1Pr*�)ݮ1���)�ʗ�m���.RD��:z~���Bз1h����gOO�^�3^��L2�]{�ǻ�
`ל��y����B�?R�YJ)z�4��h��e y'$���Tŕ��Һi�U'�}��[.:NT����������ga��c}�T=Vո�};��y妴�w�C����C�vzY4-'wcr=f�2��akJk�L�N�׈si���_���JU�Y��Ƹ��U5D{���oN�.cI�G��{�ԇ7�C�́��w����.R�������Xٮ{�ZH�!U��:�.9�+<1����,��m���pWZ��g�c##ď��W�4��S�{1�u�V�/�T�?�?Z�oe����������YS�3]Q�g{;������c3�Ûb.�8�	����f��9�D��79d(<�tF/?���j�{�^�N2��U�y�eu�c��Cn~���r��w2*�Iѫ}���0�'DBQ�/o>}�<Ui�͗�v���C�R�e�-n:��q�w$o
��+M����]q�-px�N�9é�2jդ��r񢹻T���եtq�L�r'�U��N͞~�p.ۡ���MJ��7 Y��[�&��N Kc6�;��S(<��_J�|����;	����ޞ�?���C���{(�C�O:�W��Y��yŻC�ޫ��vb���=�!�o^\���j�V6�ț����uk�K��.c!b#|�qw��^�Owh�k��1�Y�슗��b��;|�noeO_]@ђ�+��$��9�I2z�Y����ҤΨ�(�ًh���/�ޝYެ��f9��-͝S{MmB���R�٧
�U����އ^j�}�|��'�~�����ߧ]:m�_�Z:��}<���y�E��+N{$ʴ�5�^��@i�8�F��ˁ�'��,ײ
W�*.X�!�Z�i�F�B5z͘ zػ�g�
��ʋ{+�-�M�!��;���8yZ�q�a�̨Us݆�
O:��0iA0�g��b�.���]n���=�y*f��Yr�g3�c��1Q���l=ɭ+cn�:�Ǵ\e�B�����j�q*�������n7c"�9P藋��s8H�i6-��;2KJ(û��ʼ���wt�(�E9��A�m�s.����e�Y.Ҩ� mF���Mp�0�V��v���]��.;u8s�>6M�����+f�p��'"�[�eЕ,���}wN���{΍GV;/R�fo��j��}�s��AV��*�v�=V�'(��sda"��R��i���I��l�X=��$x乑q�y��4]�c+��0���쵇�'}c%���:>q�ZWv�tB�ٳ^2���t���Dj�l��tCt36N�;
WՔT K�.��~�M>�CE��7�l[B	�Hq/g3�����R�z�}q�o+��ҍ3�����u��ܫZME����I�Λ�*���������a�*s��+*"rT�԰�p��ՖH��&�5�٧V� w�抌�'dsOf��g%Kz���;���Cu����Ƃ�Zh�Y�����g��K��a**o&�KR_d��Ob�q69&4
����u7(�9���%��)����-�4�; 3���/z�����U��+8Z��,�`gK�y�~km�2+E�crY�@2;�O�Y�yV���:�{N]\��/&�A�����]��e�K����˛B�]fu�ŀ4�`�]dx3#�y�_+>��[t��x�v� ��v�e+cВ����vΕ��z�9=��a!�3��_��G^����+�4RS�KmkHEl9�giq?lC��r���4r�ITD�W6��`���1�Mh�mFر�9�p܍$PTk�QUs<�Q�֊͊`+�EOv���TQի͠�����b�&z�T�
���*����l�<ڢ9�����o\����Ԅ��`�׼�"5�g	�+W,f���B�s�If�\�[1��W��M���p�6[=3nF��|�vmTa���ŽRĘ��E�A&���[c3d�S7�.z&[��V�1{��U{���|�#���ƫ[#r��E�<C�P�[y��U�֗vq�1�Ej�2ꡦ'��;.��7Pk��J�lQ���c ^�Q�W�]-Sg�[��f��Ң�89�5��2D���4�h�o����f�4���!J};���a�l-7�xS{x&�/{������>)�/��b������K�z��Sah��(���u��+�>;��+�������|�|)�A�k6�$�C�%OFh1��s2��!��]1׳�\���+e��W�҇�Ǻn��]^���Jt�t<�����Q#�d�^���VW�E)��O��0��`n��Ͻ��e�����*�K�	VO<�Q�tO9�)���Mڗ*y.�� wOq1NXq�J��w5��^���/��7���~j���&�q���׵pVG:�N�'�O�\�a�뵩9Z�^�:$��S+W|��:�{{���&����u��0�_M�iT	��5����u�8
2+*⥕�R�s�"�YB�R�a��Y��`oO�N��U�5,�~aɋ��{ό�������Re)�ʫܭ��wv��V��t&��Z���b���K�Ňu�����mv%�wY�՜�P싯���T�1�2��q&ne�6��$��8�(d�w�/ �.Hk�MIR?�r�%�zg���^3S��T*_+�C�o� Gf)+wsS"�������}�2��PL,9��u�\�d׻�	�A.y��Mw�W��|*��=�jH�Y"F�~�τ��Ҁ���<է���tG۱W����mVQ���Q����7�����Ν=����{q|�f����t	(�k/�6�-P�a�z��V���|��O��Q-Ll�9�'����b�w󾘭�*��3Z�2�1�CS ��˭�dS����B�L�k��׏a꼁�@;m��Z{�Ȱb�E\.��y�k_لal�k�,��:n#Ǩ:�x�}xX���{��.����w�Zؗ���\����-�.{�;�XѺRq�'3�����+�Q~���9t�u.U�ب��W��Z^l��GBm�S�b��h7�"n{q�n^�C�]s}���"o^ɌAKnQ進:�7*���)�I�ښ���3�j��U�'Re�����WQ��d�2���zfыَ�>�'��*qeΆ��[��s����5����k_M�>�7ˠ�yy;['9�V�-tV��w�n��jq���Z�ڟumr6�:|�'=๐�������l����˧�¾�����{�s+�N��}����ҳ�r��J�>Ӱu�+�#lWW��(j�����+1J����Y}H*�ԣ��c�C�_q;�o@b��;�X�w�)N֪�0&��k6�;뎷��%�	�'W>]��B���R�����(R/O�z[Jg���*ji�M��%j��~�V�E�I�r��6���ښu�1��˒��t�0F���<�:^�\�=��c��IE�~��jj��w�Rq�3ݲS�\��wά��;u���Os��/hlmqԵS�1oUx�s'JW����r��z�]�h&�Mg�x��댊η�=J��[\���e��k��1�J�{�����i���z�������uxWUӓ)��X<[�2��c����Ez�cJY]�����10Q.RNދ׀��y����mCw"�i�g:%��g�80��s�ay�.fܬ��2ۆk��l-�"���N{��{���MW��K�GP���V�U��-E�x�u�W�o��Q����SA칳/s^g6�X�S�ѵQy���9Ŧ�ݲ���Ҕy%sς7�	��d[����L>t/3�/��u)ퟲ�Dл�R�r�{����{-���i�+���N-4A�vM8�/2e�=��}[{Z���$ڑ��t�R���NZ>��'Q�UN��f�M���$�483W
��ܝ.��؞W�Z�;���L4�,��<�����S|�߫Y���@�!����ZRV�E
T)P��x�����\���Jv÷�Oz���9��_6������m;�Ʃ�{d�ChK�u�I���ѱ���A]M3���7�E�����A���y���Y��pP1�S}]rr�E�[.�9l�g�z��]_P��h�y��J34�\�^H�k��"|6;�g.��[��7��v`ȋ�	>�WӞO%*�0} 2�4iu^������1�5{�t�C���,SQ�"p�5 ��V[��v}�g:��Uc��伴�������;�w'�Og�&QƖ�0͖q���I�L�s0w,�P=۸q��WTӖ*��K��{�5������N���⡞�\n�y9�=i�+}�K�T�T�M�J���9�6��/=D�x��/��-��#���iv]�Q��,�I���l-���P��U�;��@x.|��~g�,��f�\�2A�U����!����V��kkgZ|\������1���9��v�)xQ����;���4񍥪�%�
s��eg�
��Iܘݥ�=�50/�j�w2��g4��g���ȭ�w@���ټ��t�c���o^|!��v婍S���wcK��Lcn5��#n���gr�u����KR[8���c4ܑ6�j`w즻_�_H�P?W��F �x�HG쎝܎۪�jRm�}&j-p4�kCJ��r��5ݯ��']f����tiy=N9�x��ڤ�{Ʈ��:ŭX�ٔ�/ڇ{h�O��{J`T��T��w\��a
�ŗ% ��R9GWPk�$&�[*��q����ok���WP�=̹Q�Kk���R�ƿ����Oj���穥}�A����L)2�ЋkUݥ{���}�cX��>϶�]��=�}�X�7L_�x���epߊ)���*�ޯ
r���JP5���DNh�a쏕Soy��P��6uM�5���G!���@�x��z��k�),�IQWtZ�y�j9ܸ�W=�k��������L����sԺq�wp��7/kZ]�Uf>nθ\�+�4�]xW�#�M�i7<�s3�O��ٮ@�N:���xP�0��֒�jӉ���)g/�n0��P��<{�o�G��P�ȍsjfe�/MOj��o�� �c	�y���eoܧS;LV1f����.¦N�~@��F�,w�+�֭�[(�f�hB�t��M�e��YR�n'����MwwsDEi��Ġa�j��2�K�0�\��l��q�ה��7P�d���c�Ka>1��NqFO^g7$KȽ�ö&S�p����l*�Bg�Oy��ݴ�xR�!tu���\��׸#�F�߼s���^����Ӌ�]N�A&е��{��^������s�c��~])aSf���N�wRS�ê��S�W�a�~��7�i?M�9�*�:��X⣣�1��s�r�N(��瓙]�����Gs��3�i�n�{\+�rxgz�������*K*�{(]��9���s��~�������|9˺µ���1'����n𮮎i=��X�mB�Q�;�OZI����*��Ǹ�i5a��.��w��Z#"��3k���r8l�Gs���ס�w���M ^;\�G�ML��r�^�.���V6�ٻض��k�Cˬ�w�sN�[����A�N	��� s/r-n�a��gF5.�8f�lꛑ"�v��P^f�m�ot6��o�\�OW2�/-�O{F�d�JN����Uh�C��𘃾S�X�~3�!%�;Q�7e�r�u�DXF%���-C��j&�V�r�.2�)B��NQ�uY$�o��"y[��+��+YZS�	��2ĭ�����'-����uqa�G�2q���c���n�k�(�DI>A�l!OKᆗ�[���V9�Zy*S��d��}{���L�t:*uZ}�i�N�dEܘv��e�]����hή����� I�\�,_Q4�D�Տ&��鹼؜�`Qz_|P%��C�hWQ���t�R�C;G"�B�cȵm@0qrHu���!
��r����S%_C���D�me�Vnq��2$RV��nRˤ9Y���Iu���hYF��gF��1	X���-�.fv*2�[�,8 ��Uî���[|t�R��׍*
;������%�`���ui�ͩ�i��� �
�V.`[
�>�v��ux�u'�c���iDf��tY�ܳ������thu�!�x��@@�a�\
�!�弦�C��&��i���W3���z܊p�k.����`ŸV�����ɢP�H�f�y�#�`�So��Xɧ��soAqW'��BH���L9b��e]�����i��e��9pW�Eb�Ţՙ �;=��5':�7�]�e��]�Z������{%&����d��̌K���"S��3�fB&S��o�Π�]����z�K:�˨��R_;��Y �%ԏq��t���n���Ϟ�ﾻ��bH���B�(���"�����b�X�(��X��&��k�i���&�������b<�h������9
"(����Ѵh�(Z)�"�fbjb�gTy9�	(��1$P3KT�QDU���r1D�SUTTUT��UP�UQT��lj$���Д�Q5�b��h�h"��͊Z��֘�����C�<���~�J���X���<�*�y���e�p��N��|�H��,_�yn��k٫s�d�}ݐ;�8�g�%ڛ�bLk]|gBr�NnIn����L��NOa��n;���#�^�u��3ʬ�Y<tV���]R�ٙ���|�>?Z��c#f!�Ϥ�H��
��eЦ�Xh�ӱuv�L�mV�E��J�8K?�Q��,�
�W���MZׇ���i�S�py�0���ف��jϻc���X8�����+1!�Bb��FGBS�Lb>���x����U��8�mO'O��R�[5:�:]K}k�[�{FA1�;�x��ؾ��W���u�{n��'�g)��rq��Z!�tpǅ�ݩH�{�p��Z��֔D�����*��3�����	�4�e�(7��1)��M��Mg.���F)MZ�K�������d�0�5�_��e�;������9=�޳�F�o!\3��-	��8�3�#x�1��\�h�yT=~<]�k=����S�RMvs�F����U~���{Z1�B{�&R���`Ff����4��Q���d��$�Qg�5�徸�sZ���[S#5v�ǑS���RWF/?M㺺w�\kg`,�gy��E�ZL�w���y�8�w����r��ܰT�֞���-��� ��53@٬Yս\�-R��YE<i�W��+�r��#y{<e��ߩ��h�fz��T�U����Ks,�9Ύx�Z��݅�����W�{����=f�/w=�4�S���;�=H�Z9d%(h�_w@�]lΠ�����%Ksy5׻療��k���=n:�1R+��эq�c������#Z�=�*�8/��Nv�o�n�R����m�3jO\���E�V����ת![(S�@�u`w�\��76ro��(��ُ���/3�e�b�m9o6���cM��ӵ���\�@�F�WǞ��f�?n�N]p�y�t~(�gsS�j'�#����Q�{����/p�s_�십z׫6�ݛ'�O��L@��R"C�u�~h�h���7����z�X^*H�Wt}<�j7�G�XT����:EP/Wi]ze�ܙ�����5#{M�#kS�KD;s�T�������@���,�]�Yq��Y��iu��;N���h��Ws�sS��XQ�z{o�m�>U28��RM�~|i��}�ŷ!-L^N�i��eT8�ז���>�ߪ�?d�PTj�lt媧)g�*U��9��RG�n�G��!��7��7���:��}�8�u���c���3��1����*�'�q�u}�-v��C�����>/�lj����׷��g����6�m̧6ࢼ���V�k�GC�?)��c�Fwd\^����ۻ�}wV�y'oh��M�t!����c�гy����>�q�Ϗ�?9^x�egj�zzf�^JM�n���s>T�����Cէ�6����c|��W3��C4拊S9�m�����Iu!���th=/0��η�
�ޗ�^I� �?�s���χｶ�[�h�ook�������C�!���@s}��G��B��B��Ŝ�WG��m�N�}�y�)�P��-.9�6�V?zitu�:S�dw@��g�CTh��^�6�'���k�F�ʹ�-�ژr�9.����������2`iŎ���ق��K�p|�a�4��YO����|���sS��߆�LD�ɾ�R�wsk���p5d�z�>UBK�6�Ĺk�k��N��4X�<���V{e�c��~��Ё�䓋s��}S���%J5�h'���������J���ZWKvq|:
[9[Q�=����ji-���lЌ����<n�jG�^fE��k�t�Ơ�x��]̀n�̤x'
�����˻����eNb��g������R<ek�:s�ؗl��?d�����ګ�����yJ4�	t�MWS�h]8�=~�:��&4c�~�S�u8�!]ߡNN7~��: �S�Δ��M��ǚv�=��z
�=��3��>��m�V9���"e�m���j�[fow#ʦ5Fn�<g=�%��n4 G��{��}�{��]qI��z�r���ܭ��z�g�eǣ<by�s�\���������9^U��WKTx�Ǻ&19s�UΫ��,J�^%Z�*���.��`b|���mZ���mt��ڕ���r��WNP�a���6]���[շzdY��zPa��]`Vë���+d*m�gvh�tz�p��sQ(N̽͹�Q�32K�������A�����ۡ��G���<�5�x�B�Tk}W=�Ϳx��J��ϣ��ؽj�ޞp�˲˄��kw�P\-sƫ��n�O����_[���z�<�;�4c�o)O�L�	�Y,Tm
ƎF ��(�e�=[Zh�]y�Ց����^�f�-w?op|��m��D(����ћR
�N1�z�0oHO�j��H�U;�WZ㠵;�Ԛ��[�-4���M}��J���̬7��BV�g�9�^��[]�o7���Ʊ{״�s��9�w���ҫ��0e;B�8�N؂�ֱ��uyA,�B'��r��'�̾��������,��"p�0*����9�8h�yW˄�̹��L�d���������
�M�}� )t�'�_�K��e��Mq-A��K�8�f�y9�V뼙P��a){{���>�}��|u�Ⱦ������~�~R;�W�E�Q����2yg��42��&H�=�y�N��Hc�n���ϐfϭ��=��O9޲r��I�5�Kd�qņ�a����yzI�̸do;����'�l�'n���,ja^)�y.�s�Llm�Q�ܗok|�އ�]@9ue�7Z��9�3�����������|�U�1�l+	{�q�2*����ה6[(�	c��j�j�΂G1U
�_پ��k�\�16�����^nt�(ooVm��KL��|l���Ҕʍ�g�{�&���>�]R����|�ji�pU�ok��qRx�\Wν�Ʌэ����U!��8=q\�/���O������,P�G����#L�������/��8�c��TL��N�o����Y@��P��U�m-V ���/���@��aVK���P˙���$F#�~cF���F<���HC1�tV��𚙌�Ϊ^
{'e9�^|��гUh�h�ɉ��C/�&`����<`zwB=����Ԕ*��j~���o��'�5>7��4����5�u��e_%n6��8m輨�F�x���g��*�U�1*~=�ͩ�Z>�cq����Xc��M���b'�ۛ�P|��:g��z��چ����업���e�s��վ��{�t7FhS�WjW�>�DL���fg�l�`��`�ܫ��}�9ĭJ5ƥY�at��[+�r}?��~֪� G{��2�1d���I�2}b9ѯ^�I' ��������qDǂ��c<S7`�
�Vӑ-��7�}#�Mx�:�π���) Ll�H24c0Q �{囋�����*1�v}�f28�/�@�'H�jc� �@U>�Y���g�TL#�lx=��P�'���c���A�b�W��8��ٛ�����`��t��ѱb���j2c��\xw9��e��s6O�@�'�L�߳7�����1<}�,ҼU|����?oկ�\�
_k^��H�S��o�߫�:6����g�#d߫**��V)?\m}��ي��y,���M�YB)��H����A��*&�;U�{���q��3Q�P���L!�!�y`UdQh��]6�YK���(�~��Z�ʻT:i���gMtUQb���=ʕD���]�r�!��&Jᬕo.ҽ��q|�[W�v:zX+*�_wW3eՔ�릚��Y�������5�X���8F��*ڔ1�Ι�Qa9:�0�����x2�*)�O���Sd�:b1�^��Q�PC1b���&B��\�4�L�z�^�J"��KX�t����i�xM���V��w�iB����*r�ھ\��'�>R$��]���AYon�|���Y1V�ԇM����W!]+얶#�;�ާn���X��Dm�u,�&C)[8��j���sw4*�[���l:β�k��鋷i8�v:"OK���F��-v8���� ��J����2^�4��Ũ���d�BO[cefX�:)uc�W-e<�`��g;�c]#�VZ��ĬZ~Z������r��s�M8v��L�̫�gu,)��35>���)CHF[�>����s���
�흻��9#S�L�6�s.�R%�;�o%q�2���X�(>��73��e(����*���[q�Qߍ\0�z�NeG\5�u�(��`��@q��4w�n�������R��T2Zͺ�On���b��A��vͶ��Z$�=�0�lB�:�-�����zYx��F��_�_s��b�C��OD�����N�ų*�e��J�"hQՕo:0|H�X�w��n>�s��Y�[Zu�P��E��O� �;0R�����-�X�*Wcn��(֎fP�V�o��U�7�c[�GT�1
�te�w��B���kuː2r�p�Y@c��(�ծ�KSws	�M5� ���xA�"ݥJ��w��Iz�Q0�)ڕ��ĉ4�\!W���^2��m��J*���]��&��F��cM�R�P��=QV��.ҍr�K��r,ӽ���\ƽX����%���j���DPQCLA@Q�LC<�R6�SEQQbU!Al�����G����9%:v5 �G3�m���<�I+�_'�놇�VH�j��i���ִ��5���

*�[�K�ZCs;ll*�N��p�WI����:((4i��6iE���h�3CZ��*�'�<�����,C���h�R�)T��`����Zh��F��b�l�4�T1)M�c`�Dih	�I�5�T�;e4V�N�rDV�ƍ\Γ��t����4i�bJ4lg�|�m`e��h��n�Qr���;�1��f�#][��9u�������_�����N�+�3�ޘ1jP��9�aF� .p�g��-�ު�(�t��^����h����?�j�2x��k�y�ު���	���������+g�<׼�z�y�x[m�]
=�
�ԅ	�U�����UU��L�]���c����<*.�&9r�Y�<$�;Ƒ��B��>b�9���z�r�z:���na��j�c��0*�fzb�I�������Ẽ~���<�
K�B=��H�,1Q	�_{�2E�L`�յ=��,�>^cp�F�=��F��
��ɏx��ra��[��S�7&��i�~U�ׁM��Aߊu<E{���ˤ���{ts�>����?z:	�Oi�&9W��U��,躆'��b^��~W[��U�y�? 37eI,��<�i�5r�6��g�t�&T%�|�p�~3�j�D �pͧ��:Uf�83o-)r���L*���fYo_�ޯ�R�Q�� =ĈH��H��@��i�����1��v�˷�FפJ���/H�1�(�wg��'LK�T'zg'�}��׮O�O��:#7�ƚF���b���du����$��[�'x_1�裸�/=(V�Q��p����1��pzg�=aAW7������W��6����2�YЫ���=��-�*��Wg�s��o����6��4���V&�iW��Ɖ�u!>�ji��P��j�j~����A�.��B	�`֟���]��<�]�8zq�Kƽz��b���ڦ�q��dL�B�8R����|��9�zn�/)�0�lF3}n��e��Ö��٧��w��G���<�<&�uK���^�o��s)��O a�̒}٢��_�2�zU�bTť��Iu`*]����$�(m=&=m�WmAk�+���1�o����\Wܳ#=0���ff
f�N8�Q;����\չ�9�� E~��s����@��8�aNǜ�������.��� �l����1Q�,\� p�dRޗ�LM_��w�$X�s Lrpcr�u�M*!�806�\I��,�z�z<ܝ=� {�0�.@���xm| �§1�~RQ���.��3�P��R�$���LoX��Q�'�s�l򚝚^�4�\���O��:]E�@	�#ԡ����؞�j����<*b���Č�^zo�,r0/������5�	/R��=�}�t&� C���E���T��ًV�j������������S�aR���ԫ�U�\֖~7��۝�v�y>�}~�ベ��N����HCN�k}qVx�Rد��\��7jY��F�fPEEm�V	�a�u0��o��q�.��:k{HLf<��<�G��V��Uy�)�h�0m23�;���vʊ�����o���i��>(J:�ɋ��t�2^zo�<�������$�yOivk�|kf�bqc��U��O��7O&����ސ��虃*t1��<3�.c����ާQ�4h>���xh�/H��R b<��f��K~6܄+�R{��*%y�쪍��p�;�Wҽ,dA:&"�^���QUR�j䃃�@��c�^��@�����+���L�MO����|��\P�E9��Y�|;�e�&=��$	ٌ�dh�s�>ɚ�����(��1X}g��r�{��0��4_Yу_��ý]�KS�F�Q���aI����P�*����&;��9�w�џWVc��=�,~�.4$P��~��d��>���`""�����GlѮ��Y���fM^�S���`1���ǥCJ��=(�Fّt���c*nڭ,��C3�[ۡLꮒ�u�<%�#zak ����w&��_�'=u���b>�,��Lh�sVm�7�Ԁ[>g���|�n�O�G:�.Ll*,�&6�*ʋG�qH�_Ju��]�\��/y���f�ҟ�S���H���yM�A��#F�@OU��ｯ�Έc�3Q}Q0�u��aޞ`���A�QJ�'���K��U���wQ{:����c��Y1p�K�k��E�ڦ��π�>���D�0hڴ����_�ފ|P_�Fs�ڇ�~��kZ~�^�����9 o�b��<ȣ�+҄k8R��J�|�;�1[�Q�����Q1��L�����^/�cPcÕ��x���n�xq6;�xxu�ŭU
�� ��1>(Mq�	�/u�W{�˞��1��{&&�4X-L1��1D�<P�Fz߷�W>���,�y�U��ǫ_��e�!� ��1�ܼ�J�)k���v�k�h�cighY����>��j�e�%��.E���H�Z�iq�V�-��M�gko����*	l�>�ʤn	a�?H�0aH�Ϳ;�����%.4z	�h�G�ޖ+	�&l�1^��"-?h���Vn���<�Lz!ic�ڔ�6�\�U�1�:�z��:TX�s[�u�P������*�X���,��'��zj����|8�����X��$Lq�(�#�i�����������~k�B���_�:p��4�� ���@xtA���gw�=��]��=�mP��-�Ƙ� Ti�tE#���F.:����vҼO�9�*}az&pe}�B���n9CA�ct��G�^1g��<ܼ=À~8�U���d�tYЫ&D�ai�mUF�6i{����U�Dv��W(�D���x	��b��c�1��afLz)Qy`�bf]��I=f�u!�:�j�;�]'<'�;X��l��ڔ�8�S{��ja��O�����+Ia�>��iW{�e �%�����S����}��t�~����"L��k3��N�����h�=����ˬ���T!=,]�LX��炾��wH8C�����	y��\`C\��Qf:u�
gMl�^�P�L�M߂�뛟{oټ��^�ȒxmƊ��Ǯc�'޿�΢�2��������W��\��y��0ъ�8�|*��0SST�n��{c�ov�h������4Lw���+���#�\3=��~�#4����`@� ��ߡ��JH�l���ϲ�ݩ�P�u	��I�O����+H�90���l�:��g�{~�#�&j.��G������UE��HU�<���6�{��jv3�tĊU7S$V��W�*4��9F�Cc�S�S�����གྷ�� �3OZf;�o}2&ʾ�r5,A�4�� ��g���������sm�b��>�nt�m�[�����t(���J:��򪪾��3Z>2N��+���s2��q����P�ŇT���f��]�� ȡC�NNkZ:�F��b�% $��r�z2��Wy%~�Hп)���������a
�C��s����\bq�]��n�5^��za^N��jppb�����.+}q��ӭA6}k�W�{홆���LS(O��b�&;
�t�3 �g��[�z|���u�	��f��	^�������:i�e��]/w�`Z>.@ʙ�>�0�ع�s؊�:�����ǽe{w����Q��I�ꍩ !�EE�Rhl�2�gXz]�O�ow�Z����]���C ���+��2��0��o�]Z��������k���a�Ҵ����LT�)���f�y�=�)݉���J�t�q�;�^8.2n��W[e�Jyw�ߦd����}`�8�"�eقT2�/�2 �h�uI8'��fϊ��'\�������}}�>��W�b�ǋ�Y�X�pe�&#ޘ��$1��hr�
7�M�q�RD�:�VY�Bbc�^�n$Æ@�M_@o<ˮ�*3�ϤXb���}s��-��^>����e�S1��9S���(��}�����`���lX����k����`xD��zz�ϐ�Q�q���<#X1�i�s�4dR������Q��|�!ɠ�||\cv���;�ʊ�S�j�.kV���^�}^/����0�����V}��k$\4�r�Pgǣ��.�-V�}f{�pܙ��Uβ��7Ƅ�s��܇�ةm>IKр�阺]Q�,E�8!}~�1�y����ހ.��ow��� �E���^[���,���z����Gc{������v�뾲��h�5��s����J?LG3�,����'���Ǉf���	�:�(8P;��N���Yg#F�xN$M�g/�\�KOZ�s�{3s�i�W*vϑ�OeR1}D��5���� S>te{)�V�[ܝO%���=z�X���4d/UC���c��w��Y�$X:���z���މ��p�)�^8=g�&.W
��0H�q�����J����{@��ax�ɉ�쨤X.���Ђ	�ƈ����ͤ��{� �����<��Q,1I��Ld��0߮o�彼\�d���.$�D�>b����1���5u�yw��޴���i�b~��5�f;"*X"x�3s�W��nU�},��wzH�G��E:_J � V�yإ�K���S�ڃQ����ڼ�z}=�ա��:k�p��H���Lr:#����d]��ݼ�=:|�i`�u)��L"��*Ţ_h���;����ki\��H�wvl~�1��@}�~[mIȁ�3OϬ*޴V��;52K��J3]��X���\F'db�n������>,�Z�gG|�����㬛�����Ni	T�n�ܼP��y�"�� ��vR�a���h�}�:Z���F8��?'�'Q�) �i�u���[��۸��}���`n��{�d\�b��ɇ�+��\�M�0;�"�R���]�3�/JxLU������$ejF��֏��Cd��57�!X�.+�:�NA&v��.���l���Q�i�\�xw�w(�k�1c,�fL��Rir���mR��^^����k�l6�]�璌[�j��\�_�����4�k�t��V�"��#�,�)�95ܠ�,�b����H��W�>��R�V�)[t���I{�<��_����WX� G�*���*�P%Z�/��muމ�����V��z0
���ٹF��<�.4�<���Q�F> ���Z����I�2�*.���{o.8�A�bX����H�8��vu�t[�����4j��`��'��̀��/������A�G�7��/�n�L�79P�/��ZtA.���\�ĝ�z��+`<ea|E���ޛ$�-ǔ���Y���znN���e�r�:o*P��2!W��E\&�5{�h�^8�[e�`10hye���jHS��aQy$<�3Y�O�P�� ;]̭����i��YA�Q��M�P� �Fo��������S;�=�+d:�T��]:`�1�� � �c =�dE�N��1Y�X� �V8�f0VmB�1����аv���
h�2�8n�r�ʷ{��v�s(ࠒ`K��yҔ(�Y�I*e���Γ��#R�bYʋ�j�v���QazMv�Q7�� ���9��U]N����:�E�w�!�4Vt�4�K^\�X)���*tbk�9p���i���ض�5��К���Di4h�O#s�h+�jJ99�ss��T1i]4��U�41m��:J��W 6�J9��r)�[FnZ����6�9��>@rN��Rn�P�R�.@���DS���+��AI�I�4��y44 ��i5�)R���Ss.6NO)������@j��#�w5Kɡ��A���@R=HA��\K@�R�uKIN�*�CE ѡ4���Հ) �.��aR�)B���^uν]|��χ��wﾠر���˛;m�� �;d_,|�l\�I��φ.N�\�m{��ɢ����i���Q��Lc6��:�5��Avn$m���a��,uG����zcCю�Cp�2��l{�w���~��1�`
��P��~V��Ŀfx�N�������S�����p���/�~ʂx��t2x	;�gx�1�G|�+譫����<��;�����q�� �	�)?�(�)��<��!�no���!��51�bx�V�ŉ���G� h�q��p�E�*��+��U1�(u\�i���pdG��(g��Rr�f4�yO���..k��hp����ງ2'�X����>�.c��,�"����1��=�{�7+�p�;zz`ʜ\�P<�^jc<'���o�]�}3k�M�yW� ��@�^�@A���jX��b��4jC��g���ȔQ��}�.������O;ݸ��SU��Q���ET��%*qãPB	F[���*�Η�gorsa%ȋ�l�u����f��?X!a��ZrC�L<�ƌ ���_u) �s��@�^��+;�Ǿ�c8�z�3dAr��9<6�A���9S�oz�S�ʉ�=��]C��,R�>,@g�LG)��$-�e�}��[�J\`�>9�i��>&��v�� �B3�03�����nbKݾĆzt17pm\�C�ߧcK�`q�`,���'�_�ү1�ɂ��q�&�Y�$��5�*��:�혷�>�O]\��Ľ��3��lz\�)�thTJ誄�FT�d爻�����5�ԹƮ�"���=�
����L�3�~�5MICMA�@S�������ފ�l蘹��oLny�Q�x1��\��@+=��5���^����
�N�@�;�c��(r4:�>*/��xv	��&^=�dp��o����n�9�p��6��+\�AX����Q�Z�G
�.�vufZ����n+�%Aj�ݠR���t�NB���it�V˸�J�a�n�>|RĒQg2��+��E��xm�ň�w
��2���[K��6���L�q�c��H�{�+�x;ɍ�c��P���������!q{Ӂt]T1NS�X	�;�򯌯SJ���(ĪDy�����
��rG�|�*��a� a\Q xJ�
dl���S��ϵz<ϴ��1�4���M"��W�Q0��8�}=ݚ���!���%I=��f�T&����� |lC0��Q�Tz��I��4	1�4=�,�����)��~�/�Ku)�/-�cߏ�X�Z 1�hH�Cs���L<�^���4�s^��@�Q+�1�²x*P�mW\U�}Nӳ��{r�����]}�����Ttcܧ��Ō��C�t���eBo'�����k�Ě��n�؎굘�Vt��
���/��9����'�t�V���)�&�vpR���w�E���(�zӝ��7�\���.�@xڇ,D�8:����"Y�m�zb�R�敲/�Ud�a1J#DƝeZ��j<lL'8������[
�
�d�`�����\;�b&"�ud[�<7�p�F��D�'Y+U8��Td܁:H��b����48!DǼ|7�d�C��Gs����i��Ҹ���^1�"`쁮f� 1�*����+C��P��xZ>�d؟'P�9�P�D���fD����b}#o��%9ϴ�GLy�ǆk���b�.�EBi�8 F��.�Q����cƧ �Y�f�������T1�n�3�4�1�[�iKC���r�s��B���0�2e�S$T' r� ds,����o.�G����n�%�D���"�����*Fˣ33"8ob˳���0���<�Ͳ���y�_�ܷ�az�;�Q�{%̵�3��L^�<^��Y�I�|"�%���W(2%����A���F�����YH���/[��D�o�]��5��#;����nD�܁<Q1�i�S��MK!`���lrX��[�m_��M���	fC�`��j	�T��:�ʂf£��V���}���R�'�a���Ds,f�!��Q��lF�s��{�^��];0w�ߢ����-�G�� ����x�uv���# �ﻶ�arl0/Ҵ�<�	�4�q�f���o��U���q�T�C�ɔ<��Ȳ���X�2.�T�aȚ|[$��x������g3��~,�n����1)���ts���F�[��n۬�Is�c���z|'�b�7�]�*��I:�S����H�����z�ܜr�������U��'yT+�"H�� �A�FQR���^�����^0�L(�,Z1C�:;�SL�#�����ޯ �Uw��B��ܥ��T��[ ���k��\��tl�*$��&yz���+�A��ڃ��Mx$�+�Z�9#%��k7&�{���(*���C��Q��L�.ϳ;E*��V�^T�Z�����VT /Hs�L�'��(hXXث���/��,��I�s��o���mN�Ox��-��s��'E@��=8;d���g{޿ɏA�D�s��<�w�� �ڏ3�U݅h����Y� P�?M3d��$1����L	��fcr�}֮'����;��a�+�18�Q�H�f�Q�1��s gO���[�E��	����^�a|X��|�c�)�[���G]��Pp_�^ل$ܡ�ӂ����c��`��q�, ��8���W���:���8�ʞZ�UQ��k�+����02����9�Nޟ�g��C�TP*��E}�D
��pN��5�*-N�ީ}�z/C���V��]�Y}�\�m��}ŏR�]W�6��bې�mfX��&��V�ќ�����2l��9�Bb���Z�����n���E*#J�r��S7������S8�ܓ=&��'RIu���F��Di���M��O��8"��ƅD����IC��u�n��'�fs|��L?TmH��1�g�F��׶�{�u��Ť���V$�jD��;.�?\�o��݈�HW��P�+�bVK�;N��p=Dyj�4|�0���D�?��������~>5 �D�p�mȤXmo��M�6}�����uPeJ������(N��>뭻׾(������S5�M����@��$�1�s��dƮɋ �q;Bk/ښ�z��z��n{�+Ʈ�E:�@��
�2�Ls������o�{p���
,X-�����`�� <�7�W����l8�wQP�3p!�ǒ�}�QX/b%�:cި�����ڜǛ�.6+�@1>�'���¬�ʄ��2=��x+ϟ�y��K�ny~�ĝ�ʁ<V�N���2�8eH�Pŀ�z&N+P`JB� ̛�w�cU�]W����q$=%8Ϯ�1�	�]ɋϔ��(��s5�^��IUO�2�{�Gf;�{�>Юf'�`�����h�ǱM��b�q�3�P�?û�ٚ�Wn8v��+���LO�W70�f8M�w�㽘�&�u���P���i���7���}҇@�xV��c���k�v�7�?wI��&$?V~@g���ki|_�lG��$pdu���۴Oa�޵��S��rf=�\�9����1x�3ru��1�C8nCѸ�[��x�2���Lǫ�P�Kd�9�D۔+��k;��X��W����j2�@�H��g��f��B�f=^��s���^~����X�4=��n�i�m��$J1<�Z;�^=�z�q������8#��8*�X�ɋ�'p��S
�	M|N$�����h�q�F�wN�H��p�M������Abo/���ٟ��k��D�`�O|�6<��S�ᬺ7ڗz�Z���\v'v@�Gf�C�R�^vP�'eD��nf�N5?����W罵/�7����+��qm:�`�ɞs9}]z���K�4}�"ON��X��}�0�r�|�ja��,�ݫa��i����O*^ T���xH�y�{s(�d��x�:�����!��a�H��z@CQd�"|���b�9���^yQo�=����ه�{���8"ccJ�F�;nB���l�}�׳�d+�s�ђa������20�B��1ʡՈ{��߈������F�g����:T�b�>5��"9�7\���=�a o�<���S4}|�Ҁ^��H���� v�:>o��ֽ�ڵ9��<=��&�%���*M�9P� ^�F��Z&8_���^�U۞�v=љQ1�$P�C���zkM����r�i�x���ꑰo[�$��w_��4����*U�xҾį��r��Y��󲒄fr!b)�ַs$_'S�v�c6W�(��޼�(�R������yON�$?����C��3�p�(��eEؿ	d�2Đ'S��Ξ{g��<)bw&/��u��V�Q3�MN��\$ٴ�yy�^2}�LǕè�X�P��N��Dm�΂@{��S�[Ϸ��6�5�|��	͵Lf�}��X����T�g�w��|-O�ႢL��>u����;ME��S�<V���5��7�V�\�E�h���Xt�D���!�nKW1������j�N�~������t�=����^1|[4`��,�`C]۰6|W^{˽�nc���׏�uG�Q�, c��D��"�mGg���疳��w<
K�!}�Q��˛y���&���3��5%��R��{�DJ=���� �2Y����� s���iIxZ�'�0s&`z���T!i(p���aU��#:䣶�%ez�4õ���؇O��0�Z�bu��e�v ��mřh;@C��mc5���Q���Y7��Zܚ��˭�zK�e�P ���_L�5�fGrRM���dы9��6yS��۾im���9���`
	���M#^��fc]Ķik�f�YU{�v4���%c�e�*0�a�e���p��]'e%f���PU���a�eWG/]ˊ�u�'\V"�a�iס%Cr��qd�Z��2�ӗ(P�s�sqbD=�t7��3���_@���n�[���{	��v��B�']u��ۈ����٬R��Zƞ2q�yO2�t�{�����}�>���j�a��������ۃ�e�c٠�`��^Z���Z�T2q�u�n�^H�;i�vr
	�>�eu���+o��������)�؇�H�;��S�@v;������y�D{8��&�]є�������$�ח"�j�9��]�'5X���u��ui˰NK¥�]�ޭ0��Y�k��]iA�&�n\9��s���Z+/_
x���xe))�m��je��E��N���wIj�@ᰊ�y+�}"p���f�#m�V6p�9vxS�]4\�ަ�������Q.ehGv*\m^<�ZH
��EMF��5w�S����e�^�Sł�L^Z��8����8��B�.k��*�4\�0��92�c�
�C��{:���e���lkV�7PJ��78���'=F���Z�r+��9��tő7���,鯤��]��'U�\{s����$�/�{�0k� �S���1t8%����f=�T6E3U9]�G`���������ҷ\�!���wr�-�RF�[�'�b=ȬF���f�F�Ĺ��-n��ޔsu�.j�7am�Da�q�;�r`���ϝ�=s�?z~@�4(R�4�u)�
 �(
 ��(J�&�
JK�SAESH�)J�?`�P�	T44�
RSAIE4�F�����B�&�����*�F;���� ��"ҥR��@�P�RR�"�/r��C����������)����)�E)KJ1 ��41)CB�u(w߮|�s��w�\��c��5���[_�O��ߝGp�R��'���=��g�cE�F6�1�^5u��XJf|P�fuUD�	�SV���z=�$e}�I���6�joŏ���uz��X�� ����z�8�,�~�/K&&5O
71Xpm&�C/}</��os#'γ;���3f��^�_j��	�g	��+g��~0��a.�1����.�b�����Sc���)����ƅD��L��~P�f0���w�}#�2���Y$E[���S
cʴ`�tM�ohT;�O�w�^�>3��acnf7�Dm�C�8�x1_vLK�f%cѮ{���r�cuL��0&*w�Y���c��ꉳ�����N��|���(LnMq� w�S0Q@'1����(mn����{��Q��G�9TTYviת:�:���`�j	���d��W��~�Mt�ҫ1�D�w���'%�����>�o��Ш�i�/39��u@R\��	7�t��mo�]峅0D�:`�R:�{�_q&�^[�g^E��[�$�^z�,mD�cs�Pw3Nc�<&�W�_I�_U�ɝ�Ǐ��{�{G���QX�|�L�(�`��P��C�08�<��WS��6�l2�Q��j*=���p�9�A� ���6k2�^��,��a�#\z@�H��U� ��2=�x��	�cj�߳yyz6,��(�4	1l��Uzb��aAת���݀h��~^�I��g�Lï������\"ѢX�4.������_����{�s�Bv�8p��G�k(F�70�f8~^�/^�fz���xo�:��f:��4X!��+�М+OG��+��0*��y;�>�]Q��Ty���욀�������X�?�޽���yVx�f*��c��Q�'=;�ܽ��\}���F+�+��I�����ur�;	�E �yDU��VS��ܭ�	]Z0;�%�O�)�g�rAĥ�ʜ���U�s�v���t(��V�]��vJJ�E'���fG�Y��7;;��G�'�Y�e��U��Cߣ%��uo��S���GU,�����1�OCxjױԲ�E��k8O�*�i�w|v���w��o�<<+:lS;�_q�U1�5�[I�7Hn�?��n~�%��a���B*8���xb�O���ɇ�
�E��gZ�{����wQQ[+.躄5�8\�b��bi�7�}4<��;��]�>��@�5̉.x�r�w��b'�pY�^�CtzN��Z���� �>ӡ�<�*p(H�'��{�(���V�ܕ�d�nH�1��$OL-4JJ@�����F@��Ԝ	u7�ܶ=�I�y���}�c�&8-8jc��B������=�w5ޠ|�^�&&#xz���0CP�	�D�@�ֻ������sQ=j�KVh�9�?�-�sˬ<���t�/<(���k!��_���}����Al�U�.n�)��퇕�9�n�Yڌ�k�.�`�JI�q&����f�䟥����Oaj�s�c��@s��Cdk�@�:��e��#ϙ�W3F�x��@	��F�Dq��"���mg?{2g��{� S>2LRɎەF�X���"�}���{Q�u�����0{fT�B�'Cfp�y�Ei�w���ep�S��w�p!^6�C1s�E�&3��U
nu�0���k.<|=���c��C�{<=p�����{q2�D����G�zc�������z4����j����������֨*g*��Aۡr�~��������`��4wƬƳ_y�.SjX�S'ޞV�'b}�3���/8��dI�0{�������N��Q�����A3�~���yӨH� �&�D�O��W1�)�ٓ쑯�\�nM�������٫96�~>w.5���Vu����+d6S����w��"!藤���ԃthe���M��e.�X��+��0�>�����l���*�f-���cb\�`�<�`�j�m{W�Ώ��D�f����͏;�PX �Zj	�� ER��B3���ܽ~�'�_���$ �ޘy	��x=�0*6
�S���5���~R��#�5��LLg�S�~ /Yr�K��}4��x��7�,uCG�ǲ�Q<V5P���1L� 3sA���_�\_�LO��!�Lh�s��5<)�8��G��͜���2j{��~��I��>��uJr��ڦ�ł;\�����u�/=�����=s��φ�w�Ev��������� ;�;���$�|� c��Q�P���Q��
gK�1�Q*=V��z�������55�hU��t��Z:�W/���PvOߨ��ٿb_�k��1G�i=�-���]���h�8{�o#ƅ�}ar{F�l�ҝ^;t��{�n����K��&�Q�yӯk*B@���ۭ�e�]m0I:b�#�>�����x+�#+n��5�uœ�zcsަ6�H�c ������f�����Dᡜ@:^9��x���}��f;s�*��W83�+�)�5��Ɗ:ϑ�;�^< �<z@�uPbT���<7מ��7��l�O�>�粄UϺ��Q��n�c�Q���1ܤ�;�*xe���j���k�sF�%�#c�۪��P�w��Fx7{k�s����4<���7(X/B�}n���`MC��V��iz|��81/&/������Q�X�fX�zĲ潈W����c �Z��"|S1�Q�T&k��]֚��~q"7ä�0i��F�Q@�GY�y�}9������.;	90���s0����|�����g+
��cx���3R��l��7��W�SEMb륄Q�.�ɇ']u^<����찾aXR��T[�gN�����E\��s.�L�R0���(0���]�}�����ֳ�P��E9챎c��C�B>�dO9b*5���D�V+�b�\��׺<�^�˚�q��]� &�1]r���s
X"WK�hQ�=~9J{{���meF�c���v�ɍ�x�<(o��,�ڐ���v����\�u���<�a�7�_aa&*�D��Vh�Je7��n��}��s>�ba��V@z|8�UC��\<,E����͓�Q�2��W��c�i�5���[Q�@<rN��p=�Vx �>u��[�f4�8^����3�:�e����0r@�\UAW��>�T�w�{�̾5|5�6+K�b��8f���wL���������Lȉ+�*4�^*�v낟�8+�Z<-yT�S��r���E[��	�@�(<P�{M��}f���8�øm��9���5�E�г�^��+7z ��͜�FG3݆���*s;����3�]GP:�=Cpibg\���7s�E���l�>N�Z;��q5Z��~�7���D��p#��*p(H�y��dì�5�QNy�zl���H����d�sHn) ��D�,g�W�?D�0y=��zF@�eɏ?H�M�b}��&/�+M|jc��)��m����_�;��=�����M��������6� 0�1���Tvy��(�g��o��ʬG^Loja��:�1p�O� 6H�e��G�g�S��B�t�&��
j��x�[(=�����PQ�v��w�=t��~�vx{��a�ѐrb��nd0��J����IN��ߪϙ��O�a����"�E�Q3�3:h<��2�獦�GH�{{���{��PO"��1�N	���q�zf�����ݺ�Q��w��zݟ"Ǵ�q�i���,vw�c��.-���K>�0%d���5�ά��l]��˵tk��0�ꗰo��u�4a��a�,���w��܀�Em�&_*��R���Laf�A�b>ĳ�G�'��l�ӧ[�����+XL�\�j�u':P�B��hcDfڨ��U�3����i��f0K H�>��^s
�TZ,R1@�j'�+���{\Z��Mi�d5 hC$����Q��B7�3���D�f�<��1�{6*;���e� 4@A2@e���{��]nsxwW�}>�������a���E�Q/9��\�`��	�^��#�!�s�`��҉���:�� +H��3�t!~��]W0#Ԯ��K`�"�i9�,L{� r�E����+wپ�	������DO���,)1��{����:�B��m����q&:X���|�aT[�ఙ˨L�z��I�nϳ{/3�v�i�az���#��U@��tl^����>�+�8x'<���pT��C�c��|7��'$T��qG{��;������k�OjU�iY��Y��+�rR>F��ظhӰ���C\��|�eF����������<��67b�
�VY���dl�����w(p�y�Z��CO������&�w&Q��agG�*�����v��d�w���_l�4;�>	���1�{�G�������MM�k1�&+aӗH����-R�^8(wb�".s�&�����^��C*YU�󟮺�Q����53ˆ~3���/L�{=�^�ǣ�bw'�q ��1��B�	9Ɓ�1�r�7P�j�-��x�6.��	̚F�D�Pz@�qU��ǃ֞��F������"�<'�pE��{��9���)��J��<��T�u��<�4�n�f3�ScZ����Z:�*�y��k��?U�0]���еO��ͭJ�Qf6 �Vwi�X5W����WU:l�Z��������A"B�k9|b	^�,�A"Ca��&�;ܢ�--���fW5�w�������}�;?��TĢ��R ��p�A����REzZI�M�������^�$HoRUsVu���Ee����=q��Щsn���(�62�6��d�E��f���a�-�]����T�TA"C���n}���Y�����2D$H��E���p��k#��I��"x���Y�siXu�\��(Wc��$H|�����oQPٌ{Z�av2�z�ƉRV�z-��-����_)(ǟ��H���g]�q\��R������H��4K�۰y_%1D`z�8`�I��*��j�K.�UxW����g�S� �!��WL�,a��c�}�/ܥ+���1=��s��G>Y�^Q���??���M;L�+9�J� �!�qf�xt��v�������%>�0��v�XX�'���vw�����StLI�8�J�'ͅ��ס���A"Cd�T�WCٿ�y��	�g�Y�>�^Rx*uXm�"D�e\�H���rJ���b���9�k���h�,��by�?��H�!��,�ƒ��o�L�D�%�A��c0zf��i�9kx	�������v8kE������{����H$HW����*MӿtG�6���>�9�Gfٯ+��J,��]C>��ƪ=��#j��v����X�D��	ϒe��[�*�RZ�I8w�W	���ˁZK���j�zGw�i�MS�i�Lp2�l���*q�
)I�	0����2�;��l�ˀ֣���U���i�f��
�ꍸ�H���t�bj���J�m[�q�N�E��j�&�n��(�gGfVߢ�{� ��&�%I$H���{F�}{g���0e�ٶ�!�7�SlTdc}y�&%��ȴh�c��_���Ȏ���qײ�L��rE8P��n�