BZh91AY&SY�ɣ�ݸ��`xg����߰����   bF��   �J��*   ���l4��EH IJ�@�  �4    �%@�j�P)Ta�*��fU�(@�bvm��F��A�I��[i!F�P)l��5����M��5�h��)�1%�6�@�Z(�ZD   ` |�O@5�a����*%SB�X�l4m�mg0 �W�
�dkp0 h�.5GJ ��.�� �p E� P6�Z��icZ7���*��J%�C� U�ЦիM�M�4P+'c�-h���U/��ˣ2ATh��[6ƴ� �K�tP ����_>�B��6�P �vp���TS<�{�]�F���GW%���)v��}��^�ڴ�J�uW�o��v�Pr�;x��\��	�y�{ʛlk3��ހ��l�{:x{U���ݛ]ZhL�:�Ckm����)F{�6����ea�o�:=+^���g��{n��gk�ﯻ����U��<w`��W�G^}�_j�b���;{��k�Svۧ�;�=}��+h>���T�O�:�]>����U]�L;��%�EP45���T����[ڭwY�<���[̙s�;�U����}�|�XvuZ��{OJ���}7i�l(�W������-��m����[{�wF�������]wv���˹�[U����5VŰ��>j�UUF��M>���&�m)Ц�ƹ[)�+�upR��շ:�����gK�K��Vj�ή�Tn����Ҩ=�����U˶Qq�tWN���K���@VZel2��>�UUJ3�L��¨N�tK�f��W��֎��.�v2�M5ܻ:��]��
�.u�mVNy�x�(i�t���m���oxuR=Zx����wJ@�VZ�5�B��o��P� �����n�p���u��ε��;8 �R�\ݞ� x��:̹ ѷ5�U�v)X�vՕh��{��"=����k]t݈�h=���ͅS_zP�U(n��iB� �n�p��anr�rQus�P��jr�A*�G����U��.ݠ۝wk[:����Ngm(�WF�hd-aTM����B��Pg�}�
���P
v��3]h7Fh\�G�@L��v[����M�Y�5D�Wn/gz���a�����9R���Y�0h�w�R��U>���)����GR.���P��ˎ���u��j���t���Y�ct��M�g9V���j���U]]��i���( (     P � ʔ�C# �!�M& 4�T�1%QHh��0#�24����4�H�ML&��a42d� S�$�Q��0��	��0��
D�����Ț��=A�'����SH��)%@�4 �@h �����#��J��_䬕y�|j�$[������=�����>��*��U�<�G� 
�
����P [�~O֊*��o���}���W���������?��_�/�AEd�<����QU�	�H
.�������	�?�!���$� �������아��J�+	U��a)��!�0��S	a%0��0��U0��!+a%0��Ja%a)��0�XJa�E|J�!��"���C	L%0C�%VXJa+	XJ�0�	�a+�J�0�!�aC	XJ�0�#	�J�F���0��V�C	]#	XJ�+	^�V����%a%0�%!)�0��V��"����#	XF���>#	K%a+a+	L!��%a"�V�C0��Q�J�S	XC�0�%0��)����	T�)���W�a)��!�Ea���C��Ja+���+�!�V���Eae�a%a)��%>%Va+	L%a)��"���+	XJa+aH�Ua�+	F�Ca+a+	L!�a'H�0�	L%W���%0�!���"����Ua)d�Q�H>%P�WIUUX@:AU��S	J�S��UL"���S����E;	D�%C��N�U;	�% �!G�0��J�0�Tp��US	J��P0�T� ���U)����
��"�`B/a
�"t�a) �(VJ�%� J��0�L ����(�"���%���@�%�T;T�$Ga(a"'a=��a)T�)L �U_��
8��J!�J�a
��(v��J�a ��*�������:	���Q;	�$W��^B{T�$C��a)T�QL%R����UP�"�	D�$S���Q;	�%����C���T6�aF�L%
�*��*��T0�Ua(V�a(V�a*�JJ0�UaT�)L%(�S	A	CU{Q;	�!��N�T;	D�!�%B	�$P�"�XB���)L%R�EU0�T�%U)EP�a0�S	J��a��U0�Ua
��a0�SIT�0��%*�J���	T��aV+�H/a0B'a*�(v��Ha�a�! �L ��T�
aT�L��������;	D�a��a*��(a*��!C	JVS	E=%R�E�ER���0�+�0�SU0��aXJ�!)Ta�%V�Ca!�JY*���Ja)��%0�XEa)	��%0��C	U�VXC	L!�0��+	J�UzJa!!���	L!���&�C	L%0��+	L'�0��Ja)�VXEa�0��)��a)��L,�S	L%<%0�	L%0��S����p�a*���Ja"�������J�+a"��a)���Ja+�0��+:C�!��-XJVXA����a*�C	XN��a+	L#�0�#a+	XJ�0�%a*�a*���Ja)��Ĭ%B0��Sa!�����S	U��+a!����S	XJa)�xF�J�%+��%a+�0�%0���#�aF�a����a+	��"��H0�a*�!��#	�a)�Va!�%Vda�0�0��V��	:��Oi����~wް9�$����K�w�b�_,�W�#�uX�2��$�2nQ���n�Z{�^�V�v�cy�.ǔ�.�^2�մm���Ɋ������b��Hճx�Y(�S`��f�W�\�R�+�J��sJxa�J��q�u;����57tl�A�LDJh	����w;t�5���x wd^bL=���6N^u+$<f��F����Wr�E����إ.f-J�KD������ksfL8,�z}X�)ԗ/wՖ�Օv��X�M�K��e(uʦj���.�^O�$[bj:eDk2�%R���m��V��ݪ$]������n�r���m�"���L#-(XFS.�J'p�����ה6�i�VQ�ʷ�ǳw��eݭ��/$n�eܛ,�9bjA�]�b�	5�	�b�i��ֈ���y|��w;i��54Ya��XLbꌠY���]�P���4E��T]!FBѺ;��^nug:zNi�&a p����t�*/�'�6�2l�$%L��w���w	}o[
�s��(�ʗZ�&f��Q��.^#�R"�I���U�uh�ae�{U�=�n�nGI)#�]2cʶ��
Fh��Tp���.ۋQє�k4�dD�����t%X��5O2���5Y���W�Yn`�N٫���a�s��u���o^��a�w{4�;X�\ο��Jd-U�o͉G
�V:�^J�_�oʼ{0�(4*t���g5Ϻo_h�H�$�JŴ{����K�J-@��9�'HֻȬm��b"���|�j�d��/�Ǖv��/ez5+q^	���u.��^u1V�{�;\,I҆u�Ɋ�(F��c7����T%�{�Т����&+�,��*�u	(���1�պn�og:M-�[4��-��.ٯ��&����d��2��z4�ݫ��M*Lj�&�ô3q*��!P��FK��y��MY��0+�+���݋�+.	uwz��#vC:pa��vG4KD��N5:Ƹ�:�κ������5��N�j�ZJV�+Y�NPɁnĴ�<`�ڝ���9i�JeL5n��F��Z1n�E�T����e(�c0�惼�ܱ���{9�IX�E���5���ջ���"ۻv.�h�rwv�I=2�.�����ީU�3���CY��:e�b;Cb�q ���o���4%��m#Ef_k��9g5�9�Y�{�mo:���Z�X���4�e���и2-���Ht�]m�e�s5ն5m��N��o��AQ�"6ɼ�!�M��yyB�&�����[�T$9S%U��_Z���t,Ǽ�,��[NZ�Z�Kp�7��"�WwOU���{u&�mJqټ�ms��v�j�>�v���<!���Kc�T#vB�LК��/\���ܤr��<��{U(/r�f˛Pq��d��q�q�R�.��n�R�T�(�d��<xC˄��@�7]V��r�k��ب���5dM��QWchf�s��@��u(�-b��E	�X��Z���2-6���Um�fX�&�V�i-G�D�w�;�A�:���t���x܆D2S���m̊�����I�쬱�i�;W�ݜ8U�j����+�	���{Y���%ݤ�����d�n�r����ߑ ����}tF<�$��Y$���Hh��Y�J{B��6��A-�f�:�/��6���at����!U�j�F���UJ��}[y��}S��sQ��qЌ|��{{h,]�3*Tf�V���h�n�/ia*�US��6U���{eHoj�b�3瘾K�r���K�5+c���å���ճ2Ӿ[�*�L�Z�M�I4�\&싥*�F8��չ�{�XqB('j�YqS'!2��"!aM��C+3dƮ��v���`x"�o6oP�V�W��몥_}b�8q��M�j�50ݸV<8��=v��H��N��t�{+O�y/��/gW]�q#�ï�E^
�,F*Iq���$R�sUK5�Qh�/j�\<W����Z����M�Ѯ�Y�Q0�-�����mJ���C�EV0��4��`�%�YF��r�f�E��t0㱙�^�^��#�s^�t��
oi@�e��H!eU^��*��S�PmP�D�Z��p0��׶GDݫ9�R�b]�+3�u8�o.p��T��[E��휹.�[wa�bct�A���i.˛�tTyC�;݌�Iƚ�i�w�	����/D6ڈ��[�=3/7P̃uQ���L�v~��9��g
��ʹ�=�ѣ�!7v"��+r�V�}�Mu	���l��	����᝚��YlݣKّ�j[��1�`�\c3]chm%��oP�	�	㒻f��Ĉ؂��r�dʧ�>UV�+xMЏ/iѧ*�£�L���ڻ�XF�����}��T[1\Bv������Dr��g9l�p��M�(�j�c��,C������LFyu����E�|��O*U�i�,�e�k*:��sm���
�P�'�A�w�h�Ӳ����������Ž�ֵ:����j�Tī��z�0�I)����1��iТ��3��{.�f!���,��ɪÉ��j,/k16��fL�M�:����ֲ�J�N�V�-�Ԫ�)��a�h�40�Z�f�,��2�+���RJJ�|��#lҳ7vٻ�p�۽�GK;5/\���Ch���f:Y	��W��ll�YtgU"u��f�2Ph�x��Kn<VW�i�ǣL�uv��1�cEi���ʀ�͎��^�!���[�*�bkr�cB�z�)5�o)��E���逊�Pc�\YUJf��M Ә�]��Ҁv�c5z��"�<���6�NM��k��4���{[W�o��VXhQG3e�&6��Q��Ub�V�l�ԥ!\�X��{������VYq[��Y�ȡ�9�Z���9�K�)
�/+%�����+YۘLwҪ���M]u��-�-��pm����!�*���rŶa��5����:��M�׃M Rf���r��4�z�P��Y�A�&��<+��Bޞ�vF��T�u�a�����C��GQIsVAN&��TOM�Y��t2���I4H�%�����-hf���re�Q˸©+4:�����ywe�B�82y�!����r�ӆ���V�F쨰6��c��*�{Oz�6���u$���6��n%ג��:��d.��V{.��疛@ˤKͺTq�&�^Ă�5\:�8�!k,���i�-��2�b�2�����U1��םfɒ��M�q��nդF�J�a��`ӧ�5�̘�B[2)Q�m!��W�Nܻ���72�1b���͙SJ���'^����ɀ�U��2������¬�\��ZV���0�Y.��/L%Fff��+�u:��b��)���I+�uxt�̏*�ݷNcH�m^cF�B�=�%��^]
V�uR�X*��w��d�l��K�R�.���	��ʽ���ѤѸ��Y��s7),B��*��2�b�h�؍o���#2���J�A&��3��kin	�L��n�
��,��lVYՍ��ȫfnA0f��,"�sЪ�f�S/oyd��A3��ڼ�#��0��İ�p�,GTV*�Mճ��X��m�n�cddr������ԧw[*+��j�n�Rn��Q�n٪-�N6W��!�&f����x�����������1G���VAyD���"�ީ�t�:t��Z�e3�f�Zx�A��D�eɱh��KKvń�ĸ`�3�M����rӵ.��#�%��μ�7�e*
TӚ�RLԲ-���q*�eJ�$�qy4�Sl�&T2�o,���>j��'8�[�uD�W�l��5�
��[ӻ�̡q@�ĥ�3i��4��ɸ��%]�y��	l�5��Ȋ��+�a��Q[�2]�==Skl�ЩM��h��v�Y�%�s��9P�J�%'��%U7m��+�Vp*�����v,Ȯ��q�ƜE���ݍ��Uk ��WYE�	fl�j ��F�9uiշGQ����u|��J ��e>!+����)�4�&�9��%u�B���.��5Z#%�n3�b�ڮ�Ǥ���2,J�7d���t[��x�s40�k\
m��\�w�PZ�U�Sͽ��㽗�p2��"��H�X2	�)�ڹ�:��h>AK�\��1���*�/*\U�t�;P�J�wV�A3h:v`,5 .c)�Q�,�n���gT�skp#���[�l��b��.U8)*u��Кܧ�KU�m�[�i�m�64D;V7]E��S.	���C�L&M�p#6K5vn	�D��H2@��UM�d���PI�fi��0(óp%)�te��ٳ����$ܔ��r�q��AS�4:��PV�&���+W�cg0J8�D^�a��6,�&���AMܷ���or�K5�WNf^-G�.�!��9�B��P����
�}�N�]���2��7*�!�O"�F��JM��o5}j�leW�RN
[1M�8^[�8fY�8��N�7�2	��!�sM��qfn��z��­����w4^mѽ��)��q��OYӐ���&7*b�vѬ�ӱ��G�lQ{-�%��va�smj߬IV�����3 n��DGB��l�e�4�/p���L�UCn��T���X��K�X0$km"5�M�3�S�	ǌ�a�^�)�X���\��a3t�h!'���$��[��a��#S�Ȇ��5��B�͓wJ�j�b�u�=JiJ���4�ꔗ/l�VJ�TS�A��G0+�J�h�S���'G/0���j�����.�m��Z�����P*0�B�� KM�i%�1���V֚`�n�nZvjΓ{���\j�c�T�75luYI�uV��ܣr�im���0���j�e�;�7[#�R7�i�!Ja�7����얊�͗.���0�n��+4�n��j�NTa�8f��XۋJ�8M�EZ6��uU���/J ѡ4[���\����"��n(�Ui�EG�E;�����7��cI��Fk&������T�K�,^C/Uޗ���2�`�8�̧��W@��(�������*s�Wc2[��S��j̚st%OoY��*��*�3�Mo
���iѺ���C�+���L��ҵ@m'�F]��Q�ái���˻�$��R�����B�1!k]��Z�%Y�a{"X��W�V��p��U����ӫ��%�Z*)J
J�fe@�,TE�wI�RG$\�i�T��f$���E�)X�H��M�R��y�q�U��[,�El�4f��0�S�b�غcv
�u�Qa��з&+� �L�]-Re��Ul�L�ڇ��F8D j��o61yjj�:l�V�I�:�Y[WWh^Qv����.�'��&ed+Zl!wN�G1��ն�,J�,�fZ(��~¨��c�pJ�C�J��*f&:�N������^7V�f1.��\2�3��7Uz����^���P�L�e)n�t��e�8�&�eV#��J���Hb�o(FR&�����Y$l���/"E��rMڄ�+fʨ衖�ݛ�ܼ~�Lf�QR��+&��T�y��b�ۻ劎f��'�B%m��nn�V���iE��gc�1��ک�s��d����^:��/d1��+�z"�!|��7AbU��^�a�wt�J�<ӏhN۵����2���i�&�*�Ub�7n�$ZpZ�M^U@�3w��;�xk�J���
���Ƀn�kV�X�zV�nËk�W���%e�n��ٷN�v�(:d��EH�哑���÷&�2�n�Y�4e��s-N��%aZbV�Ѡj�B��^��|j������l�l#�z.���X��$-�~U�-p���kq((aT����5aGθf1��Q����Hf
^x}�[��c,��aB(&��
�6�p��&����5���FR	`�Cd�u���O)��1hŢ����-�n���-h�t1!x�g�F�%}��U�!M�
,(�E�_�2(RC���9�C<�ˁ�1X�E]�$�@ߖ�,��?j pr"\hnAo���B�
D����.��c��x;��c��`���ŏ��2؉�\�J�����B
�Ix���Bg0b��;�F�Hc^d }��*�L"��7�M���[������S��^��$
����<$h�C8I�q�{~�xr���%����2DO���b���AC����l*C{¢���\X��Z�q�8�0<����c�(4�,1���3P�C
׉M{Hք.н�!XN�Zc3�g�,l�m�`jD6:�g�*=���V�L+��XS�|)��ãB϶�uhp�5�l��(
*�<��j��P[ �H9���`��Nx�Ň_z�$����+��ō�	T/H���{H�﯃c"ތ�/@��=�pcD74#C�lv����*��Ƞ��0P���/�&Go�w��$�}��0W0�� N���g�������1ع�g
����p��M��ظ�B
,k#x�M�LY�wyׯٺ.�,�����<�uy,�uh7^��]���9��:�1��h���
��LfP��u�X!���~���}��	pj�(5pH�puh塤1`I����<	X��PR��r���Z���%�x
ፌ07�X)X��j�bC�PZ����óA��^�""��Z1�S<`j�-�4�n�`��8"�%�X&!C��X�~��)������<��b`�푻��V1%�`]HC�U	�=Bk�-��

�1LY�j�z+��C�	���G����B8!��fLm{6�A"�;HU�iy�7��J��A�"�!Ɍ�@���a=~�V����1C�`���ƛx3=kְne��A�0&G^��$a*=s��C&z���j�z������%{/C�ؾ�����#a^�4�q�-�� �����e
���D;PO���oa���]��8<�hA���	���Q��	`�B�¤~�'[��Ǯ\���I���������П����������D���u�
���m��m�A$��M<Ҟ"�m��6�m�m��a��m���e�m�޶���۶U�U�껻���Wy��W��E���sr�\�US���'��$�9 ;/!�dU/�yc�(�Da�'pt�G	vt��.��dV���y3V�Z�ԑ�`�f��4��j4븬&��\\��0�ɰ��m~n;��6���ط�l���T�%�9[�Qe�6�S������Y�
=V���I�vd���FM)@o1�Ǒq'"�qM��G6�&�����m65���ZѧaMI²�䨊�o���uǱ�&�(��{�ㅤ�B�"�])��h0�9��Sw@�Y�D��n��*L�'����;�r$�хUu�.�,u�}�r��̤��-�5y��.��WGbά�S;y�7h���)��P�)��"�LZ��8	���wW��vDP�Y���7;t�q:]��6^[�\Ȁ��	���θ	WV���v�,h���Q3a��p�,壷�/��i�w�}��y�e��.��"���'��fp�i-��I'[�]Rf��{oldZ��I]��}�d�1�6����M�T�t�*�y��ەx�!=�6�mm��]y��LV�n����W�=Җ}�]Qv�l�EC�$��Р:޲"S��aۑQ���*p��tsZ�i����FM�b�"�R+d�i�I�^hFv�vC;*4ط�$6��u�����^�t�ӷч�-z78_W!T2fK�Q&d������X
�;.�]����@v_!��Ȍ��[X(n).�8 ����Z*�ܘO:�UB(��+g:���}�&Q�R����DS՛��΃˩��U�o�B^��}Ƒ�R�"�vӅp
��Z��Z�%�*U�\�=j��1���㾿~�.'��w-L���村4<�i@�7vTeTa��J�c���m)lr1�}{�q�r���i�:SFM���Um2F�rd�sd�ZU�:g5Y.�Yy��<�OI��a��gV^�O(�p����9���]�r�n��)���iV�d��G���5p�ov�����ZD���V�Ew�.�"��:�	���޳���m�ܻ	��1d�D��E㘨0��Ц�{9�8���j�U�[D�������'��Y���x; � �ù}�up��tB��S���}b��<�:���֦唛�14n3v2s7]�x�bL�ӻ�*�9��9��qU���J�L(��rh|��	Qm�<��O8}aL�V�^��eV�᪦RB��^�2�M�傒M�ː�-�D�)�ϳ.�2̓	
VчO+��TLc-)Sp�������;.�zu���J�.a�e��,��CAvS�g��Z5���;Ň���fKV�L�y̐�mH:�<��Z���m�ɍ�؝5��Ng*	5P/[/�[f,�v�gCڻ�M����^+秦]��e}R�QW��EXg�йO+������uD�V�@�귭�N��ڄ�T�V�ټ�w�BZ*!
�,x���m@Ğ�w�M�dI;7$xk�x�<�����Z֜�qu�!g���\��]E��nV���sv��FZ����zMY�k�j	��d�YY�ȮY::�W\�y��H�X��S��x�.�X�f:�Ub)֍�(F�=-�W����uMх��wHJ����,�6��=��N`�LDB�iY���n�s�I
���}��
g4�F`�fFC�U�P����M��k�5[Cxd�QAj�u|����*(���-��DZ�����&��L�j^`W�s�E�v��;�W�2�%���P.�CjrwCy�}H�ǽU[�C�g+�h�v:�s2�����,i�O�&�p�Nd�E���y3�D�,1f.d(�V��"����tA-��J�1�q���e�HE��u��.g�Ǌ�)���^_		R�.��uյ�gc��pm*l�R�NmP��EC��u����k�]��|�Cս�����p�����oN�u�ӹ7r������\�[/�MƻQ�Xl=���؎�X[f��Y(-f��njN�O_i���56�S�K2\�+�����0>U7��oj�L���
�u%�M¢V���)[y��RM֎�w2U}W2KS<�C���U��0Xfn!.������JwC���T�O�U��!@Z�.�&��^�H�e^Ͱ�wb�-V�c�5�<J,]Y@�Z�<�ʚ�v+�K#�ŉ�����m�K�m�����v�D���D��2�ƨL:�ٶۼ��
]��8�VS�t4�eڲ�h#�K.�@��뾷�猴��Y��=Y��'h�u7Kۧq�&�yC�K'N�qfU�j::��Ѩ�Z\ʙ[¸��g�To^�N�!K��ڻd��#$�N��^�Q8�MSm�J��Y��*�X|�N�)<�&�Ǥ�9wop��xʄ��6�䂕Va��ǬZ�fSѻ���LJ�*h�7�Q����s�PfH"�����%x��uu��n@7�����^���{Y�3-�inV貹���;�T7��`�6&]�F�^��K��J�9���bE�x�Q�6{"P���J�xN���Dou\F�\�v��X
؞�����đ7me�C1Z:�c]�oF���tm�{:��an*�:!8&�D��'���nL�+��[��W=�&�M@�����d�<�4�+`��jص�
C.u�ur�e�kmN���F�Q�.�8��CVZ"q�]��\�r�Kx�dOu-��Rh�ؑwG�:�{X��c�Lb�͙�����V�s2����cV����4YˆIN����,n.J��Y��Y��Ǖ��6��ڽ2�&sa��b[�켔d< �Q	m�`�34�mQ�of�ry��6�oLaK��|B�o
yk�ڈp���Y3;@�D5I�joj�;U��.�4����NL[��۰��w�t�V+ۇ�����H��u�{�a+;|fc����+��]��W�e��XW��IB�z��5�i�k�҆���]�nU�{�m �Y�ͷ�h;��86�۪�S� �[W�O*d�Rz�c7���%���[{e��\��lc{nJҠ���ur��;U�\�����Ǎv�%_n,OO�Ѻ���U�g�161N��
��Z�܉նa(t[Y���:�%FUkǙ�W��B�ʗs���R�K:�^\�ҍ쨥�5��`�X�q��:���ذ��z�J�[�*77{6�U��e*���a����0�5��,X�86%֤j��U�nv�W��s6�ͫk�K��17+��i�1a4U\�V*�\�a3J>�h���\�T�����wV����E(܁�]���E͗t���)��ˏi��f���W%&]���2\�R��ŵ�W��egs��Bis���%�+e8����y�X�}�u4m�WU���w5�0�*���e�^�5w�\˜S$��=R�!h)9����2�P��ec�X�iu��vgh!�aY�9���5WC7g����/\�&�2N��%�ֆ����j�'Y�äW���p�p�:֧b�����"��i�<��=��Jʼ��,u�e�W�dѭ
Rf�<�a1��i]���H�̻ܼi����]�@j]m�QUZ*�ޞ�j{ɚ��z���;I7�{5�«N.x��+2˻lKy�:�2�[�S�F�x�ah]�,ګ��gVN��W�Oe�W��rG3[�_u�z���y�^v��������&�U}h��$LΔxKVՔ�qL\1�3�JѬ��lTuM���b�u�K��1�=�}]��y�z�8Rf�+�ȹ)5x6�*2Hշ)[��j���v.�j��rɻ�3���:I�3����i��x�53�>��oY�W��Es=P\�'M�}C{�)�G��s(�b5W�ܮ'L������G��鳵�v������P۾7tVe�=�υRA���^v�Y��n�c޾�x���EfRzS��q[��I���UJ9�,�r����݋7�����6�	��)�u^����p���3�gJ�N;t�H1/�QG',�rr�彝�	�5�I�YS���[�6����(!�a�`�a�	&M+;$��5�&���z��y1�~m+���[8�$o[�.��͕��W9��evJV����)N�7���dfl�u���8�F4�NÍ�m�X+~��M�Ƭ4����6oQ����SWg-�ť5��AWSy��\�P�ժ�ʽ`��Co���'v��{+:�1-+>��Je嫵Fov(ma �.�7Y;//Caf��ʸ<�N�
�wKj��{�ho�Y�g��Hj����v�b�6��� ��}�9M���ܷ��=�:Օ�E�r5ą�N��UCm�Q�r���LDm�sE�ujC��+N�3JN�hO��7�d+���}x�z�A��dp2��1ue��	���f�CQVC�h;��䁺���KV#n�	/4*<2k��p�5LU<��I�`�ԃ$�Ȣ�EJ��V��u6�b=��'�*��S�W��p��a�k�+I��9,��q�\4e[{��Z�+3�LJx�D�$�u���EJDU�gIN��hIbl�Ĝ�'aU�,�X���򪪪�_sum�L���"�ZZ�%n�����[��gV�m�Q.����v]��\.෱�K7�,��6͐�m�3��͢�&�S|薩�ξ[�ۙ�[={��G,)x�"/)�klj�����in�ݲ�-�[p��&gm�l�O-VQQB36�p��v+��Ӥ�M�wVV��
EY���gXc:����᧷�g[/.�ʝp�Co��塻�si��Toͨ�0���.�\,6N�WU����L0x;CWo�0V��q�]������gM6�M�V�g6��T1�S/]�:�Ƅ�F��;�(۹����h��U�ޗj�-�vn)Ų�,M]RU���[�ټ�Æ������e�J��P'�M����w�E�5uD�j�R��e��B�أ�[�QE:=�
�wmW-p>+lnfAj��,�R��0Q�d��2��;;oh�������ZGf�Ͷɘa��3�WP�f�Ԫ*5��KY�,.�N���+��(�;g�+�1��Ku"�4�ӯ��ˬ���JvvTj���[O*L��D������GR�'	��a�{yp�|u��͂R��EHβ(!)��=I�˙���W���ѩ�L�!Y\����[�9��6=\�u#V��D%�C����n��+�L��wp.Q�A۵ƾ����>�*938]�y�*��$���>u�:�Q�D1�n.��
�nAC��{jA�(mKu��#|w ��G���X����fQ��&�ǖ+�����
[X����(�K>�Z����é�T�����=����ٟ����f"�λq:�PMM��df,���W+{G��L��I^�z)�.�"��C.�j6������}NoD����%u{N�ID�u5���nQ�zu���q)��[��i�.�u�Y���u�a�(����&wC��n�[�Z��Ec��m���ֺ���������E˪V�W�Y���W�N�pf�ǨSĊTNa���fa�mg_���G�lݚiN�cN=����Ү���Kan'H<����g*��xW[�vl,�rQ#
&�ϋQI��2oTދŘ�����#��U�G���-5�fi��w��`�P��6㻾u�|��8±{cJ��Mak��n�J�T�A%v��0��x�N�z��r��v��EŚ��'N8;�ooCOh���T�M�����1X���t$���-i��r��m^�ZMDV�"�x[i��m��a�z�:��M��m��n(j��"-�x��um>q�:�o:ǯ�ƭ���󨏝q�x[�N�բ����DDz�^�[�׫Dq�p��#��խGKG�u՜uh��x�z��x���GGQ\q�-u�8�eDz�-V�8��B�uj�㥺�:�:㎭�[��u�:���-n�뎺�n)��]8�ձ:���<GQ��"��ӈ�����C��q�qV��ǎ8���Ǆ<[�*��t�֫-q�#�륭�:��[���:��Ÿ����z���>Dt��E��ޣ\W^<q��e�����Ћ[Ÿ�~qӥ��G�8��b޼u�[�-kE��8��-Ǭu�ţ�z���:q�:�!�h���θ�zx��u��=,�Ǯ#�q�ޢ��=z=x�Q�q�#��ޭ��ǋqg]|�GO��u�>x�-�8�GQN�!�Ƹ�Z�[�0F�1B�S�u�&��VӢBT�&��)U!L��u�"�<tZY�]@TD�~�<|�HYi���yB*�)��d6�d�a��!�Ϗ�M�!�h78��A�T������8�S%2Z$#模HBH�U�&8��	>�Z5�(�@�*�I>>�$N�vJQ�I&�Ag	hB��TL:�bG��e���Щf�&��`*ID��&|�D8n�06�.���HD�͟!Q)��T �����=3/�2��>�	O���ZIC0c2�*�횐�L�"`H�Q�92R���R�a���#fZ�o~q�p��
���}X�� �G|��y��|v)����;��T����ǿ>����O�k�����*�3�q���f*|��Y��M�/�Zl�90����+%U��7#k�q�Md`��2�q@��Ò޵���)�4�*�ű�yYvI:C(�yuy$,0�ʺ�C���XEwM�c ̂S��.�2&�;�yD��An^t�8���.vu�_J���.�STa�;V���;�]�=��.6a�p�wwm���E	ֺV�\:`��'Y!�R�V����e����8!F�=LgZ��=4R��Y����D�O+U��Vl�A�S���UNݎ���~��*�	�n�,q+��}t����<�\0RǂU��S�);:��r�0U�i�r��`ڎ�|[��{ZE��oma�v{U=�%y�88j!�i�����T]-g5�̭׋�{�n]�G���m��}�9G9�PR��������+���K�d �-�ћ�M�K�/Uf�{F$I��㍳D�^�feǗ-N�DΰE�B����f�U�U̝�-����m�3(��ܸ����C�u�6�=ՊN�����ͷv�0�e1Nf�qg��HѴ:�5chH,u�o�Z���BK�ō�(�v��=�*�1<�n�e�Yjd��ۋŒ�x&·qP�c��t�A�ѵ�"q�k�R��sID�`X���4�M4��M,�M4�M4�!��CM4�M4��M,�M4�O4�N�i��4�M4��F�i��i��h�M��9�;��ƶ�q��Z#Y7���7��"ud�\�ݫ�ͩ32��0�}��ur2�;*5ݕ����TС�]Cf���'��M=8���OƎ[&��7�f/v�E�mD��K��m�8��H{Y5������c�xRm*{1A����VV�=R�*Bvvu���={	�OWs�D�#Z�u�Σݏ�<��Jի*֧R�㩡0)@ǻ�M��zM�n�)p�*0��X;��Vk�f�z�5��v��x۷��*��̓��e�`YgS�@�W�C"�;f&�{)Qpg^�2���
n��#n�["��ÌR$��23,��Z��إَ�m�[M���v�)���zj��Rrx��ܰ���fނ�p�7a��׫N�xtљL�ʃ]��ayS��sʞ/1W`809$圉�1�^�6R�u�7s�,c����D��K�pfm^2��̷r��g�s��nu�2��犹g��i6g]@+!`P�ZKinc	<3�3fJ�T$��v�u��ܛIw	b�rŋH.Ѽ6V��I:�okc+6�pW�����aJ��m��o��o�r���ԥAH��n_Z�����kՉDEl�ʍ���ZnXlU�!/�8z|z0��M4�M4Ѧ�i��i��4�i��i��i���M4�M=4�Ni��t�M4��M4�M4�M4��Hi��k�|��9����[<ZD�Hb��=�Ól2�n/9L�Q��7}��\{kG�����V&<sƖ뇺`;Um��P��o��T�����6�.��mI=��ں�9�K�Z�a.Y��k2R_b���/��ʠ�����㨥�y���A����pU�����5��L��a���J!�Y�C��-ff��	�{�N�tt�t��t�`Sb~�{S��Vj�Z�47M�^�v⇏�[�m'u-��U��L����E�-"�:��{*�9SPm�H"9k[��
Y�py���A6u)|�&rʭ�ee`��T[�DV�GcB���JX����!�|ީ&o;L����龂��ث�m�6��&���*W��g~�Lmu�S�̷�����Q���`D�j����3D��L�Lٙہ����{.M���U⇢��t�`����l�HB�L�������f���wu�hgG�hV6�JZJ`b/2�]��VT�g[R�Z��MCjU+
v!��U4��m�=�����-�TՒ�]�d���q�6t9���{W�,�L�b5��ɐB��em�NZ���&biF⽡��x -1�1�tة��zݒn��F�Jee%v˘./\�U��C���Y���(\9���ņm�{F��h¶����Ϫ�bq���K:z|=0�M4�M4�Hi��i��a����i4�M4�L4i��i��|i��i��t�M4��M4ӆ�i��zi�h��h����z�d�b`ҍ�z�,@[g66�����1 a�铭�Z�CMq,���%��DJ�㊩�g�!�Z�2�hݱ��V6�H����4�d&���5G�j�]i�Y�[Ӂ���
��+K!wXUs�0AxR��o����^e�0��0!9�Y��>���J����zWo�<xH��nc��h.�qgsa	[*�{C��^V�>г灞��3������!�O�z�r!�۲iJ_ ]3C��Q���❀'ԽxA�/��f�3�i�1fRPNr��3��R���!����E���:�@G�j��S*�Y�����n� DG�obu�=}��`�~�eM���W@�&�u�r�)��7�o`�QnҀwx�N�ǀ
Y���
���q�,QǸ#=�&���8��ܕcޏ����Y�{�&A�>�֍9��� 5�L�yK����9��ܐ��ʎ����t�"E���\���AN�'lYZ�0��mR&u�	v���p�Pc��Y *�,����T/U���{R��� g7d.LT�K�橉���L�"��R5Uf�TO�����{j�:�Ә8�����
�0i ��+^�%�]�r�#��r��#j��Abm���J�]3j�fu���ݲ���ِ{�5*��R܃�꩔+�Z�k���VJ�󧛕-��[ �����C�K�.�l w^�����F���=Ӯ��*��`XzzC4�M4�4��i��i�i��Y��i��i��4�M4�M4�Hi��i���i�M4�Ni��i馚0("ݱ�1[�C&QT��8nt�{���g<�S/uە�^P`mr�Vxod������u9m�5H���=�T��;e�i�.�Ѻ��0�����ӎ��"�f�[9~���Q�EK�"�u֩u��V�d�"������z85_�Cގ����
�����'ec�bs[v�Eҹ.�N�5�;F�n}��	��Ս�tpuX2�}%{�b�u !��m ���mˮ#�H��� U�{��ݨi
�i�I7�h��2su�����AA�<VcQg>��v!���B,�=������Wy���R�{@�!�M��x�lP��ꀢK�O��|�G9u��%�Y��X��^R��W���@ �����΍�ISD�R�$<U[n�͝�
�N8.����
���x���,f��ہ>�5J�
Z�a����t!�
�V�sDI�70�;��;Ptf&��P7'3��6t>]���1��uw���IՕ�M�W��8����ï�����;�.�RY� Tc=l��J��LR�#rȈ�.�D�Z����g��:�S���_Iz1 �tj�-�܂u�x���Jhz8,��������ָnY��Ǜ�V.\��ɷ�(�)�c��,�cH�)�����d�Xh����sr�Jf��!�mjma�=��6[���S�n��)�:���uTf�aY;��{��l�g=��0�����M4�M4��M4ᦚi���i��Y��i��i��i4�M4�L4i��i���i�4�M:i��iᦚi�M
�H�F�aeTB���m"�Mf�ž������{&��A_�����u� ��v@� l�v0��5Ҏ8�K��p��s6����
�%jGN%��%�a��bd������	·Km��uT���孶�P��7-�=YF�å�>Z��f�p�S������s��.��]r	���:�Q��&��Lh'U��[�o]�c=��Ws����@
ӌ� ��=�#��p�y�y�&�^������;��/%�nP]tP��3hCٖ��)��wR;���a_N��O &;����'-��K+%��.��b+beL8S��;�f���G�<e�������6�ל����q('�D��u��y�X�c��)\ ���ۙ��F�joK�²��ewm�Ld�wo%�Xp���4�k��)M�WS�����g:��L��V��K���MU\ ��s9����Rƣ0T1vOդ7��!Ico6��+w�9��R�xA���k^�/��ɽP�lr��`s��[^�U��J��ݹ�ݶ�a0���Ջ��r<`Btxn�L[+��0{8k*0�A����E>X��a9T]>�n�j�^e=��Tۮe֎X��*���uy�,�$�ˋ�� �Kuk�5Nvӻ+�$�T�,&$-b��BS�ޚY񦞟p�M4�OM4�Ni��i馚Ye�i�4�M4��M,�M4�M>4i��i��|i��i��i���i�M4�N�n���������rI�P�)�]��9�n�h�}K�����"�U�Թ\�̛`�V]���O,�㚽�r����w+��Hp�ެ�&Uie"�6�lm,(R�6��	��-�f��od5���MHl�e�[Ǔ�}���қ+P��껨�r؃i�D�*�57��ܴ#a	t�r�b���w�k*�s"ɴi� X/n��8�Q�ȧ�J�EI�_==ו�m%.�R�Jz1��B!�dLD���D�Iy�97d��Uy��n��Ƀv��wz��[9�;.c��'��x��e���1�87J{W#l3RjA@��b@�m��	�U�g_:��4%l��9E�3a=qnwK���Ƴ(aP���T	z�&:�dWO+�x8��W˱���ۆN��}���r8.��Z�B��)íܔ8�*��"�pJ��:&�}��f���}]r;3��V+e�S)j}}^S�k@�v$�U��v;�@d�D�Ơ��u�e>�ފ�9�Xkv�l�F�K�D*�(>PCN:Z��y�*�h{S'�z���x	��B�r��L�yz^�*h>:b�%Or̭��z]DX�u�vqy*==hfet�&�p����ԍ,9ˊo��7y�����k���O�R�D�#/-6�.�wOQ��"�������4Ӧ�i��i��t�M4��M4��4�M:i��iᦚY��i��|h�M4�M4�!��i��i�i��i���gfZ_�Ͻ�Y{�1�{h;�	�tV]j�M��7!�;�BdT����nѧV��*�U'Ox�{��ks��M�uu!;a����.�9����a���b���g۸�X��^��ah�В�&Ъ�e1Ah�Ķ�!�#NZ��rm0k&�Ġ�L0d�G,��� �$U��8N1�n�������S�q�*Q�ܢ���[�j�I��`��DaF$�6�-�Or���*Q���:L�z1ef��XlW�U��
:���r�m�6���ָ�:�f�����	S���"��P]��>Vk2m�}�IV�fʹ�EU���M�Ѕ'K��M�g��G��\J��n�L�Z�`]bT�U�6)����v��:a)������*��pe�f)�[���Ow]�3����m��cB�z34k�pqüx��osNbr.����J����B۱davm7ˬy�V3��f�.��xo"��{�맃,1}R�7SWK5l��X�jSq榽ȃV��'aBL�d:B�mEK�n�x5Լ=������Y�Wi�N���V�̜gDi���FN����4+h�f�EdG�
��D��u=+F���}��y�:i��4�M=4�Ni��i���i�M!4�M4��M4馚i�M4�M<4�i��i��h�M4�M4�!��i���o8��gg�rwk�h/T=hn �na��ؤ�+����h��u(�Э+�j�p^�!/on�钕�ҲO+��ۍqA�e3�=N�]�;������Ǟ�Z�X�n�������+��uZ�>�	#���>]"�n�u�1����UPmUn��e�)��ۭ���40��QN3D���:�Hs�w�K��BIt����2��*i 1b��vގն��������W���R���Nc�����l�̂�%�7
LT�j��I��Y@̠f��Yv\`f��v��{�Ue�PP��%n��;�������p�nc��s�Wkwj�`��[��;ՠ4.��AR�$�5&��s0�"D3W9Ys'2l�GZ�Cd��B����|���sk{=~�z�GA�M+VA�`r��v:'n
[pJ��D^���Q]d:�Ln���=W�}��X��O2���2�P���n�4��Z���;�v[�I�ud2��s0��}�1�/f���5	�t.]i��V:�'<�����U&��n�L��ג��R���Z+/)����̜��5�@�mL���e���t���s]��ՅՔ��X�)��yF9�U6'wB����bJ�j�ɪ��gJ��_f�h�q�Q�-��\��A� TfM��Bi�RXm���a�]�om���dV�����n�q�4-��51(8�ŋ���\�+fƹ�rB�"۽uB��7%������m&�d����C�Vf���T]���{*s�dV��Ύu��E;{�iH��utVاa�M_�@80�U3�Y;�ֆ��]H�mc@���@𷲣�z�Uʎ�q�+wm)���,���+���=@�gr��AfY���.�5%
���:�A'V9H�κ���k��.���AGor\����O5�X,D�Z�|&pf���ѓc�WB�X�XM]k׵)i)i��˫�e�����4�m�U
A
v>�A�Еܥm�Jr:�+^:�h���*݊XeJ3:+7&��R�4�u�ѭ��m�NȅZ�:-A�UW�p��#:�pK[�j��˘���9����6��!�ؾ�Kv�X}e���29Z�X��6�J��w+:�ĥY��J7Te�\�}e\�j�y�U�Q�����k�Q�d�d[U�5Va�P�/�@v
�5T�<�*�ë4�XUyj�XC�W�4��*��=�rۗקnS#wfG��yp֐�<v�]���qŧ��ߟ@�+�����~-��!�O��"7���0�.1սV[�q��oy�q�l7�1���&PF��	�!�Q�����)��e��$�G ���~*�W΅����OE�d���W�϶}�9��}z�Yژ�! �U�[nv[���ff1z��FV�e�T��˵U=ȷ/+mnƏ:Se��ґ�lV{r�c\��XƏ؉�͜�bd�Cia�B��:�1)Z2D:�ȨR��VZ�Zj�,�AQ�O�۶��D�tsT	˘D�8����g%�f��G�8�����%nܔ�Ү�]Y@�0�̒�[�ͪu7�,V�{x�˪�ܬ�dCrR�A�E���Ǯ1��o�_*m���tv]f���%�\;�{��S��(Uh[�b�E	�^�3����3,*��V�:��D��g
�h�&�A	�ܝe#����eS�&71ի�N��Q�Tm-�KVf�[8���,���&��5}x�͎��v8��#iu�ʹ\�d1G��9�t.YwT�g�u�!m��v��:��2I�`;�.Ϩ�֐�;ݹ2����&�PH�Ƣ���j,n3424+wLY��z�%~�w���,֪vmYd���omBʹ��ֱ����2�Ԯa��L�$f���"��K�t ��Ղu<oO)Ə�'�f�fru���u3y&�1���"Y�T�����E�J�lEٻL<�n��-,ς����g�q�-�Å�G��N���E��[Ŭ���8Bգ�t�^u�]-[�GqY�Qn��q�\u�]Zp�N:���8�V㧋!kG�-��qku]Bȷ8��-���QX� "	�)�F�17��l.'B��u�aF�H	�%����?X��~`�Q6��ઘa�
ȑ��EO�A�U���*�o5�5���|��QAEA99QA@TUIE�U��p�IRD����xxxt���jݩ�&Jc�L��F�lDz12����2!֌�v�Ext�OOO�4�Ȼ��`�Ŗ4aC�DYa��2�	vJ��%�\E�DK��QCAa�Cc�8aaƜ�$"$%ŉ.�Z�Z���M4����*ȴ��jB#��\]���BR.�rȞ՜�b�ʴ+�U��DHQ��Z�� Z2��r�� a2�(J((V��(B.����rޟ�ǧ���~9��B��"�QR�R(����`��50�FN
o5�������s�,�̃�9�P��Z (��h�6Xd.y�j����~:i���?vFG8�")�S��y8�B��9�rлX6``Pb�փ ��z���V�E�84&E9���d��h�哒���Zľ��H�_�����?�Z�xX��a�p����b`�0�7��h�r�"��-�G.J�����K���,��Z]�H��Vyg8�c�M4���ƚ���"1�0�i�b0�*�p��2��0(#F�a�4��q9%I"o�M4����N�<A�aXFAT�6Z(��%��cTZ,�ʩ(���M�C���`z֍dᘵ]�փ�\O��TH�C%�r��?X��&�q'��` �cm�ա�^b7���/
_���lne_
����U�;�d��
��eG���s�gK����dx��z���뮬�� D0 ��~A�H�f4��"$E%� �RAp+G*z�� ��?ۦ��٢vDwa�f�'oŧ.\�(��W݉|�._�����En�`�?:k2(����3(�ZH�]V���"j�t1O�5V£���ɧ��z�i�	Ü������1T|$�0AW��z�ʯ�[���O]>�y��6ҹg�&�Z@Ávɐ3c�l���.{k�kk��������򆹛UV�.����Wa��e���Blg^Q�R�2���y}��˕��v����lwv���5i�&t\��e
���k�|ή��͌�.���������}�\��=��\�Q-���#N��t�N�"qG�vL��ʼs_*��]ϱq�#��z#3�������>��G 3�5'����[)G�0#��Z�vy��!�z,�Fc�ԯ/<��Ay8���OR���!94��O��p�o�F���W��gik-�j�:�G�>��"-��7B���t����\�����v�4���y�F�gV7YkP.�nF`�`a�	�8�/C�;.�d���a��7ү�oT�:�o��K�o��'�����gLI�6S���O8�r�l|�ܡL/�|C��?P�{��n5͜��F����;��럳/�l���4~���HA�z+����ɊT]ӳ�ݔ��	Ĺ��:]�P�x2N��6���t4��N�}Y�JL	�|"^j�,Ps�ژ�9�w\�/'�r*�F��\�^sI��&������k[_u�@[�Gq�k���[k�9y��	��Y�vw�X����'p��#�9^y��/��Sy�����mr��h��+��V��[Y�"|��i��)p"RΘ���Cڥ��Olnv��jվ��Ho6��Oe|ok�@F�M�X��O�%������s���{���t9���fŖ���}{U�n����S���v_f嬔�qb�n�^,�M�s��V[CFOF�]c:�Y2]G, 	� A MX'5X��jn�m�B���5���Q��N5t�8�n�%�/_+g/��bGz�^	-f�y���/�N�vZ%�"�z��&�!�t��s|J�;��� �ةP�U���==F�t�s����V	`�s�iF.�<U�������n�P�<��k��S�{TL�D�~�5�Z�p5 3e%�ܘ�sy%���<�:��韫�b��[;���S�KFb$���n{雌�.�Zs�,`�UP���ⳍ����r��  Pc��c*�ɑ�K�*_]�_O�7ۈ�}�s�ST�-�� �zW�k��;q��
U/����rw�C*���Ƅ����:tؒƻD�W(�#
8n���<߰g;��a4�S��UvhҎَG'Zr����dX/T��~N��`��8p��`\m<3f�,P�a+��i�5�=����ձ\|�yP5S�w
�H��OlT�t]M�G���U2�ᘶt�,]����9�͎����e4���?|���6(͹�We�U]�5������Zy�T�9$K���EE�MRa����2ݝ6і?f�ğ�ϐ�=$'qY�m��e��LPZ�A��s;QP��TW����E?���M�=�% *� n��B���\oZk��щ�6_�.�� �4��
;��2h��0&�h�㹟���뱍��m�b=��A��	̾�φ�[rOUڽWj�t��ѿ[�eN�lE,�3i3�]ؖ�oZ�\�V��b�\���m�pn.�7���1	��3f�Zw�7Ǥ���V_r�M�Pg�k���n>��W&2E=�$3���	/��d����9�{٥�צ]�����3�\�3P
��+q�'��3-���v�]=}+o�fV���)��I�fى�c}�pP�,ښ�J(�^�Et��=2�Ꮠ��X���ܤ@V��C{돍��x%�e�{x`���r厢:,��ޙQ�9�p�^�T�@j���:�����
�]�D@Ǚ(-��1ͨ�.˲F-����6��T'xm���n��!�Y����V2Y��u��AK�.��ƗN��5��zy�&Ž�WS�g(�.�;yp�Gi��*!e3j�53�
�G��]8�e��>_@��Z���ź���w��˗-�	�������4P�6�� @��a&�a{�����4O��0�`9�}o����c:��כ���rux��l�	}�g�h�z�s��+�U��Ww�/�D�|x�J�뺷Ù��Yʙw��SB������/L��(4pA����S�l��H[�\���G�܃`� �;���kXX�OM��G1FX	�R6�]�E���/���zNv��K�[}O��X����7����]��X�M�X]֯i[��uJ]F���ư�<�.� ���ȟ��8� ��x�W)��;[��;s�p��l�ݪ���d�SW,�V8@(G_�U+��w����n�ހf�u;��*r�Y{�W_v'�JX	�����Q����@O!	x�wuV�{���v���{��.W��0��3�4!ڹ%���2h��.�:v�g	��S龕�`���-����,�'�~�hN��O��ksrӪR���fЅ����83�@A�1��WT]"ݷ�q�� ����F҃q��d��wO���k��L���a,f͹��I:�r[�w�45����j��WOPplʪ�.T���{7���燇X��X�M�N#��sJ�w�{����}�~�+��x˒nK��\��V�_V@�k@���vμ�p�@�ri�˨������ �.;=-\H���nS}Ϯ�a���G�S���L�{/yR��uj6m��(��[�����A�t�3�$]�s�z�[��Χ[x~��w
S�So�����bT����#�u���ixXʒ�̜�� @����J�w�y:}_N^�����]8֘����}}�]_IPI�bׄ������4��K����m<�.Mj�4��Z���y5EP��x6���Ă���LL��=P��w�Wg>�Os�D��g����"��Lc�W���a��꧱�adun]喴��;�Sռk)]:�j�@��`���4V��>׶S' ��-6�mgi��;�7��K4K�ǣ�O���_S�E�Ώ��[���3n=���Q�-;;������)�х����ơbYq{�����%�Xo�Y4�LҸΰ'&]��ˢ�>🻯N��y%|]�{��,fl'����G��`L`��R��C^$a�4�I���<;q��|�9��k�y���4��q)��7��yz��>���;=ܔ��t����
��P� h ǵob|��n��Nj~]�3I=Y=��L�z؇��5J ��>cp_"��W4��w��`_��IG��э<y+��CΚ��J�g
F�Ǖ�2 O�'O�	k20@��cc��e���4����bz�� � s�� ��6�Nu�EKz�E�_VAE�MGiW��5�f�NXHD�d��lT��O(�f;���]�� _b �U����妤������������ǅ���^r�[]�U���� ��XyvxX}���:�LZ$��쾎խyK~�C{E�x8wJ�F�ɓ��n�vvJw2��5:0"�,�Z"�hs��܃O�ԧ��8�5	7���#�=}B��T����4����;D7Ms}�Q��6��dL��S�XF׿I	�Sז��\�A#���c�>Q4ډI�r��.�nu�s�dH�@E�] Y����sb\��qc;+t�;�tu�:r(��1_JΑ������m�N�aκ�l��B�/�V'�	
/w��=���,sz��`��?�Fi7���܏�-�7�Tj��G��P%N�~���Y|���r�����ǔ_Sb�V�H��L�}�&�`k�7btHwF_ۙ��7R�@��q��f�Du�l��c�Al��6l��#����F���29^�)񎜮����  f}K���k4��O�����.`�NFͰ���1{�$�`��������ke��Ϟq�L=ˉ��E,<��6@�;�y�u#Wm�,�hH�f�.xep���GݯkM�W9��	�fk�k�τ��	�:�������w5;ic?�[ox&�f�7k�-�wN0Q��2��%:�A��wb��*J�Ry���cD ��@A��
Dહ�׶$ĳz��\Aخ�k��w�z���AŎ��˼2n�\��˳HJ��o�NtU��׎-Ëqp�\w�;|w��a�!yT�������<3����yb���c���]:?d	�v@vnf<��4�y _�C5�\Jiwo�U �=���$F,�3
:��uԵ�Í^W}2��@v������G���퀴]@�h(Ǯo4�]�o���Өt!31��ʦ�{'M}��q����7B:���M��=�w��r/���� ⼷@�}���`^K-;ɭ�G'��=lu'β2_'C��@F���=�%b�(wl=��:[�����in��q�.��o����������+܍d��
��v+_��yb;)�ڛ,�}7�ؔ�����C���LP�M n�Gdf5�/�|�[���O���r��^��+h��:�X�{��c6�J4��4 ��e+}{�B��2�� I�Z�HE�'��^�8zvafYwd�*��e�:�;$��ǱUv��ɹ�U���w�"l�js6E$#~Bh�M��z%l�n�7I����� ��F�a[4�.L�7oH�Phk��p�M̨ZK�f��U+3Md�:��ٝ[�ZN���CIn�ۂe��>�c��Kvr�K�_�S�×5t9ub���l#��ol��]q�O
o/nzܮm�����F%C��H�1D�$
�����C�8��Ԗ���h�i�5���>ͭ�gY �˞�#:w���Ek����~)��91�u�����gY?>ݛr�g.>|�����_��ݚ��N�XL#����|�`�>���\���Y�<	��]s�@� v�F�>��'��>�B��K�Ɯ���K�g]��LV�96>Dgwfv}Ý! BD�-B�)mt��*qS��2ʩ;�W y�>'VS�ȁ�nT�8�k;�-'U˅����GB�f��':��|�A��p�&�׸�.涮�1\�.��vਨ}�V׀�+ښk�$��㚹��8�sC���VY�u�#���5�`�xH������Xh�![@�+6����vE�=j�^�v���VsRv�sWZ�O��ܟi��/;h����JS{[��t��9GA���ݎ����9���$�ܸ'J�vsU��LN�E�X+95�fV�X��+*V؜�]���{]�j���
�.[ʝ�VN+�.��k�3��	�tm�B�ޡ�V�Q�i�Z�7��,��Pq�z�9�W|d�2\��֖�=B�BP6��qx��q�;��L��jme+��_�S���X���3]��%���hx%J��mzh�M�;E%ƴ�}���lK�ղGLGS�J�=��A�uwOL�q]�1l�����<�Z�R4r�^�-za��iwr�f+�2o"�m�����c6�9���}��}�.��K�8T��b̶;�x�Kǡ=/
�0Q�O�J����n�+��X�Y	nfc�2�,��2gu�^���\euV���-n;���K�˕��A�9���b��f�KI�u��ɵf("�^��s��\
����t��Кv���[q<ie����\�� f����W�n]6���o31�v2�u�N�
P�Ru��v����l�X���}��#�mm�VmQ��d_I���q� ��L�eQ)�h��m���:�c{SЪ,�Y�v��Ez�Ww�W`�}�k;�&�$m��¡`X#41a�(0b@�s�`u� c� #�	�`������RLGo	���(�����Rn�b�$]�.���T��o�E���`�Bڬ-�K=�9gs��L��+��9����Xfm���;]H�ҵ�Z[����U�9�y���mY]����q�W ��Ռ^C6�E#
��9a�c�����������f�!�T�j45��s2�S�.�q�^�%�z�(o�uE���UgR�Ղ�լLֶb�*Mhiۥ�m!k %S�Ky�ei)��!�ݳxXfJ�kE��nD���5�aUN��U
�: �����A�j1G+rm�29�5����|6J�m3�Ð-@�sD���Ε�";�}�4��	#�)��jͳ���Ȃ��g,�B$�O���,�ӛ�|�y�4������=�)F�ż�a�Z�U��2�
��!J��ז�IŒ�����lS�xF-<��*�N�Kv�]ݣ��8��{�A�n�Ix��B�ã�R����<U�m֋��W�����֍�ۡNʪ���Ƕ�=����N*l];�&V0tI;���L���Z�E�;�.톍7�]$�S�*�iE��.X�uZ�m���)�!�-Z4������.>�x�7�Ȳ�b�Mzy;�z�r���	 F��A�&E*�_���a�;�A���������a�TYTqQF��>>><0������;˸�#�ڨ�	�����)������:]Z%D�[V�f�zi�r��ow$�QUa9RYDfMHQ^A�%"U}*C��t�����N�7P30rF�)��ʈii��rB���:���<���g��PR�������,�h�#"��Ȣ*I!"�S�r��0��x|~��������J�B$�� �9*�����������lu���1�ơ&
Z �-Z�,���^��8���qUȩ)r�&Yq<.�DII)"@��݊V�i�Ǉ��u]@�J�D�DT�(
(h
VAQn2MA�B� �!��Uz,�	'�I I Q�}��5=���.�O��-X�͝��,(!��܉p�M�S��a��4v>�/E�����M�Q7+ygw�����  D�`�o5�k��{��9:ف������9<���}C�>3��@�%h�O_ԟ�9�e�#�#�S��,��,ex~z6�΁����'����o;+��o�̏e3�٬���=��UA�C���|����[�/w~��!Ia���q�^�_��}��-�P�{2���тw��Sx�X:%���O[�X��x�H�_½����Q�!�;~�)��`U�#d#>�{v��+e�eŸ��W��	�~7���p$7�����t&z���0�X;��n�ʒϕ5d����Q�o�Z �N)
m.�[��m?�d��x ��6�D��e�f[
�Y"�b����Lt3xSV1��~����g�%e�l�J�l��`[���g�{��2�{�_�Z��\����[9-��v\ޕ�;�W�%�͡�xӦ���XH������1�|���m_K �1:c�m0�y^YV�Y��PAPA���n�C [ŀN���ǽna�$Txk4z�C2N��G8�c´Q��6 �#�WP��p��.�%>��l̽Iz,�ٹ�?�`a�Nޟa4�Ù�����C&�Q1��Y��Op����`�U��������\nw�6�*�Q���{�J�=Ni�Jnq:C0��<ӑs���N����MDM����^3������{L4�Ő�+gky�/
�Z��K�����"0`��ӽ��'n�bu�:]b�>fQ�o[��8p0��[ݧ�=-��*>_T�&����KCxc��y�4cf������~n���\����x��u��uf-�gH���{�[[��'�*�8oW�!~6@$�C�皼*<��aב��p\�iM���|��-��D���&`O�d��|�� G�!��Ϗ���R�м	�ׯ	gX��{���2U�K��m���ù�����5@#�#����"� ��Xc�`�6��b���mg:�u��
Z��_i�t�J�^s����^�����K��x�|#����Ύ��7.5w�����Ǘ���#���`���< �;.�ǎ��E��q��M	����ٮ������4���~���U���\z�/fǂo	s�^��%�>���/�g@����-��g��*p}-xS\[-m���uQ����x��3x}�H���3�Z�����;�MQ_�y��ϔ*���ٹ �r�y����3ns� � 1F<5�fǂhi�����P)��NC�91N�� T�F��W3�l1���o��NN������>x�	������_�za�/�-��0�n[�������0���������9Ur������񟺩'1w'��V��f*�k&j�d��늣�JDk���2�mƛ�SrlLo0�
�!)�n�!���PC�oMf#J��q��m��C�7�ѕ].W$��t��{ÕFr���γFI��c��Ёk XbD �� @��nFTf	I������V��j��|z���]w��~��q�E��r�*�{q��xA��_�V�C���J��?p��zvh"���q�����1�1w���镤l�ǌ9�9� ��[CLx;a��m���x[H�%Ǥ'�,�(	��-Crz��;�6�K�n,�wɭ ������|+dd a,�`G�w�R��̣#�@-�>�`�����No�����t�5��PYl�=����o\kR�m/��G���T6������s�]<����Y6�d�@�����_U�K�ؐ���$D@�����`2����2e{�q߿?ֆ���3�&mcV:1��Cw|�7�?|8O�s̾�)F�]�hO�����R�a����Vx��sF)��֠_]�{��a��=�T����s�|(����BK�>]�����ƅ7���y?��#��2��%�����wDv��9@s�|��u�!�������C�y�� Ĉyd�@?�x�C|'u��
Y��{zDL���y��l0�і�.��C���޹��}d���N���(H�/\��q��za�$���C�R�+eÏ;�#z�f� ��c����`{ ��M
����
`�0��Q�8�vs�T��_1�f�%���R\��>2t,�4����\3�X�;�Cz����[qxM�kd��{y2r���˦�mҩ�5�u���`��X{��[Ŗ�dJ�}�.�sf:Z��C�u�'U]^Xʾଓ�^#{&�&����M��u�F��֤Ȼ�$D��P���'�)~��o�px��y�+�c4w�������)��7�g�B�����K95�5+��k}O����m]�A��?4Xq�G�J�Ӹ`p{���5�K��$� ;�ʾ�Lp��|;\� �+��Zׄ0��~9xD��Fc���=��ge�����.OM���UG�,�<�%��ݞ�A��"d
�O��K�&G�ΧGÿ~~��0	 ��M��<
���-��n��6s��Ƕ鶿b��,Ĭك�>�Ն�Cк�� ԀG�lt�4���K�|"�%c�M�:3;1u/xG>��Zk���u#�a���Pq�'=0���/���?@���pJ(��2}bok4ϼ��(@���~`$p�W���/�;�������5d!ޖ@��� ���xH���M�kٮ�s*�#uQ [S ́��>��C�K�*a7o��X�G���ܪ�,���5F�ts�����Z%�o�����Zɯ���k�/��I��%�6���ksZT?���US�js��o+}�@��/���Ax�Y��8��x3��N>���z7��_F�N����y*ZT��{0^*��JJ��a��.�l��-<�S9޺�g3gN�����2����q�@�P#����
Y|��
R����IZ�*�n6����'s`tS2��Ъ��Tz��R�A`/�uMg3��<���?���J�dT � Y&�0���ݞ,� &�p��(?��@�g�
Bx�i���Tp��O�ȏ�����
w�X��:ѳ\�J�|l��`Y ��	��A��?�TP����K�kLgO�3Ɨg'jnbh�-=���{m{<=_��f�X� !�H��"�͑�#��  *t�G��� ��V��f��O�p�@k0�z64�Q���_����=�'W����q��N�4��g�3�ݟbyr`�$@�(��<��@^>DK��1�ߗ�1��}B'$�Qd��c;(v�T��� K	��v�C�<���q��`5����A��g��Ү>����(��1��̍�p#�A�;
��=�~'pӠ(�I��4�Cl��xi����;=����Ļ��;�4�;�3�Ϯ����������^���0�ͤ������֊����S�h&NG'�M
�aҔ�'�vb�YS���jU�����
3l��%M6Y���.���4pS>���l>�iv��oii]x�����@D�C�SH�4h���-�����
~�10n�2Dze�f�(7�*=+��/!VH��Q�TD�4tn\��LΗ\Κ4*娮f=�F;u�%�FA�bom�� ��Pה��1i�͝��z >���'n���x8K�GLL7��`�p×�N��Q����L�+ʼ7���J�����\�e¶�\���}�s��|��UO�P��]Ҭ@� A"A8�\�=p�-�z<.����?��7J�Dx}?�ڭlQ�	D	kҦ��ʜhi���]l�x�fw�vs�P^��ݍkg���@3�Hl$B��>��16���h������(���N�6utu?@p��}Y/똘�sdo� �A8���Ͻ�P�?u0:�=)p�lɤ�䁁/a??�"Rݗ~��YH��+��'�z$����G/�!/��S���N�mE�3��b�AT�Mx��+������,���z����R'a���8�ҏ�&�.pN <2[#삞��&-C� �hXO�Љl���w�]�O�������T�MVz�@~q�(�eH��$�ldk��cՠ��9��=��o`�A�f�Xmw�:�76���E��P��i.�`f9N/r2;dy�	5� ذLcc96u<�MA̳��g5n �|���4��ǀ��3���Eq��_{�^�������ɹ����aO�U�&���S�)�yxy��b�Ƽ�8�͊^[Ø~�ܽ���9%����E��qgtx���*���
�N���t�,f�YW�ҭ���0�]����)��ms�s5mn�*���w�|�.�Q�0���I�t�K�R���]�ln^3��4�II��f��:��ں���XU3N�#2Z�����cV���*���ѣ����ke���S�@�p $�0 %X!2SU2B �8�8���{��~�Ó��!m�p>� ���9�gO] AK>(i���o��T{���X��R(������4�5�W����c�!-$����;��3�����?�����{2�)ڍ��vk3oJ�@g��:�����gh���F�K,}R�_|�!`tk�{���J.���;̟,�|e΀W�O'!}Q�)B"wҍ8�zb���t)��Մ"���C����1��;=�:v��� ����5���薩0S �
���4�,5Ȥ���� iyN�_{,�o�R�PG�ͺ��=���b�|&;�(񊜇V�toƓ���^�c���⵾^��� ]�8�6s׭fP�	��w��6��E�H��U�x	�����N�oaٜA�a=ڷ���_��;���zJ)�?`*}�j��59���.2�FA�I�:���0{a��x��><h޼�-�+�k���� G��%2��]	�l�6���)�Qʹ
��;s��X��7��D�U�OP�mőrz��I���=Jq�{h�s��/ҍ�;�
���a~ZT
��c�VR�c#\Ǳ�Vn�+�c��,��؞&q�36TYDf�_,�׽Hwj��*`@% p���Y��m�Hs��YY�iȦ�Y3'*vΧ��T�:ru�Q�)�L�zmY��4�`X�on��0VX�f����`�`�N�P ��
P��$F	�F�2Uou,��9��HC��e��#�LD$�`T�E�6-9�^AOe��_���5���4<5Mڈ�Pض@'f���|����Ɨ�}O�^YMNW`�EH�,#w"F�tq��\u�@�od[.1L�A�p�۲��@qΘTƾ�?&|T�l�O<rv�A?D�v��^ [����a���4�>h	��u���?q0�~��92P���W���vE�w��e��$�+���B��������Q�  ��tZ�L���~+��"�i���	0"j�	���YnC%�J" ����x`m X�+ ��#���:�5�K��5�vO�
��z�y� I��x�����1BW��[���d�q�#�: 3�0���jS=�m�:Tq��(�v	L;j��4�;��-�xa�i�&����%!�h��Ɂ�GCwmy����F�I�o}���m����jT��lٵ�K(�e1�@.{�DK?^�aNXl�Ɍ�ե��n�%�$�O�Y���u�j�f<���S��
If�·^��~^Z��s��q1.	[�dQ_(�K�Ē��u�.
��gYO}�`붾W㶐dN��T����(�Ř&�p�k�
\P�Uk�|A���	*S�O��uYo2p̙܋Kh����%&+6��Ҟ`V�.���k��<��]yƵ�0~H�Jv	��H�`B�� (�@�dCM@	B4o߾����v�[�º ��'��B�M�h�1Oa�8ǕY�z_��A�Ɇ�����:c�g���C��[��t^D�����z�%й�s�t±+���m�Sm�7�!�o{�~�2_�o]���Y��hx��s`V���J��8���L��~l���}A�'��_�T�u,�hU�f@����vƨ�lyO��� ��=�)X�9=�F#Y(�|�#K��8q�7�~���A�	�ڹ�(��1z���yB��t'�F��u!���7K���v��ՓkH|��ݼ�U0�0����F!s�3�o��n�xB�/B^y�!>ynlAl��1~ݶGcjW�-��o�M�4��u�`�`ùƵ?d��{06�BN�F鬸�s�,��Y�~�~�C#"7�xr�9����W���!<xx�D�k��!��*"�-�zP~r�z��B��O~����`h~���S�w>O_ۡ���B�1`_'���9X[�w
�It�n�ϗ����2y�a���pO���f�#2�FG�@^k@�����~� �,K;�i9)jUN-ٽ� <�(�R��`#���y�:쎖�U�^F��\��0 h 1�H�8�>��(�Q[rb�\��>�Kėe^����qv�pra��;�|$�V�N�V]�]7�ʉ���������(�H&H8)����!J��!JRR�@�����J
)������	C�c��T���;�`w���=����/�;=��{��h��� S�_�5C�U�c�lC-P�1���ީ����N�T[c���R���Dw
��x�&���qDNv���!B%Æ�6>EA1/���2=�%_ݭI�!US�QL�R��H�7HO���T��u��u]=�!:���f�@�!�M9]4.[T�ie
�SnC��pˢ]��߲�[�8�Jՙ\��4�P�yqT:4My���m�&�t�V]u7�K_�%8��)�Ɩ�WX��#_T�d*�F��! v�M����@�!�T[	��q;&I{�P��� � �r#7��3c��fuW�~��cU��ꀫ�!w��̝�����5��U�~`k��z#1��S%�w�&�2�dP����'�D�|��2�l�ƍ4�D���TWw�ܶ���?Z!��r��Z�A���7����>����ZF����'�zn-5�Aٍ��QoT}����4���y��:d��`N�3��H�L��%��3�>�a� {��	�O�u0`l�}7J��Vh̽[S�6(u,�{��G>�y�)�y9E4�%��U��Ff<Mfkg�z;��L��rc�;�7U�	#�$����!NTRĊ��X�;�5#W��ʜs�q���v����T2��f'o�inѾه5,��-��)����M�WO#�Lۧ����҇(k��i���	����@�����1���T�a���z�*��p�)&���B���G��h�o{ٖy���+5��3me�n��������'Y�2b
��7��Vp+	����Z����[�S��J�V΅J]�,**N��Ύ�k�IW6f!X�
��jWϟvI����4��i���yA��l->\�����KV��I���}�����SN��;�h��j_d&�۰�rc�5<�n�],	�p�IS0�OS�*ـH[Fpj#^��C$�(m�Ŋt�&h3�V'��K\S�٢orr��X����]��u;F��ԪKs�J��1��u��2Yp[M���U:�Fe�ݍe��]<��u�
-S��p�\b��f�d��{G�x��R�w��2�

V7};8�P�f[�SF^n����nXE]>e6�[�uK[K�щ��L>��O3�Ĩi��	�X�5,Ӄr� Y��1F�	�4
0(:uX��	��"l`A<��~MO��{�>^���m�W>�8�����/��Y�u�t����9�+�BC����>�Aؤ�������sg��MD��hA�C�A�">�DW�I��<y���r͆��5d����s[�He�[�}�*<�=�������3F�q�w�_Y=���E�`�I�PvSV4��[���\��T,������KU��U}�ޥ�^WXo�[�"b
َӼ���w1n�N�������ސo0�'Ww��Y�#7ɋ ��e���p?�g�Qy1�<�kmѳ�����5
��Z3oB*n��Z:��.��A�wD*���`�"�P�NC�śjۥ#R�z
��G�ݮ�5<;��^ǽ�]�]�]Vﺏk;�N�8vL6[���R��K/v>f·�"V�wk�;��Br�K쩲�V
����n����Y�[N�sd����j��C���ƈ/�skW-�������8�L�b�w�h��ݧT�n�R��^�b��:����7ͪ9�y��L�''dtyT��[vx-[�w����m��۳l�\���i[��E�ws.�IZ�������xW�ncl�`�z�Bٚ�ad7��IA;9i$o,���8,�r}��n&x���Asd:{!�t�.����Ot�����m����M�8���4�\�r[�n�+
����x�t�J�{u\7kx��S�N�Pke'��N�%[r�1�.���4kˑڜ܄\Cs��!#E�$0�,h"���N8��Z�սxp����-�x��:���ëGV�:�Z:���|��<x�N8� E �	F���6؅,&�Jw%X��!%
BlB��*��s�u�q��{���&�&i^;�u5�̦�b��#ՓEI$�*%,���O�9\�u:�� ()�-�2!�iJ�U��%T��f0���v���4���L�iJH��aP>�M�9'��=��A�z�nB[p2j�&���2P������c��O�:Ur"R��IL��$�HT��)fa�L0��7PQ��Լo
hZ�����
D��;C��v�A�m5)�����R�E'l�!Q$��[(��i���:z�B�hb&�
i��'Rj��RQB��:i馝W��e�I	)R4��R��L��	����d��mTFE�D�j���F�VK��*#ֳdfu�ދv�PR0����/4��z%X��U�S�{��L�{Y=@���y'O�策˭���sHE\�ɆJ�b�X��Z����#�#�\":@� C��	>dH#m�	�-�޵��f�@	�$ �Q P�Q5*�@;��R�
ZSeUQ��_��g�~~�1m��~ �����n��)ib��^�<��o������{/�Ij��{O�;5���~4ѻ���9��y�y�C9�M�Lpפ��$n�N2�0���h=�k��575�-uw9��I{ld]�&�vg����0(�����<N)��Ӕs��ND�2���j=
�{�I��>t#�����&
Z�0��|�
x���.6C�}�x�'�FpT�]~�tk�Z!���@��
���3�@Yt��y0�Ո��;!�n�~Y[����KTL�]�d�l�:�������1.�L��恮�q��Θ3q�P��"�["�嘑3�@0��wQ���̽/,лc ���^|�,�����[c�m'����M�� �>9L���l����5�>(g�����0�5`R����E��c�6�x�9��j�T.���c#)���48fu���6T���;���ݔ{�D�e��PS�� `{#��5qǮ˕����p���~�\��d�˔�V����a��C���E��mE�{�/ߗı�3��o��m'�6��G%�ۍ\�31+=�2M��ss�R��\�3	��PӖ���)g*YuG�n��ö�o��3�!����_j���T��N�ɭ�(Vl�-C�'gl�/st�V�Yl�+4�ń��v./r���d]G7�cˋ@X$��� ?�> �`�;�S\��� X z�=z���z������ ����/^�\��,���|w��9F6t�n878���g]���0P�p�u�^K�ye����H��r���!R�6"<p����#:�M�V_�Pm/�YZ2L&����EJe~Ԩ�`�c�U��53CP�e�Ja�Z��	�J���۠9��x@UK���*�9�֠}�����<�qE6��Y��A�[�F��ބ]�8�`������z:SL���b4*�I�/'�/�z��2�O����-��f�Y�s��*Sf\� ��;pv����}�:�=�r8�}�5d��2	%c�;ݜ �m�K�QpҵP֑�)� y�cwр\����� Zw���sj�'����9��F6�Y?E��ӝ�J��|���us[͓�/��θFsC$�7�������3[����0���p�o`�X�
����uS���nhD{.�u���r�]���+�g'K$�����!-Qb�|��7�e/�{,7y҇�e��+j'���"9:�6���"(�Տ� ����N���s�r��n��jB�[f��GWE䵜3�O��P�	"�T��ʕb�iH�1j*�i����è�%�h��U��+{
���J�u�vpه�L��)L�]���=qe��߿�� �{�}� ��@�U$�X!E�L�W�u�����^����ֺρ&Ë"w�MB�<\���#)��0���9�ۓ�w�X�RL����_�]# dh��p�+���o�Ը�W6�j=�!�����(��V� �z��x(�|pa���������QdQ����F����s��+�9''aX�כ��y�"�y9� K�qq�z���&)�>ب��f��f���%��Nsj� �����H�kH��4�Cܑ�Q�@���U6�|�M�@���1Z�	\��G@�z��2o��#K5�· Z0y���a)?�N�(�~��(��a�-�X�	�j�a����zx(��1e�W�m�h�R��?
fӰ�9Jn�s2�0Q2$=Vl��{}p�|eO��y���	��D�����`z�> /���`@ϥ{�~����n7&������zF��zl�C�b&rEы$��"�!6��7��ڑ�^�g29X����KH���J���E�R3�3n��t6D���у�7�+y����ɝ��|8`�L��]���9}����@����\�{:^�����lF$�`<�8�j6��\h��z����a'�6��Ie"6�&���Ґ=��ogKu\�����%������"d	H�� �����)N@��!*����B9������W�����wsi��4����|nT]�7�}0�o �`T��H#������~Z^���߶m�H?r�Q£�v�^���r�i��PGq��u}�����.�c���$r��i]{$��q���}o;��1�&6��`tzL��V"FE&e����ݓ�>���������D#��"8ΰ�\��>���'��2�nFS8-:��`�{P�Hg����-�k�Q+U%�_&`���SR���}~���>�d����^-� GT18�ߔ3
bH`4g�����V�������u���|�т�n�~)ژc ���z�Jf+y3_uG�!�+m�]��-}�
��[e(n�v�6)���Pz���4�@Ɣ6�y�kgo΅z�E�4o`P����ywq!�S��:9̱l����h�?���1��x�!�B���i����q�x<�H�l���=�}�j[�Zǽ}�Cr%r�`lB�ɇm4<���ڣ���%��Y��6L�{�c�{�||��v��fe�b�7k2��L�6�d�;�)��Կ^��n�X���l2�؛���ac�1��0c� ���	�+�"dT )W�U]��x���m\u�k�k</Z8�U��o`��5�V8K���c�cn�S6�-���P�� ��0�lѭ��������A�A�;`W  P��V	U`�`��G���ԥD`0���w�ʶt������45��=�a��d�k5lj�Jw�@}=l�j��df�����0㰼bVF���½Ψ�9� ��[\��"~zc\�?/�������C��w�|7c���#�FÝr�s��(]1��������>��� d��ϯdڷ3z0��UʶiS+^R'�f��Goy1��.�7-�n\��hD�W�1�v�����n."N-|v%K��4k����/L���V�n,�z�kz@�~,��(�_ό���I�����k��0���,�����[��Ɠҝ���n�N�6vȣ�nP�n��&�0����ܜ�%G9C��"�䉷h��$io� a~���gg��Ě�B0��c��A�mL�z�V��1�6��������b���}zu��FE�ԇ,�ᙀ�K�-���j��8�?N_`���b��P��:�_���#Ǡ �9lsΟ��M%u��j��(^���1��������_p^�M���g�"e�|L�.�I3n�:<�c}�N�>N����_NN!j���a?U�0��:�kWhc|]G�yҽ���W^����nB���̂�X
a�ŤE��!������Gq�v3�#�ĤSW:&E=Z��%%��wsQ:�׈�<���{}�Y�?"<��(�J� &@��(�d �!d�U!U�O~��3����?sv�ƛqL�W�\��2���!�t�$���{��6��L۸��J����&;U�>��1~��d�=�6&o�B���R��AOM���f/�&䆬�Z�jV
f�B��v4������z�
�}ۈhʆb}=��4�T= Ozc*O�	G�7�4��D�y�7�mYOh�Ci)�p���A���g�F��t
�q2�!˟er�>�~�(@�V��*���uP1��>(��X���8r��z��qR>�F��tW����l�3�ð��
J���@S
�����j���r�G�\�}?^��lgT�s{�W���=VU*���;���#E�&���@�@Mmc����{�#�:e3���-����O6׊��()�g�$}�臕���^Ӫ2��!4���9ם��*8��S�/��K�� L���t@�sư�ź�yۡq/J�rB�i��|B��
�2���'�I	�_۞�hUS�����ZFC<�-5[��}�#�!�y��	��g��,�w����4x9�/S1��^YH��oA�*~ϰ���V�
���'}Z�����uK�p].�սsm���l�k��´,��Ż&��7X�
$�P�3;i�[W`M���&ä��oV�T�Yha�9&����/{�l���#3�h�2���n]^��Îu.�R
[����3�4lә�� �*�&H�� ��A"�A y�{��{����%vGqW���&�����*>���;�G�^� �;Ԙ�{�@��&�ux���tt�/\n̨yޛ�L����ϝ~ HQ�o)E��o�7�,'" ��ZI���~/��؋�5�{���8�]xK�~a>��R,�N��,�',�8��|g�uSS*��R+�B�г�i�V���Ȉ� ��ބ.�4��L8ދ*#�a� ��Vň���*�F���pӹ��m�����m�L=���`�,�P:j,�^8�� 2��N����߰+���_DEf�\%!��3�����a�@=3�S� +�F��E�P�q�)��>�=��Й�iE�h���kݤUXp딋g+���_u�7>�ڜ�+<y�9�zSmP�Z�����6�;;��Ǟe︝ǘ^�^"Zh������5��,]�0kVگb%�� y��J��J ��6�A����Β*t?�c,t-���Y�^	�D&9h�
r�Bئ�>j�^�D�jC
̔~����sT	��y�X�����>�`��#�6M�4��'M6�Ja6���Z�m�~��LD����_l�!�k&S�9��,,�9N���Ni��
t�Vf���$�N�n䧜 &���I�n�B�)Hw�杔���{�Ȧ��D��u�F�rh�0FC�z�]�~ww�z���Y/�f��H�H���A($�A
�(A2�� � ��y��~�~��ڳm|���e��=)�p�-�*���s����O���-��2��ۻ��WyL��.S��ԁ!�O@��<c���#a�h�xb�����ȃ8�+�i0)�#)�:��0pvxg j~u�ٞd�<��T[kP&�5�G��&~a~���n�X��ݨc�pj�I�OqQ�n e5[��
~n9РBƩC�4*T��>��O���/&0]b�5�0y�	yg	�h���y�&�{nR(׸��:s�*� ��r	C�<�G��+Sd���reO��/�n~�π���3�(��0,}�]������r�Q<r�b6�1Wz�5:wh"_ch/��c�)�&:���B��c�/��j�^ذ��K.����b����l̻BȆ{"4 \�KTo�� v3���7FW�KF�Y��{"����摢F��qO�.��p�hf�C�B���Qw�bjv��~˟wn˰��5�ӳ d�_�o;0���c��5��9x�@9�MAa
,Z��
�=|�T�lO�=�GuVtj��&�{�d�Z4��Z����x�60����7��9�ϻ�X�P"�8����!�I�f�.chc�����/�����'/�=J����m?>��V�-\��7Y���
KɅN����6�����x�!�q��ʾK����^^��_��{�p$V	���A0J��*�]f�s� ��$0����5Æi�CC���~��d�,}���4�y�t>�E}�.fhl@
e�/�,\�O5��=]+##oDZ�e�BW�t�f�P*@��"G)F�p:k[��#�{R:�� U-���i�e�d�2��ҦN}�P+Ƃ �@Odq�J� ���
�d/\��;� ����7�[�&�j��ad?2ӓ>�opR�g�<��Me}=� 8�h�}9�WW!��[ޓ,�m���Tۈs�ul1���s���<|x8@�'�~��}	ڽɞ�9z���;C[��G) X��> Ș�T��f�=r5�ʍ��Ak���||��W��Ŋ�!B[#Ýc���A���sS!��)t��:�G<y%��I� ل�iib�:�_��mֱ�������x��b�dN<�0 /]���~��ɫ�zy����Ke{�Ǒ���ԥ�t1o��Ŗ�@`�O��r�� �rz�� ×��0'��� sVwк�kz��A�vq
�J6ݚ�ȥ��S�� �����3�%�X�{|�iş�tc��c��d�)|R��3b1d����Bg)�u���>�]0����o��1Y��g�}�s�Ql�����0{[�U��#�D�y�<uW�z�*˶��Eg*�U���(Ļ�t�m�1���/z��|��U�n����ջ�=��}s�ۜ�=������R�e�� �J�J� �*D�@�tJ-#G�u�^��{���~���^�w���I�ⷒ3�?A_���q�g��J�<mj4�H!xޠ%��r/��
�L��&	�D,͋��)��F����[��ts�_1���nϠ�H��?�� g��	EE�1�C��3�����	��w'�%v��ks"&<VC�}�@��K�N��P�ݧ����:vק�#�u\l=�=%3߃�zX���<5`���C��\q�A�l�<�hQkۻ���������r�T��|t��� ���F����ޔX�P��X͝��S���dNYE�40�^�.Gg���LLmD|ᇠ,�
�������f1��ޡ����T�2/Fd(�,[��	 �/y�#$6\]����52��'����s�l��~i�;�N|�g�ž��/ܣ�q[t^�+��.\�|�'h�1N=�HON?F"��C�>r�r��V���ej4�ec���w�8T�f��g��b�S� `����L��Z�N|	i�q�چ�����ɂf�êM˻<��[�xG:ٻ;2�j�k�Z#�Γ�m�{q���H�F닧�2M�IEo�6w8���Ѧ*�,��'��k `�Z�\;��kvL�Ԩ6�]���B��%SU�yyvLW�@��(��^1�*�8'*[,����ݕ�,��a�ݏ{%*ꪋV�ur���sV@�BEc��4]P����J�k�8*�_fђ���=�wg�\�ӵs'SN��9��P�Q�`�`�Wԍ�^Ñ��F�Ŝ+"�s�S+d�<�h�2%��(��&�ÙB��!,6#�3�{��M��6��N����X�]|oBW�hkdvVmڮ���bU�US���S��!̪]�N77o�[����u�wM�u����ǪWh���wJ[W3��n���/4*Y��*���e��Sh�85Iz�'���ެ����ӄ���UٙR��N��Q�x�d]�Ƥ�1�e*U������Ɏ��<��8���:�svT뼅�G^FfnQ��u�IN�Q4т���͉� ё����z��.��Ɩڟ���YBVRr��C����7&�"h�����T��|��5ƫgb�H;�4�=�&(1 �$��!��,]A�]���|z�H��B�+,@���tc�1�;� p9
@��H1�����&o�����ſGjЍК$x�K1=y���b$���n�zP�HM|�4Q��	A�ǚ;l���Z�EIo�i��.eΊ��]P.�v\�b=O�Ӻ�p=�+y44#�^겑ϯ�ePB�ޥ�F��m:C��u!��ok%v�Dk5���VS{D#t����7V�8�.�#��gb���/�:X�fQ\��z�<�Y��c�}�o0�8�*��`�b�� �`e`�g������{35}���nW���Ul8t,�}�ȡ2Kݝy3m�gua\��T���G����VV�4o#8_UF�T��DWo%[��w:���T�7W�7`�ޱ���c^Ø��^��yG*VSrE'2��\E�Ǵ�����%6��ޛA<^�ۼ����Fkڙ�V�Y�\�b��.���e�CYƙ�_�paWU븬� d��V�����{�WDNw��WV�U2{�ʽ��2�{�O-��{O��,s��LEMN�,f��b�{��9{��P�Ω$��U�YB��Wx��y��y�|k�;��(<V!�5�GB�*��W.�l<S�R�۪
c�,��iS&�2�f���E�7�>G/BR�	^��b
FJUĔ�Ur�?0���}�jGp��c(B����,���r�����8ð�v�0��DJ?K��ER� ~�����������y�Uv$Q�(��
���;g�L=0��UWU(��!iI���@4P��(l4�a��9�����/�\���`d�$.%Qw�y�z�g�����������I�����`G�r@q-*w&INÀ�zt��:�%J��}R�T�'6A�(w�Jjh8��)3*�+���ç�tvP��2���4�R�H�M��V�
H���c^$xaD�y�R���������89b﷢R�Ӻ(�K�Oql�I�$��\Lғ��[̴�����89g�G��֟�h�rO��`�$$X!���`� 5 ��\�o���M�;|��MD�"#l� �\�����&Z5(��J���֝qv|�z�M�k-�����&��;��5�so>s�y��^))��1�8�k"Oh������iu�[�L0�;q��A'�+�	D�"=����nB��3��C�k0����j���'��A�z�,Dᖡ�C!�C g���Q��L�'�%嗡v���vZh�g�ѴB 1� A�~�?s��~��	�o!�����v�0���8��	�9�E�cBͅjGf��3x}@5]F ��OFZv�zU_H`�������ϕ�%���}<<V�:	��� G��-D��'�z³���	
�h(.[�Y<;���KHX���k��wy�eː)�~��ç+�!ǟ��H;����L�z)(���
n�w�X�=��@?����W�4@�g��~#_}���^\�jR �q��|g1L���V�_ry|D6.��*(`��a \�1|bM3(З��"��D��ݙ��U���I)��+%y��{׋dO1�y��En�wg�:�˩m�x�%b3�@�/\�����w�-�-�L ���Fӑ�6��n%>�"v�d��$ʻ�>�O1Xu]�?o!��;��k�n]Wrǃ8�0��V�K�+B �H 2 p!H%X%`� � �N����=���|���8��Ʊιod��D�q�&!�:��1a���3� �!K:����F��&�4e[������(�'����Tk[�@��x��mٗ<�a� c�w���^��$W꼮��u���m��0 ���=��4V@R5�ND&9~F��u�-zU�0�<�/&*tWKE9��|���;�ӆ�2>��������}���K WYp�mM�N�o)�%R��^m���r5�JGLʶ�ئ�u�-�5�r�c��#*��ܐ�tX,��L.��N�����l����jV�~j
�3@�n�<c���)T��5vo�#�9�'�5g���s�� ���T����b��dn=��_��R�D��.���&T)�ʺ��{cO�;k�`C*]<�n	Q�^*9  >�6�A/��llX���({%2��@q�grU玹��(�Q^�*��|M�"�3� |yx�F�����W(�$L��`�T�ʽ-�3*-#�hk��>�B_ ���lB~�.f��B�� `�ܑ�vW/�Tsā�*-_y$n'��m��^�� ��E�z�jG�v��	E�U�b�;��T!Ǚ�b��%fno����H2#�D���*V\S������V���K���qa�RM=�Ө�R�?0�N�b��+��ͣh*L�{�."I��*�k���w���ϸ�X�x���[���Ff����������T�x.�SA��p!$�z�m�J��Q;������1�f��8v�;�`�,(C��!F�c�P�C`�C�N�����w�97��=K������/���[F��&N0~lc��D}o����d�S�� "Y�{B1vh�]��@6�Z	�cJ�O���@�k�ū�ԡ�Vrf>�;bo��Y����X-F�/k/41����R�Hӟ}j;��D��ɰ kS�i�I6�B�9Ǆ����-uJ~\��NW��M@��|N��N���p}_Z˦$�Նl�=/�~0W!�@��Ɂ�ChNa�2>��ؠ���� ��:�YHoz���D�#��唆��ɂS<w�C�h��_D�2ƹ�����">�>�Ĭ{�&8��K�,�N�n^�u���������S���XA*1ׁ_�:r6#�!��2�~�y�Z�{w��opq@Pw��!ʲ��iu��c&�kJ7=�u�!��{�>����8��Ռ|��8�Y�a8�t�2������n��H8`y����M5��4�������tt����ƮԘfeF����+�7����uѺ���V�O%_d�&)1�:GqS��D�x!6�UZż��O��aZ{�ٯ���t��ƳeT�'5��O�2�Zq�Lč��u�Z�Q
C�t����3o7^���_�B)	MJY	�� � ��~���~�}u�{�:|?�&~0Wڀ��^�l�u� ?~p
��N�f�	vX���x�>0ƎT����7h�cj���~�"F<.t�y�4s�l��218����{���7�o��'�hD�e���yӵ9���.wC�h#�pj�480�ȧ����#s��P#Z�鲨! ���u��<�ʼ�A�5���	*E�% ��j%��ˑ�o힊�@�}#k�T?;�K�U�s�(�g^��&;f��^�fŅ��e|�� �* �$���w�t��\m�y$..x��ŝ:���7� ś�d-؀�9������z$Lk�.͆^m��;TL_;Y�����dNC����3�i@f�2/gݭ�ۮm�zS���?���W(����:�-�^)�������R�U��M �:Đ�|�4s`0�~�$�l�J'|�n��u��)�1���,/����Sr��#.��
�8�Lx��l�=�=�^i_�'RR��=[>���Y?	4�\c����(��l h�P��zQgA����j��������J}� ���L���vft:l��1M���P��ip�w@����Qt@!�E4�n��/�ۖ��Y����ņ�gu)��Tf�`�Nla�Ym�dL�eM�dPX-��ˎw���Â�P�N�xˠ��J	`��X%{8	�g�s�z̨?���i�Z��HȮ̉���`$����P�1U�̧��:on�j��vo*g��S8�Lrpk �ȁ�h�ZL
�<�
�@:V1�0ouF4Ô�mmN���7�G���L�lS���>_yO�6ۀ^C�t,o���|��q��.BG��c�M��B�}2��E�A�
���<�����2��b���tj��̈�������9�
�4��(`�#E	��%�N��inl_%�2���iH���)��ڒ�O�0�v��ԩ���d�zMoԉ� 4>���ͺ�@^L@M�6'��-f8���:§I�]��rm5�ݦ�F�T1R�`0u�M�_-a�M���l[/�.�a�`�T@,�؜1Eb����9�{�)���{w=���w��,'�֡���:���n`���LƧ�8�A��Oxz�{f��Q�%��C,ti��0=Q�C��G��6g!
`B������ѡ��3 �-w7�!M=00��d��M��3�u�k�/[�C^̙�(A�B�.�c!gբ���GڦML�YW��M��vA����H����I��&���)m�u�-������.���\�j���e]!� (��F��n�jO�oV��\��h��#�q;��y�R�:����eA�-�n��{'U9y�S۪���>���0�rB�9S��C����2��ٯh?��]q `Z�rd���� A!�_��(�CtP�[�q=��~�
Z�U ��2�%�/=`O���bjs«�?�C�+�� ��g�	��9���a�/�#Իi�W4G$���︽�E��H&|���{ԨD�H�_
�*W����H���Jҗ�6F�n��|�W�eS�)̳����9,�T8��&��P�T��#�`@����vVB�4�:(d#�\�T؆��'Ǆ@i��<��p��B���V�sh(�-�g�HG`��hy�l��ˣL�� (��#���(nyۍ�� �⍨z;�hԍ�J�f!ze&6< �6L�%1��<=��eL_C�6�F�#�x�j���Z��l*�GM�qq��ӐHY�S�I�ۊ�"S@��lh�Y��.6d2O ��K�� �n���Ϊ����U�.�,%�e��a?E�w���F(Z̡�R�3j�aS��tIm�G(��aC��<�iJ�����F�<���͍:�����C�����C��@t2j�r�BhӔ�v���U=¤�w�QJ���6+4�����:u��T��M�T�12����g/^ix�)Y�N��n۪G��u�W�P�\9�P�f���;�6n���n-�/{~{��ψG]�E�g�W�!	��&�H&&	�O<����ٴי)P� q��!�3�57���-����b�:T8���>4�'@{�oX��}9>(�Tˡ�'PP�,�D�o,mɈm^�"Z@�����?7,� ̵�Fۆo�il�L�z�aW>oK�AE�/�����(�S{H����sg|�|�%Pހa��T��G��*n�*���&!���X$9��˃Ӏ���ʐb�`�¯��N䎆��:L­��y&fa����R̍pGS	��� k?sc�ϖ���~csͰ-��HԘ���k�)#�T��_Ꟍ��B�L��3�D���o��ɶ�.	Q�͒q��Cy�T�=�z�K�ᑔ�5�v��0�\G��i���`|�_ �I��Y�2�O�}�(ͭ�(@�8Ԣ��x��_x3�0g���B���	��d���2!���� 8uD:���}b��qԢ:��)0��* �U���`�-|��ʄ�c��Gw�
�3fDD�JD��#���X}[UI`�ݝ����o�gvxT�~��W2�b�����a�����2����-�G�{ؑʛ�؈�ה=f�[�d�^�9*�غN%R�g$be	M��BDv|������׻�0�����+��,3�"C�0)�a�f��;�Xϒ����eW\�	��zQVU����i1L렰E�T���d��[{�e�9V�*�^+��� �����	�`�	}n��}�$����>T��n`���MW�7"|���HX'$l�z��r�^2X���^�k�9	�㓾���A�V��W{jM�;�O�Ћc�"�h2Ø"�_C��6U-�h7Y�&2�t�u���9�`��} ��/r�chF�#�Xퟘ>"Ay��� q&�g���Nj�;� �1�!�.�j�.�qz��/���MA쇫�6FVnt����ɲ"T�C&�ɨEq�n��>�*V�0Q����ZF�`c.���:���~�eg��}x�l�����ˇƅ95�#ƹ�7�ez=v�<����ھ ъwlHOdX�~���#A�CI�k��~�_��t���ߣ6>TW��t���PA���A7��ۆ^��a���:�������jr} �C�2u�$�5��?ߗ����:Ǩ
F�y�~��ns��QN
���H>�����GJ�p�K�0!4a�w~�չ�� �㱻[q�U��@0�[T9=z4T+���,:�,$ĉ�{�fs�@i�� ��vL�3�7�s�ɫ���.�K4��{�IZ�+������1���v+Yk2��h��f��=|n�#er��+��su86�x���;�;���&�y[���y����yqJ^�\�w�}�=�+�	ڥ�r��3{��}��@!+"��!dB!wdY?}�w��f-Q��T ~���a�f���g%�zS�ɂ��gO\��<xb頓�	���	��]|�%f́c�!߾X<|�S%z��~\Iy��3;�X#%��Z�$�v�F�7ր�����+Β�5�@���طP�Wll����y���q/t�#$���xA��Ը<���cc=ѭ_��h��J���E�� P�W���g�.wҖ�"�y�����v���2��.�^[�,�B��L"�M��M�U����9CI�~�x!��;���(ig�>���Ec���y�!�ﱹKg� ���q܀����#T�=�¼ءJ�;����5R�{������{ll~�c!Il��S�hVx=*��ܲ2^����3�t�VaD��bY!�y�X����F4-�����{L�"�P�>��\صyw�e_��?p�K�|���âk���f�.c܅���C�Bs��!�����L����Pzy���7o3�3���1k�T����`3f<��x���V���6��#��nd���<�)��������u���Q_����#YJѭr�Qǌ^��SKv�j��Y�^p  �H�����,Zj��b���uոYy���W�5�,vL�r��w�JS��xq�ݘ�n9:�㯅��{��� L @�Hd��\��׀"��|x�2E�w��X�~(�`��1�I��"꫽/r�VH�Bx �����m %��U���I�%�ގڔ�	���"{�cB �,{��=�?��wiz�5���\�P&��=�6��/��׉*3�NE�0 =?��^X�7D��{d�(WC���m)����8��",�/�#���f�\�,�):Q=(_P��,9�l�=ߪ��%-�e�����&�?tH�~L���\x ��HS
�CyOf��'��첰��:�|�ǚ21R����n�D�,��ˀ�\��}pnq���cG���F�n�$�w��K�H��0�6��n�1�@mLd�s�Q��8
��]O�����_x@H ��&�qƸ�� :�CO��pcD�+��Ǘ��ꌋ����r���ߕ>]���Vi�!5[�R=>�" y���	�5��}ؠ�>����%f����3�"�#�e�q��ry��N|����������7<�d�cנ�l\�m̺��_`���v5��%����>����a�ܳ��t�IJ�3�k3d<%�j2�l��5oUV�}�^�I;A��TZe��ȼ�y�������B�F��;��w�=l��V�o�Nze!X;��q�h�n�{-����ܝJ��� E�nfw�V�Z|7˜�TSm�zΝi�;�F^9�SG^n�k�BU�Վm
�p��MoY�R��~��:���2��V��Wϲ�Ɯ;`����u7r볖�ѹsŝr͟����<6���"�Ik����,�n�9^���4N=���D�!E���wv6fӭԡ���9r�v�Yz����C���-vrmb��Ѣr3�i���T%1��û���9X�r-]�w�k)��&v(��SVڤ��ڦ������Vƪ�4���@Q'p5��)肭���.�n���y�m�n�Od����ֳb�0�Bof��:uoL\�?jOC�R�\ڹ����:��g)�4;�VRV4<�[­k]B����Eu�~ਓ�c�A�A[�qt�#` ��EQ�fы�nrljj�{,�LS.i�.+�o+�Q׍jݪ��A�w�|��GyZ���U�h�3K̜kN��V;hփ����诂��5xt對ky�X��maaǅ�.��y�t��:�w���uv�;8!� �X�]� ��dU�0]�d����v�vz���!��c4�HLMT!�QA�$S�@��,([�h���4*Z�J�;�e�c� �"9nqLb����?("J����h��h��!��'�+�b��PZ ÿ���X{��saH�'B�GRA�e�1�	֯*c�·Q��B`��-�z�n$��dԷ[VFĪ�&�n\e�".�Wn�E�'zvZ�}��������I�T2���:SQ7{�`F����(`&�'�mժS�+T@1�F�J9�,��˸L̫�$Z�u���y���ˡV�֩��FFa�&�{q]!mx�7�S�܇f��f�a����eݞ��wi�(�<�xi8M3�Xke�
�AS��w��7V��W^8?�u�F��WT������!��z�oU��}�^�Ŕ���{�Mཱི����,'Jȵ�]�ˬ��ǁ�y��1[���Ȇ�LvBa��TAP\4q{;�_=�ay���g;���V�u΄��������������κ��)5Sf�;���T�0���+�f)f� m]r5K{/k�a���Yk��)�q��y�N5�tηW��7=uf�71�h���ɥ;K2�}A^��^��6�R�I�ӓb�f����B�\����T�r?<�{�,���{T�iAch��3�S�(�ut0e��O_*�;�ʣT�Q:� ���[���umCF[����q�խ�<q�8[�^>u뎵ou�׈���u���"+��C����qj�u�uո��G�玺��xuň�,��DG��ē�s���.s�(�P�TF�0���B�mH�6a��-�!�ME�K�Z�n��))�a�����%��7�R@y��8B�m��h����R��<?���bA$��C�&f&@d���2��E�.IW*B�I��t�ᦚy�O�fąy��y�@�C$�OaW*�*Z���N�<4�<8Rd��'�]Hj���� ������ �<����L9��eT��u�d�$Z)�,̆�8� ��<�����i��ȯ�}˥I%%�ȥdj=�N#�\�-H��ΰ9?:x~0ê�*��H��,F�$2L����XS�M�*H��M4���M0�ǒ���F:����DZ�!�Yħ���������~��$��Oa��	��5EEMj���(�;�F������!2�h�2
����QMj �\�  Z�K1��>�݆|.�E��$m����CMK�E�Uզa.��gxx^�]��;movE�ɺ���Π����T���*�+��@A'���O^��<-�Z����H����U���B(���*�f����,�'��ܻ�����00�#�	�Ym�%Z��f�P�K�b��1���o�z�Ƽ)�u�-n$�ɩE�H�:��l���������͇u!8��g�B`@�T-��1�[�h�P�Z��[It�@�vc���S�\c}Q[q�n�,�o���w���.hLE?�=2S�v��G�3J�ы]��"\$�_?���kj���J��P��H��s�(���2m�1^����I��\Ԇ�-�D� ӞQ��b1�td8J1���;�=���4�`o�Ѐ�_L��w��oJvﭼ�|%��kvy��*8��屁L ��H�H1������$�[N~��O
H<����� ��U���ҧ8Pϟ�gkցI�װ{�3��RE�Q���yqu�OkNŀ�B	�0ؼ������$��)�U�G�a�c���z�2Կ�A
��9���@��B�C��ʉMc��;36O��a���!F�|c���%:T��w]�zs�y���yTx2�/�����:`	�@�2f�O�I�> �޹�$wzZ�\m:/��/��-��i�L�M�W��j���)��trv"{��������Tq��i�,��rڋ�{���!��{�Z��+�kZE�I:)���s"rb��6N��w������6ޭ��j��wbfY���@���V��߉�͗��z����FkG`�"�\g��/�{�KI(�{�_&^}k[V+��[�>��>�jt�w�����0� �?l�,l2��hFm �tX�%�����R�p��պ� 3�!sy
��I "�=�����%?~ί��_q���,
����\���s�e)�NǛDG��~�&���QLT��4t��H�!���q,X�^%����ף��7��l�םr=(-�w��pǢE�x�/p��A�:�� �R<U�Ǒ<�X�j�8fY��Q�&9At@*+_�a�M�R�[���ݦ��v�{@�ف��hj2�R\�g�Ɏ��`YM%<C��SP�� �hJ`-�yK*��Ѝ�xC׎Ǫ|�l aS�u1bgp���u�.r(�r̩O���ҹN�q��w�FƉ)<�4s���T�J�`rs����:5'ѧN�c��0R�d��C�bҞ4��v�_6ak���<��1��v��<���4�������G>DA�� ��Te�4��P%�
��zP�5y�4a��z'$��fL����+M��{f2l��T�Cqȁ�ýɛ�z��cT�����x���]�<@�隹d��e��~���C����_	b��^=�es̔돋��Vj�;����r�!�2�C�c2�D��i�nU���K�;��-��0� 0`���]&>^�O�e�6�f��c	�G[�G΋�sp�d�Q�0A�s��y������5�Ͼ~�o�O�}�R�Љׯ	c�X,����d#0�'�eںLz���+�n�����@��A��e	�k���,��� �O��3�>ߤgX��Ts�
�T`[OH�.��������e��'����RVƒo�$�E]��>�@�bм��{� �k��:}ʽ�Gr�l�G��b����y4��������t�z�;�T5��4$9s�z;Ƴ��/�n���4�p[��A� v|ɯ[�8LY��h�̄���_S7�X�X�wt,:��~`+��n��!������*� b[��X�XF�Џ���]�=���7Sˢ�2%��M���6�/��4�ߠ�okX��()Q��q��Y��=�/b��r��m� c���1�ܲ�9B������|W&b>�˷P+����fA��Zϡ�R�@�u���t�M��>�-�6S�qI�f��V�-�����}-�H��ڏU4�V<yk�����,\��G���Q���ѴqZ+AR��V�E�Z�Aƹl�[GL��?@@cu�R�i�t��k�t�k��Ab�2���ӂ����.����`�ƾY����ٲ	V�񾾯��� &Ѯ�D'�|���=�t�ɥ�,������}ȥ����<GθeL�zձ�*��U�%�s�nÝ" &�0#�N5���E�h*��� (��˟��g4��u�Q-�����/:T���g�ck �VVH�'<�kϓ��0zfo;Sr{�/=�(��͛;�!�7/P!y��i�
�؇渣�25�GTLa4>9��)�Z2/-�T���ZP�=k���tbX$zq����h�?j���Z�zb(�zj�mq`������͑��Kq�����;�I./�I�^����B�[�!�(�#	�>���w9{W�w5R��ye1�[�0�C-�4�X/ 3�q���� `.d|%Ď���6�q�|�(��n �=��Py��`�Z�=sLSׄHbCC�ߐ����	���t�ڃ���\]S��C��̓ȇg�="=y�A#�aXVz�<$�k
�M^��Qv\�S��F��EO����5�`=*T�q�>�v���������yMy�%��)�L���š�lp�b�w	�Q��ud�oVYpd�:U��[�>���T��]�{��W�jE�[�m�Qi��7�';Il����U�Y�v̤�n�r�Jɗg]w^n�����XXJM'����䰯1��Q"��B.[���jsz-U�{�����^y׿]����*ŀ� �h=Aˁ�$����9>3�,6�C�M3���@�M�1:D`w�`No@�C'��T��p[\/�g���A��0d��>Y���0!�t|ܐ��W�h��>�#t�D��B�( ~2��:7Օ/���iC���7����@x�'{>��p�4�X��uR��v<��=M$��4j��f�Q��O�1����I��0��oN�k[�^+2ş	s��y���`���k��"X�J��
#�c��#��U8g��t/!d9���|�� ��-�z��7�=�c�m�j)�i�b y64�}rD�%�+3'�OR��ʻeܱ�_9`�����4qu�>ޔ\��xe�ḇ���G	54{��5�&��!�%��ltë�t��_��1���9m�[�*������� ��7����u#�q��{z�],A�H��VX}�L�oH�MPi~S���b�̍�)�l���Q���2pv�Z�?ol1%�f���ة�ٵ"Zil�Q 8J ��ӑ��cL��^b�aXz���t��*&1#5a�qYx5 W��w�� �Z�=;%:()P��۔��Y�W+g�P�/�RY����gɣ;I����3��4���K*;������k��9�k����6���$v�-�ۙ�:v����@�� !�%�}�j�����������ã�yh�ң�y�J6�J��g����^�x�0^H)�mlg�U�:1 58�?7���1�z�I�K�a|i�e�Ȇ�[�{���"��FMe�� ���:�F�92��W���!����HO��+��ɵ��f�a�ԃ��&ƟvlOv��0����
djH��'����C˿~uqx����{������͘��c2۠Ar.��5xdp���{F���טxkhg�'���ȁ*id�Wo,���8������v�b���O��y� (���b6�:";���[>݁�O�=ÂH��0�y$t�{��@��:	��*����ߙ �_"W�v����uF򼍓�6�M�è��#mW��-]��Q�:�_�2І�>c��; ��*C�����WU ��ך��[kf��l�/�K˧hi��&!�@�Q���<e܌ˌ�^FtC����<Oc=+��-��o<�{�l�T�=��a�� �l��]0Y�@S�{H���6���˸��qor������j��!%9Ы�2�5v zmU�m˹76�EU���,u�ƹ~��H�{��r�Xt<�y62�1����ţ�����9ka����[P.ݽ���d��F����f=oc�G�:�(_����?q�N�M(��kS�Fk�(sJ���&&����ɦ�7/�E�����ڎ͖V�~Q:���J\Aِ=0q����e�����d��}�	8��gVN�v�اo������k�r��z�@��Gq��f�������P��ה�k�w�}�nO�u�1(��t���^v�wna���(K��A�7�A:}��z��*���_D�G��$bd�f�p�4G�"!��܋l��8���|�sa��0�� ����|љ�����$^��5�[ȋ�龊���}Gr�Ä�fǫ �p�uޟ���ķ�Y�8l�L&,��q��)��IQ�MdI:M�n�fO�'b�~���c"�^P�U�}�(�@tp�A.Lf�oū"c�V*t��緈�A�v�ց%{i��g����_7�X�,$&9띛f�^�ǘw�<�.��z�ƤP�f���!�)��sY|1M��~/1����-�K�(�Uvz<����m�=����G�����1���H�$/:��!���^�ꦋ��C�~<I��,�Qc�.��'qA��v���^]e�t��#�9��n�+w<k�\V
͗>ͺZ��J������I�׷B� ��e�� O��9�����{,�R��U��I�W����ުe̢J���d�8B�7�>�ٙhޣܹ}�1�O�]A!
���{�~���z>��:���z[];�˛�|�+�Ϡ�ɿB�N?܌�����>���MtP�x������Zb�߉�w��G���f�`��t��6<�B��n�q�8�o:�2)����@W� q��1�VGȫ󩘡�`�e�?'��]�<;6Um�f��a�)���yR��+��<��Oz[����H��}�1z<���1��ن�����+b�a�q%�4
�nl}�y|�S⍭�z�-^P��m�*�:�3~r�9|�����>������8+�3@J����Q�`�6ȹ��}��u��=��&�;�i!z��;�!��0rJ�?&~�X�~_�x�D�؂�L.��=��(]͸��su��~|r}�~�+��PuV(C�L\�Dٯ^O%�Z�:��̚���#����i��*�?�G8u�m�C]݄CC>7H
#�_s$i`���܍E�yf�*�s U�B�qqR� ��c��\���¡�j��n�!�_-����=CbP;�
��Y�1�p��BrZ��wwһ�c�ٵ�6�P�q���A�]n'�ܜ��=bp�T�H��Do�F����E-��L#[h`�X���U{w�Q����;WIT�҂.�R,d�M:�Έ�r)�zmk�x��qC�Rݜ�}r��z�H{��
�п���[��Ø` ��>^#�q�7�q�������dl�zF"�e�.5�z�e��>��N΅j|>������qϢC2#�vx���;a�>0�~�+�R!}�ƳgL`�d�-���}�Ovm*u}b��lLO���K��5!��G�,��3��q�1e�����hQt�f=����KJ*���'���4J���*lj|fǖ<_k�����-���қ���g��%����	��� �9�	�=ѬRbY��%��W�yfvD�c�(�T���}|�àcr �`���٢��0!�?��o�n���ؕMu+(溶�}~�"X�ƋyO���ݎ���3��ذ{n��n�z��(�Z�]߻'���I��G��L�(��f��|���-�ؽ n%�&q��I�b%�׼`�1V�ZG&�c�S�HI��jf*��0}������E���{���#�1��Akr���aF����3O;�9���ּt�Z�%tXz�Qy0/�>�8� ����Zh 2He{�3±CƼ⮢�_�,騑������YU�i^�s�]؟9��\�q�w.����܆��fq���< >�8�!��F������+k�U�w[�L�`��A▥�N��3&!Z]}2����b���­ɗ��ˑ��3I ``<��=ٹ�%�E]���*���H眣y���ހ�����z@~2�����Iݔ%��!��	�-� 0�^�����?6rSB��ͪ�3A��������Z"�Y����j2~�2Έr0�&9d�O�D KyQ/`(�e��F���\�:��f�)��,���:)nvW�.���w-��M�@Tlʑ-K#�}n	�Tsr��)��\fٚ�y�i��Л����cA��`��w�e��r(tǝ(��Sxn>�Zi�8�|Jac�e:��ܳ�f�pT��A�,�=��މ:o���]*8H����ɖ�r�+b@�"B���~�_~�?W����`Gt����� >D���D>.�>�Lբ�ktxZ�Br����hn�@����~O>��>�������`�+��G ��Q>(��w�j�H��=�ߟcOš�?G����3+�?\��ic��K�F��Y�'֍��X�oޘ�"���C@n׆#)�����+��s�`D6�8Ȑ� Ӫ�;���x{��޹�l4�W�;c���*n�ҋe\�!z�d-����ِ�v)�����e�0�H�k����EK�ۛ�93xq����w�މ�6��WP��|&hЏN%q\���������U=C+S�W&�i����^�C�9]e�J�u�r�I����T3!�z���i7:�`ۧ͜�R�x�����b�Fdyм�7[г|tu��-�����`����%^<[.������\ǒ�g63N
��ђb����ۙ.S�a�1���j��'Da��)v�VW[���ܽsgE��r�/:���u�F���jkιf�{V�Ҷ�o�΅�����n7�Vj��i��a��v)�q�f��f
2�
S�YL�Xt(q��l���e�;}Q:�+u]\nZ��m���l��߫�ʦ����3�lM*A~��{��Ɓ�{0��^��j,�r���AK��bj�(�0�C{Xhwk��G��tOc�R�j�c��U!B3]��O2U����K��ۡc�-)cf�H�r��/l^���=��߮6Z�;�՘x�h�����+L�;:ڽ�Z9)�U'՚�b��Z�V�;�	��C��l۠N"�3kF8���q)4�L���!�ՅO\�`8���ʮ��c/$�����ݷS�i12�6�XP�Ǵ� d��^�+�G hN3	=�O�i�Ip.�h���z�E�#�8>A@����B�����b`DL
��	�LZdP?PR���c��:��f��"Ș	uX���  ��X��B	��mN �A�""��ãI��c�=oύY[��v���р�⩘A�q�����7���+3k�H�ݘ$��cO�`���v�UN�6�]�b:�Y��]/�9�pCW�ZT3�)�k(Z���]��+5����(�9+npa�H�MCU	D����M��$��InK�Tu�p��q(,���CF6�f�Q�g�E���gLd֙�X��\��)��XUʰm�8����rz�]!��Ƀ��^+�ެС��Y-�1���R�����Ҭv��)NӅqSU��x��A

A!�E��k�Q4�em�L\4�K�OZ�IC.ќFUE��`�de��d�u�&��O%uڱ&���·�Y�T�`78m�o�Sf,xsk�1�N��*	�[ �мw�[��فa��a�Š�i�7��f>���`�)r}=3��b��[���P5wy��b�Z'>��D�[%�1e,����̭-�<�l��lfģ ��
��V=�v�,���R��ZE6D��ؘK�B���0L��b���\��h�;z�@�����b�L�9����S���Ő���p̈m�z[���d����ηMn��}����";0�5a��OP��7�f	F�sX9e�4yk�F�������ç���<I"H���I����ݤ*�@w���\�r�!'�L<:xa�؜Z%ʞ��x�Z�)Kу�[�(�hJ'��9�Á��N��$��y)p�U�I�gPa%�b�UBr�`9!�������W�IC�NUW- Rj��!�&��fJq���������~;Jy)�ۗj.H��"���&�f4PUceE^_&�:t��M;<��I+��@�Pː�E"q&EAr��������:x|`�8������jre��+��P�AJ`O��pÃM4��I*������.�5d��T1Pj��u�Z������Ȧ�Y�a�KNu��*R�Z2��aⲨ��D�,�����n8YS/6��;fqKy�I�9���[3�����oXh������� �0�pG�**��/��'z��V����T����mgѝκ1|�.SWL'����>�u,kCz�iz������G� 0Š©�>F���M�ȭx�ӭ���/!�0�����/��?YI�"�s�J͏��Z] ��d���딇WmEm)��@1T�Ǥ�^�Ȣ��b�m�R�����᦮�8D}���<�-tN��I	�UMnN�V`h��b8m����b��
����B�^��&�kj@k�
��@��N�K����e�^�i��Z��$�'g���O��[!�$�Ż��1��'�&F��7d2�x�f�_f�n�T����|��\��3 ��>茻��)�����VS�T%:�s�ٶ��ۼjܱGb)@p�o�1Я�H���	�i�5���:�'.X�@,<^({�f�*b�w�H�z�xk׷q��w{`��>K�t^���'�㐦����l�\I�J8�}d�^G�x���8��w}�	/C���'��ڟB.�����3M�WZ�,)�Z�U~c����1�"�>S�5u�o&3L�W����li����A���XS.|��wώ8��������J��Jkd5�Qt"]q,2�V�p�Y"'bz{�0�x0fܶ^�jJ�����9���eCz��p�:�Ȇ�Dy
冷���	]3K��X�Q�γo/���\h�O"D�uo��i}9V�ͼ�]��,���)�^��*�fV5�+0����x���I��z&0H��t�7�Q�$��`�c��oDC6��&69/L�ƙ<.�[��g�|z�|T���	�a	 ݞ����RFR�C�d����s�i����k�Mv4�q[?�0I}"B�ޏ����jcޟ[�^w=`�m��wmq>1"�1� ��a��KIO�����_�~�	���)��x܊�o��DY��:�I���za��nC(yp��n���Q��Φb��S(�-�y�HxM�t)�����KW?'���	�O��v=�M�;Y#	dޜ����rn	!9R�<�t��}���qx�ou=���q �Y��f�H�;�{� ���=z�M
e�0�#�WA�C6��з�qL�\����[d\\ᚼ�z1�������J���4�&�Q��V�U}P�I��׷�����Ď��Q��/׵:����ćT)0S~���NC$ꪝ��3������s�;��DX[x�cP&^�v��ـ�H��]�J�F�g8XblT�pk��+o��":׋uur�9-�O<�r�/�r�F%�����(�pM6C�a�N7c��ux�b�~��3�N��{h��e 7�(S�e�C4&C�f�p��E�f9u^�%�0���EI�^���*{��?(�����,D!P����5�֋�ֽi�e\��_U�-�C��6��ԧXq���(���%lSkP�އ癐b*$Ül���"+}�7�v���uʀ��ȾT+Tqq����`��|0��ⰿ�	љ�=�s���g��&��pY��4x?BO�K�)��oH�U�v���z~@`��g`q\���X��{V�ɘ��k5(M��8h�}@\�,���8�-7��d؄K��4�M�<OB�{u*)���6'�v׏/ߨP�Myʢ?���gkߟ�z�����sȬ��\�kA<ǡ�7Y�~�gy�xg�5��E	S��k��N���
[�6zZL���=Z���ɹ��=�c����e�tA�\+���+T��-������x�-{Uf]Ob��MF�˫����(��N��4Pu�N`Gr�!��Z*+��N����,�;���Vh����u����V�0�F���������4M�Ǵ	��a�R�Ne���ak\}-���t�ܾە��q�!ɻCb�N7e�	��(l��ںͬO4D�4��	�b�pN0�b{�3�����F�h��JK5|������H�$P��Z�C`��t4��YB��˱�dR�2����En�{~�������ϝ�4l�M¤�;�a��%ת��`�ʚ=���ڐra�4�+�d���xn]�ؾX�d3��� �* �"c=zG��?eCc��³�{��&�A2c�;�X	}�H��m��( �Θ� hY���A�X��	�;yǼ^	�o՗����B�-	�J�7vl�5�]Xs�(��S#��?	��� ��^Y7>�%g)�=6���YFt�΃�8��R}iJ9�(X��@f����A�L�*b��/x����N">0�~��c���;uҞo_pM"4r�/@�k�ۤ���]	�n�<��{yq��E%�W�O����/�z�Hr�?x0����[�TQQ�آb��E�ֻq���r�< �-2@�{`��]8!⣏-B��'K�?g)(^�������(�	a;�*��@A���V��0,�PTP��h�����{�Z�g};��'���V���T���%�^�F��c\�߷� f�fvKU�c�T���du���ӗ��JH�=��w�X��_r�[.�+NC�獒������k.��*R���c�uPv��]۝5!p+�J�oD�ͻ��P�S��[ �f����1RAo�b���s���'W�������'䉶o,(z@��7xEC��uX��)>�1~�]�mk�ޡ����ƻ6��ol�^2||���5�o�L�r�y[�V�U���K<�$�OO5	qܣ�0����H蒢��� �%��I��/�ʅ�3p�"uӻ����,xk�:QR��[���-�����x�9�H�q�����·�W|����0���P���?�{E��B{�	�jycc�����������QW!�4�M�pQ=�~����6%G�Τ�ޖ@�*�}��.�0̈�PJ]"��MH�\��D�;-
�;���f��5s�&<ne�+�&��\D�6��}ˣ΅�|�Bz�If�٫:k��b�C2�<m�r�^�Ȣ� ���
�u�ʝ�y��=������]��}�0���l�`��=�$�6L�������o )��\>��5�������W�3� �{h0z	�KS������V�5���u)�<<$�X�n�mYͱ���8�̡�����Z��PTp,�K�Ѿ�aN땴rCԲ���k?t�o��Yr�ʂ�T�]��� ��B��%9�k�7��W�g<�l�F�7W��N�*�R��45�w
)�����ث�2�a��%�U_�Q A���	 ��?:ݏ���U�F�b��xC����C��������Z��˹��Î57l! C#ua-;������l��^� =�4������]<.z�MƆH�{N!�g9e�/�-��p���G��t.�Z���(�z��"[;�]�C�fka)G���Bt_UH�#;�nQ�����t���g��nO�k�o����JX~#B'_��#P7�@����>(��v��^YK��Ǥ���#���A�[�#���J=b��xu���P�U�F-�4���w)v������?s^P^ ��	�2�ό5�0�(�L�ZBˎ����k�]��8m�"ˇ�/|�!�N.���}V���A����t,O�2�Y�=�>���Lѝ��ܩ��6Vs�vE�����`~�tџY�W�Q�^��s��c[3."4�tOKK�~;�MQ_� K���^��9�Y��N�6N�bչ.��-�憓І �y�Ct7�)ﾖ���5�{����߆ǫ��0�#t`S&�T��(fT�de��Ö';�$E�Y!��Rͫ����I��i]��:^b
�42-�%�BLM�/�ۮ-
���/��^$۷e=��n���7OHsmi7��k�9�jj�ǱcY
�cD���㈇��]t�ܝ�s��;n]��c�H$?�,���~���}�����4X A@�&$�0A�y��pR�,��TC����kA�\���z�V���E󩘡�c#�Q1��x�v�v�[=����H�0��x8���	i�ōx��H¢��te��0�/D9��c	*"cD>��N�@(+,��?��\xt��,c>9%y����9⭸�M)����.��.�m\��ߗ�� �ˋ-HC�ߺa����u{$Hj�����Pc[�Ok䲞园X�F��v����^[y���"��f�cu�B�K��?"p��~�?/ƃhL0�����COdr�t��-���R�iR[S��Q,�1�\��@���=�,&��r���[��3e�4k�,�e��.(�������k�����d
 ����_hT�6H�ʓ�^uy�vo��4-����_ۢѡU�x��y=x%�2�RXN!s�",����ֵ�(�(!T�`O�@z�܄<"u�46�y���%��sz��*c�K�HP��D��^��{���G�Ҏ$s ��6����r'�%M7�.��S���@ݕ�j�_�	3㉓�^�QX�u��iF���$p�D�;�'0�SN(l��ͫ�̼�ɧ/h��$�1�K,���#l=�5Z��ԅc9+	�چ�M�*3h�m�c6�[u'ǅ;����fu����[�e�bȋ�v�l�?�@� � ��ի�,�P�#�#R��� �ȁ<:6q�&���(�-�'�	�D�<^r�7���#s�v� z��؟=�W��4s�)���!aj���r�GRӋ��W��W��h�Kf����6`i��\V�<����gq=�4<�l�3��I�D����MZ^��.�	��wQ� ���~��E1#y,��ݬj�6l�z� \��]]���g���W9��k���y��!�^���P�v��/����mf��;U�� �U��}V @��EAA�*[�#�T1c�
�꡺�c��*�qx�����N�����}�a/{g�d�~+6
Y�j�tK� 굶��?,ͻ��/�����yb�<��J_=���� +z.�ӽMh�E�ٺ��V�#�q�=�9����'�7�5��O��%zT�S��BH�A�m�r	��)�������k�Mug6�Y]�U�h����~i�0
}\��,�ʚ�p3�@J[=3��LE]Ҫ`����ikN�0J�mT��sgWrc:��Ef���ky�ܬtD�o�bRJ���!?Yp���DJ�h��t���K�?�s�O��
'�`龇 ��`����;��<zV�I��N8eB}�[��a�8>e�<��
��{��XU�{5�|_�}ǣn'��p�}G)��>���w�Z��������o�ZIؒ������!|dj�;޶ \�07�HG��u7Dd�޻a�a:��7�YyFYg3CYV�M��G;��;1>��{cD��5��2�� �� ����k����C؀(E��U�;ٛ���D�ס���<���82���ܶ����Ck�"�'�>����9��硵K�<�cR��%�}��{�{����JĞܷ�.t���{��v�6�|	��"r~�R��M5l�������H��LFH����^�`�7�d��}�4�7�|}�Ki:�ܞ6i�Ljr1�SJe@y��2�Ũ�w	���;��̨=]w���f�h쫈�v�E��	1�������lm� ��i܆�3̮�2몬Ԧn�̾�*���
�w��85#k�ޕ��k~���i�������ns��uT�w�\$����`�gv���*>�Ϻ��P�dB�g���ݱ�͛U����1yD[]�u�l�з+��Se+5�ycQU ��p��My��C�E�H�{%^��@�`�$xbj�^� О��ݯ��%�rP����c��(5��o�tt�-6��ʧ�n1uˑ�Z�[ͭ�In�<�.��2W6_�{�႗��O_$w z;6=3�����t��TKxIS �d��Ęp�ׇIm���]j7��k����\f�#r`V,Ng�J���eSJs��ef�� x�W���
�zМ��=�j�	o�ޣ�eԿ�'��u����]���K��K_5�,��@J�x(�P(��r��|��Fl�I*%���VV��c���6���e��h�Qi�?+}�x���>��>�䐜�=TR|���=���7�@�,��?G?�~L��u2�(e�6���֋�o���v%��ܮ�Ɇ�Zb���Cvc�,n�-�P3X���tv-��"�ba<U��j�4�,�y�7K��U`[)@z"V�UY��ᣗ��ly�Ã��r>fP�9�;�nn���-�qK���c\�p���zW�sY����n\�6�0W=���U��xīth�U�����I�yux�2�j�T0�9�������³zjws�N�g!\,�K���Yv�8zY
{ϖJ�3�|�`��!O#��z�Uê��of*YS��6cL�sK��wu�ݫ�Q(�wM�wsj�YWLۭ����m$�;���[s8�ΙH�Xڳ�x�롢V���Ԗq:�sn��f$�ӭ��Η�9a�Z@��w�.�/�����|�4�bO���$bhp��H�r>Q��^5X�i��!�
�]UW���P%�R�6U���L:�.qʹd�aUl��062\ks1m۫Z/�ݬ�W�Q�%�*6țz�[��a�ȘD��N��;��{C^�uM��PbU�[c��{�����+��w����hd��En�����g�鄩�}4�<���*����U���&�VM��{�:�ZMm�����k
��b|�5��,d�X�\Dr
JoJæ��s�E�4�䋌n6HV��ci���m2(�;Bb��;Eݩ�TS�!�Z(`��j�X�u���H.Iu�W�+�#H��A$h,"�z���>cFz�E��p���o�W�L��.���+��
(!"���}be��B�t��f44 ~����|�Mn��|_[�!�fUM�"�B�(��7a�\2�z-�-]�-�������U�~�%;�Ot��x_z_�5f3C�g)V�6��)H��B���e���ݚ��b�Eӭ�׼��2�i
n�zs�NR�LZ�e:�ع�݋�s�W}�Խh^U�����lU_j�if�lb���W�n�=è�)9��T����-�Ĳ��ո{�P��En��n�{��|��n�tb:f�e�0n1"���'N�t:��F�)���k��_N�L��Ni�q����8�Y��W+���;�[^�Ȩ]���c�7:�S�� �״t�r�d�����\�R���q ��k��sT*�d�V8AQ�98t�X�t[��F���:ˢރk�	)J��;y���j��n.�עq�kY����:�]9��,�1O2\W�E�qh�v�Qm�Q�f�(�ϝ�_=j���k��.U��Ȧ���W��.���,�P���;�NV��`��o&;��*\��f)R�n�I'Eķװf3c��LY�[�YЎ����WT��oe��s�,a�1�x�2�4�3�oa�F��0��(
$0�!|����Ǫ�[�q���GH�8uh�Z1�p�C��㮸���N=[Qn�G�!  �|�a�g]Y�BaM+ƣ�UE
	��H(F���q�w�7ɏk�|g\�̜��C�4�w�@TI���uURR��W	$��N�t���þT��ʒ�(

:�u���z���I�q��F��"��OM:t��<�^J-�(f�jL��#$2(�$�p.�����a�yG1�+S�Y eORd�	W�x2�"����8�34!�l8��6�U<N]ϦMDLEM�4�d��م�I+�M8t���N�W�\�32����"�rD���Q�Wxa�ç�aﾝ�=�NXTELDHVBe�1�J
(��,*e�C��t�v��QGKT��f`��2*�(�ɧ �r�){��8��;)�������SEFs�S�2�+9�KT�����*)*�*""i����xj�QT�ESUNXUTQUE�.�uF��f��Dl�"��q
��ޮ�����6ғ�.����d�[7&�J�[R�1��coQ+%`����=��f�������-#���]qn���x��<qe�GqdI����H3I�"d��L��'�
>$�|]�d��-��`l�YM���x�����	��y�J���T�id9�@�oxt8�3Vج���� v�uP�t6)�l6xsǡ@u5|�+L[T����������T�3GR,��[L��a��"�xc����a¶���ә�j�^D`=�'����X��k��&{������I��/�_��$�B�����,
v���z�X/�t�o\_��:qݰ',�P�d�o;��br�����R��*n�d[�Q��7�3h�Fb_ͤz���S;n��e��]�b��߄�C������r���fu��'"��b��8�M*�n6�Y�v���w��G��Sx�KG�-�O^3�?L��c��&�s�/C�,�,�J4m�m|o��Q�<$f��j�n)�WvlBz��yT-��bq��XɃ��<���FCp����s�Z����'�����j訒aa�:ʪ��D�Jl]��5pHA�ۃ�wrr��=,��7��Np/�nQ�-��6y��hA�"f�.�gF��b�*:��C��gi�u�����(%��7�3;Qҹ_V�+d²��o $����������*�&~u�k�
 �Tt��k��+�7�Lb:��Y�vB��;',��8 �"�y/!�#BI �tή:*ʒwV$mb{��6���xԍ�E�@0�k#L>�u�P���Egi�l��/���9��6d�T���y�S@le� 6����>d��x�Tw�T<�	dT.�3�.ǜ�y�o���v�3-�_D(��U3	M#|�)��ҚÁTFgC*���p��`y����#a��z��<#����	�x|��܏�c珅4��݉W��y\Ik���mc�2�̷�)L��n�>���RNk}y,��!��h��.��9d�2M�c�(���s�$��Ϝ�; 7S]��S�ZRz�zs3g��g���� ������?����q��C:��1_c��q��`W�ׄ�w�����4|+F���tCJ��ZJ���!�ˑ����抇&��H!V�v����#ۓc^u�J�Bqsnc�CU�c}�i,��3�D��y.�	�	����p���C)��nTKt0=`��Aձj73a7��b��sk�N6��C�B�!.������6�})��i�ϖ>�[�l�F`y����,2J�eP�����:$�26���wy�/�zG**��N��VVlh|ә4���ݥ�5o�=�7���טBr��L���Z�]�J��� u�5�if�zs���*��Y0�4���Q+�V�G�K�i��]��Α/qW4��@�eN�]�P�0b/� �[Mj�f�/r��w
H[�6 4����i�"�C_hw��up��n��+y�Ax�Ϛ���O�Ʒ�&	��j��s�#�J��<l��"�ڛ`�+jO�9m, ��G��Lzq�S�v��>.q�-�c�]?�g!8��{��Q�f��Š)el4��w/�z �0ܿ%�3�Z5���UkvF�i�.A��|�re�kl]-��{�e�rY���׭��%���d+9��>��
B95M�Lj���vf�����[�uӆ��T��\y{U7%��Χ�!ek�J�[�c��ИC���[Q�u�M�=��JJEȂ����'e-d���������Fw�(�����Y�UN�{g�s ��Z��H�33��h�֨-�b�Ka�mpj[Nsp�P{�V]ߘ�$�>�{>c-��0YzS=r���m��&pʖL��	��L�k���ހ'�����H-��׺��2z~��tּ4�蛖��7z��-�[]i�IqG�OtT�m9�6�E��z��C�D�|�#k��y-������5`��P�{�'+�d�-�y���`#᠁���O�aZ�V$�� �skL<i��@;���'�^��ƬgH���BΤv̒�ҜFA�Ȗ�$��=�Q�����L��+}����Ĵ~[6�-@���sgkjӽ3jW��_wbFb-@]�!�D������E.�٩ʶ���%E������]���������[�=b!���+�>6z����@����h��)���u���D�}���$tc4E��]aq����n{��9"i����3�5fU��4��_{���)���v�sƆ���KN �tt=��v��'�1&�e،��jE���biP�hOB^:줞vS��h���hS8�S�ln��<��Pbj�Dk��!��6��oY��������y~ec渋cçV�=x�AA�@�*B�7t?�{���<<����۫���P��xi�����Jd]��p�;h�*B/���5e��h>�j���"j!�3L��a��YB����ȱǸ�OI�.�}ڨ5%L��sނ��Y�I�r�>�X�5�"��R!k�L�T��:`�x�r��ݷɡ�C�]"��ţM�q�n�#��1JЄ���=��p�6 �:ǈ����6��3٬Ig.M@�0��[���-l�px�z:�T:��6��@nj�w8�����l�y	e��jDC������u��}2+�6��䯣��[�����Qg��~����z$y�����]��7��\��q�ь��ޗ��x$nq́�I.�':w��p'�ڀ'��"�ɫ�]��Yy��.$١'�>�y����z�@���18�P�`&�&�K�Ą�����"gv�1�OF������-�j�/wN��@�^���,wL`Ab�!�����dH��;ݶ�gwn���u�1�y&�6ʄ����Wj�m���Գ1��r�|�Ӗ.�9s��b�2���^G[��L��o]�޾�3x���k���n�bm|<00fh_WX���#��˯�Zk��>��?xB�����L4�m���7- �_�ކ�|�b͎�L{�_�2�x�xZ�����5T�Mo��v�9$z�p%߸zo��.��3�����2��
����)b��FҎfۗe�R�nM��{�<﯍��qs.![�gOB��r �/���kB�O&j��W�����]_�jB�~]S���N�3겤��Z6��xH;\��qL�t�b�Θ,H�x����6E9��6���:f#V^�P������扶��q��d\�%���c@<��:���qa����=�]��K�O�^�m����[����S�&_[a�m�wh�i(gMmY�9�I}W���
�/�z,��B}�&�i�g7z�x�%"���x���5�^�O)�$ȼ&/'mS��ֺ��̑w1�ٝ9��U�RIa�25�e��˫Y��p�".V�����0J�7};�`�E� ���ↅ���Q�b����^���M�w�`Ŧ��ֺ��~�x�H>�@Sߩ�������s>zP�"���q�� /l|���{5�n=���ղK�d	b�>�bo���m�2J���
��Rβ^R5�fojH����;/����`:�������^�y|�b^��p2nز&�e�ԇ��N.,ӽ���9��:�*<~އ���B� ���I���Z��ބ�8?�vB�5t4���Lw��D���ߢ�-��\�ОB. Z��ʟW�W[��%���RU����.#��^%V�V��C�&bN:;��@[w�T�+���߯e�&Wr�'�� }kn�f�K�2��X������{��~��+���H��&��'VkAK�.o.,��%X6���*z��	;/��a�G�b��&��k��~O_�`@��q79�ן���U��}�H����m�-�}�����'��g��nGY��"I�E�LT�qv�ڎ4�ca($��!LN�D�*�6A3n�9����Ξ�f��QEj�?_"���kD�|�������".���c��=���(oz�WR����D�r��c��qo䖖�2����gj���u��ag]ڶ{n8���ip��;� �nZ�]&�V���=K�+[3m@�1.��M����g�xϢ5%"�u�F)�j{���n�%_/Z�������f�<�*�<���c����=��0h�A��D|E��^���H��/ۈ�Z4%�-�o��+�7Sp`z��j���y�m��� 7ihq���^+X���t��pJcE�P�C�N[��m�����d��Lq�
�c��>N�����v{�P�pdo�e���q7%� �Q+|�l�{n���:8=t�"w��P�cH�ƚ@|�s�8��
�S�{�k�z�p��
���-x�pz��m���h�q�W������;/����Ӹ@h��w�-���V"��ʭ�e
�f!+�T�&Z���������K&|����}SLyL�����v�G?z����9��#y m뛑��*�=�8�N8����5Ꞙ�V��R"�Cڶ�Y��=[�*)�����n����j�J��K�Ǽ�b񇁮����kR�BR���?"4����F������8:ƶ�[�{eD+n7"��Z\�L7KR[t���y�{VvF����L�/v��(^K_1j3o` �[�q��^�<�|��rq���) ��`[�e`3���œ�ↈ=��00��H���&_�����&�	��@��
�R�������D1<��u�HCz��J��c[�*�ԥ�����W!��LF��U��ݲ+x��5q������~���<�N`�:XܯeI�7���}�=q�!@ZC
4���8zގ��KF_ݴ��cY�0�ٰ��M�qG:i�Eu�%�f��}R���0�<�Xb�М����D���gClWP�fn��+�<����۹z�����؂[\�b�.��u~�ut��\\�YB �b�{�ߪWQ(z��j���$@S˼2܁�z�\�rQ I����enӣ����+��mg6����M\+�h�F�����]��!���s�-^�`��<,�q�ȼF_8+�dLs�D��ٮ�ݝ2����;��paD@7N���N�`,s�1�,w��2����~�k�5��6;���M�r�*�ڍۂ�k	�S�;�%o,
M����ƴQ�h;���z�2�z#YP�fJ;��r/j�^XNl+��F�њ��R���ɜx��^�����o��M��M{K��i�$@��!��v�v�Kig�ɓ��K�G�7«��f�H��/}d�ތ�\|#�a8͔<�'���Z�$W�$ŤM4�+��mG/>�7�E;����{dt��;��,����q7���T.Y�O	�e�t�G�YG�����f:�B*=[�~�]��x��[x���v)�ݟ*ث룤ټ��ާ���#��9��{�浊�z���y�Im��jUi�����o�Wr��ljZ�g,�� ��e�v�>����o-�Ǫ ��8w�8p�� X �I�Oh�2����){�!�˭a�#���E��E����v�b�NA��D�Y�l���m��IO3�f�
�&N�u7e���kB2@x�ڡ�*E��Q����`� #�c��(���m-y��na��KdǓ�r���=h�Z����� ����4_�q�cS!43������{�渧93p�����(Ǆ�mC����7zf�c4��a�F��1�OnCǪg`��ݻ{�^�r�+&���a<S[d��%ln�ҋzw,ň��CD���5{ �)\�Z`h�l;V9H��k-�75�.�����Ct���j�(����G����jCb{ngowD���\�����v�)&gXU6%;Ι>�l�7v�EuW
X�WTj�*�����"����[gb6�(����m����H����G��L��HJo ��%�#�.�f�����U{��[�ω�"�d�!�ѫ�;{dqP�-f��aB���ц:�@P��uy��t+�V=��\�
�0�V���s� ��|�
:�|�,��]�ُ���VНc+-*<���C�W��vl�Ǔvv�V��#+M�(e)-f�wN�U9W�{v����]UJ#�����,�u��;��]����ϩ��C���5�nޙ�mdQE!;;2��7ƫK3B��t���}&1��
�s#B��bXbv%����գ"�6��E[N�;S;���7��j�1,0��a����z�U�d�ԇV��R���J7N��#�ιX7�e,��I�&�{�C̃��;��Z�ꪻ|�}J*�[��ˆ��.^Ӽ�ޒX��{������~og5����u�,P�m
Bb(�X �L_���,��` �B
�����"�Ѓ<�X�Dp"��njL.�Yƞ�W�]ݳu"�Jܪ�tW�$�c)��U�\�y}LUکr�Dw��9M�B��ng1l�uY�	��6�KN�M0���rȝa:�)fj��l��x(��k�^�._���osj55E�P,�mݕ�8qn������8)JmN5�*�Sۃj��g&�0ݰWd٧yfzr��U��=��^J7�j��h�b�7rvv)�!gUQ8f^j���6UX�WX�N�GY3H��[�d��vK[�1A�����ќ��%�8�Ur�,E���E:VC�R1	W���R�0Ct*�����r겄w��>}Y��w�6����q���8W+�hi�@����w����@A>��H���˛
7a,�9dn�.����5i��	����hkJ�b�(威�/vNب�)��i�]%�p�yѳr����s2Mل��K ^���s��)���#b�ags�}�g��l��ܣu7Mr�@�R��R",���bD��'T鍨�#��*,�n�J�jv�8��唁/#rM����욅�{P��XdoC��6�Uۣ�v嬼(4�&یz�b�FLA�)k�{�Z�;Έ���%�꭬�F,��e]� �zp�Tţ�����o-�خrMT=.�{;7���3	�La��{@ F H���4T��W����I����xשׁ��ʋ�^�4ԔfkȒ���"B%>:a�����~�4Q�9�9e����EA5PَE9fSv�a�p<=0Û�*�����G�Y��P�C3;��8��;��u��*�H�����4��x�i ʨ�2h�̲�*�f^��7':¨�<O��9]J�܄���u%$z�������ՅՔZ,R�$�H�O<<=4�<���!q�ITP�M͑MSLFf4�M9�ǫuE%4t4�����8�II$!�FAqSPVp�W�rd��R$�����~<<=0�w����D��%>�Zlp����E�d���ȉ ��"It������-*LDTM�*j���z�݌EQƱ�ubEU��5�YU0�J�dj5�M��K�(�*��+:���\u�~��k�j����˜�ԩ6�Y؝�Pg*!��$�`MVQ184�%��]�'`�W� �. @ �84s*�J��+0��Ể[y�2��3�����ϝ��'B9K*l	q�[��x�S��uKV�K���%L>�}���(f���]�=n��kۃ�HP˖W���q 33�_� wáƻ#��Q�s�Vs]�/�� Tصr*�6�{78O#lE|�wqD�>(I��q&5�����3�̊hVA呇dX�����<%���7��X��빹0�ۉd�h �2|�/W�A�x�K��H��{4u�Q�q�S��Y;X���B��p�@�U�n=�d8L_'�*�<�,K�tD����N�"h1��ƴ�/�|!��Z*�\��US���U�C�Re�Zmgqy�X����T#G�����un�4-�[����4$<"�:u��ҳ��M1�ʢ1�y�)�i'�A`����*
Ǒyn��}��'�}*����HgV�Q�[yW���\�>)8�����C��6R�U�ۗw2�[�ܲ�pv�Wr�H�B$}��'X]a���+)�+\��*��oIk-�Z�t��FrrC�,�Ɲm_>�bM6e>�ՉK˝�1��v�cR�.���/�|<�?�����d���ɟ:����k��%)8ZJ�e����]k��d��*�f�r�V�p��Q���[˷�U��m�Ȱ��&c�����/����Δ�3 솺�bn�%tW&�M\Xi���2󥻷���� ��r�V��=��/S"뉸۹OP;/H�=l�g�M��u������U~QH>��x3�x���Cy)�`�d��fAk��q�i	�=�j�Ү���'��"`w�7:Dihe�[��_w^I�\�bp+ٜ���m�@9��_޹&�0ɰAlԉ��7_ޓ�0b�`�߫����/�Mq��xo��ϵ1A�sb}lo�a��Ps\�	�Sb�="�2o~Dv�^����vR��=�hO;7#��T����`LM�5�{t�"\XK�gv���&]R�
ڎƼ�AUۦ��n��"�jV��F췒��fܺ9oaBiyjy�O'��U�b��E��5��p�x�.�1[�yX���K��u�V�iv=p�Yz���;O�Q�*�]:k*�U�c#|4_>jL�``� A�0h�F(��Yjgw�>��/�������V`"|���a�{ uQQY�2WO+7����|o�|��g���=�I������u\r�F2A��v\�x�l�[
1�v6��u�3uɺ[_K꩎0�Q`��~O���
^�]e�M�}�Hq����	�N�v�u4�P�����&�+��rVA���f'���]�qW��/v�����`.[W�v=�M�ɫ���a�~k��u���M��s|NX.�4#��	�1��0�I��=��@X�
�n�YB�����P7�h�!��h�`Myk�TtǄ����k�(����=�ΐd&�E�B���'2^m�/&��ߦh��8�m~�i���䟵רo��fg�v�)5����[d<e� %�p
Fg7�x=�'-w����{������[&*�՜��{�#�>�yR���Gk�ZӞڢy7�Z�A�Ueؽ��/ H� ��$`���T\�e��+6ӵ�1L8�iQ�K ��+U�k�[�����ck&�-��$���;[FNw�� @��.��5NQs<�H��T�x`,>c�y^��V!L�uh��� ۓ�Q��/A��ɺ�ӑ ��|}b7�/-�V�}^�6�@�ŖDlC��]��N�eN�Nhd0}�0Ëp��B{p�
f���k��X9i1�¬n�>��� 0��9��d�y ��M<T�D6�Wf��;��iD�{(գ���^ +�P:Ӹ�ۃ�˃kn�����ݹ�����Iף��=�N\tv�ta�t�-�S�� �I�<�Y�
��S:^e�끠+Gp-��y7[^#�Ss���*z�u��鷎N$&z�|"jG�������ۻ��_�r*3i�A]�uAw5VU��H��1�+~��ct�����yAd�SW�Wp�T^Cz@5��mn��>��K!G"�q�Rȱ��K�
����ڽ�B�.I�2���uEXR��.NY��q*�.^��FE��\=�/�w¯�.�[���zq�&�8�w��F�8�.Q�Y�����Ǉ)Ρp��E�bjv���
X��{���P�{��Ij��|�����\Ɩ��� �}F@����u�"a�G�(��(&�?��|K��hjJ�ˌ��p����v��mDL��Ԟ��y�qk���e�}kq2�]�F@�L=���]��G=-j�gM<�#�ˆ�l�{	��-�Tl_�����<��S���ݒ�߅����5���H"�{NN�fe�L!�|�pB�=�}VCF��^k��	��a:Do_i�����kC�������=��$0`�[��u��M/��]o	t�)��ے�^]�j�����(W�-�Λ��_M�X��������N�l����t��k��R.SRy���m����%^�쓄��Ow�0���h���o:H�[ԦE������]�6��M�z�Ox��7�0��,��A�W����,+�2���>��Z;�Pw�mi��G��d�&�D�4;|S'cs�U2�Ht`J+[NI� }D�M�e�gB+ȟ	p&����8y�s��i�sr�֧i�P�O\���0�����Nu0nj�ņ�аFh�����7c�yt+�EFv��N�[ͥ�5��zJc�����UT����3]����G:w�&�dʨ���r�*�]\���,,�+l�fV�`��<y�m�+�)�&�蚄{�敓"��4�24�p���*�3�^�5/��s ���S�6��,#�)ǫ��m7��7�����)�hc�*ﻤ�v�aݳs�Y V�W@���IRK����ӷa4��H]Y������A)���K�?F`�=� .:ď/+/��zy�.�"��7Ϸ�ݩ�0[[���^�+���r���`�	�Y�-��� 2�徆p���h�j5W��D8{����d-ѝӷsZ�N��*D�x�ܣ���\�@2�� 2]ӻ듶[�+$�M�kD��s'=�i��x���<g��	��q��fr��z�ܛk2V�]m�r&1�:I�Yq�7ՙ3h�l�E^@��zqn"���jZzq�t�PIh��8��9��`D��w�W���Y�cK�;�7��j������pd���v.ܝ�����;���v����v��h�A�@C`0 !x�$LҔ��)�|<!���,��s���w����,�8�H��'���d ��$u�0@H�M���^�zD��ճ�\�T���7���p
|V�_MŰ14#��h�:���Guَ�l��g�s�u5��f.Y�ՈҦ��'���
�YFly�툴���Gt	�ේG�[ d�!脦{�5��7r�MJ�r�-�He����4f�<�X�Nf�1���s�4�Ϛ�5.�g
~��4F�<@�*��js{�,�a��:����t%����>A��oS)ۢ折�3�u� �����%n]��[��w�f��l�h��-T�[ �5ԬV��pg��d�ڜ ~����H�����4�����%HY���R�{�;�iH�� pDM_F.��Q�Z�u�oi�cd 	�^��l�V�ٕ%����[&��x|���eT�z��%�G��;�Q{��<E�ͣ�D����s�2m�ԢǗP,"�ʪ�E�$,CX��.��u;R�!�;O��pv���V�s�A� q��n���b��KH�cw7]�)խ�d��JU;�� ?��3s�b�0>Nj>}�V�Y;�{.(®�����b�r�z
FAT_�=&�yt�=@<�8Ƕ�����m�j�  ^_*�Kܑ��J�\��o _Fn��QU�ٲWA��]=)�7+D�yS�E�[w���`�<�ÿ.�:�*��Kv�l�ȉ0_5��f5m�Q$O��.7�3�HhˈP��h� s��xn����sWT��F!�c�����q�0�"����ZS��T�A�g��d��g�:�����>=�z�AD@am��n�����/��x�,� G�ѧ���\��~�J<�Eh�����
�0s^hB�s�*����]̟��=Ɗ����>D��g3JQ�K�T��D���z@��D��x��]��k��k3[FU���JmL��7`��+Sx�iq���ל��	�5	�E}+�}Z��P����}LvdY�gڋᵿ��1:�5 �ςU3~��EHF�Kj�#Ui�{C�L��1�IyS\܊h��g]��t|J3"���)�V��V��19ch������gu#��;��ٴ��x Z~�w�ya�'�Q�仨��=S�-���UN�"DG���9q�I��Z�xޫ�-p\}a,���̨~W5t<�f+�3(S޽��i���H�-'3
]�4�M�(]���qdϜ=�{k������{[([��2��IdV��
���zc�?�ꐱ�>W���� (@���!��������uk(	�zZ jy������Wq3#z˦���=:���գ�_ ;� f������sg^`$��Z-��i��D�)���� !�@��N!�[�:��P��}
�\�
'4z�b���1{��)V��Ս@�����z��b� �z��N�҉Jw^[�*wh�譢l9�-�����TΛ�����pggl����#�;�-֛�0Z~߸��޾�*XL�@th�	�A��h>�qBv'���3(Ҳ���&��'pTF=j�5&r���z���n�7����k�U�1�{���f��`��X�l��kt�.e��EI�d9�a�ݼ�����6ﺯ�Vei�+�.�r ��wQ3�L�n��M�3z�y��7�<no�&
{���>�3m7�89��;X�_�`l���}5�u\z�V{����KJ��1d���½�!��Ó�p�4;��p�R׳b@�A��	�0N>��~��%O�_@n/NK�R��t��-8t�`�`����3���*3FHk�BV ����5�)��� �G5�ѥ���`qi���ߚ#�txR��^^�Js���OB�Zn���~ԍ�r�o��׶Z���Nr�]�ƛ�.%�ss!�sG��!���F
C�	�]�7�rx��|oR�1HƙM0�^n؃���S��2�=_��rv��))d\#\�v��9�n̉���%Gs#!�MP������{u�D$������WJ�:y�'��Ms�H����"pǫC�����r�pw�_����V�:��Ty;|��H*ŗ�[�X�,��*e�<:]L:�2�u��m�g�_�<|^傝���c#�U�Xh��������Ct1d�V�vᱫ�Yf&�k�L^��a�µ;z3+���n���TE��!�X�4(��K����;��w����!<��*ܑ/�ޗ��]C8&�ՙMRhP`�-�k'k�f�'I��늱��+ʆGS/5�Mk��5ujS���1�Ji5����VRD�A�SJ�Z�DB�
)��yYa�t�ː����]:�y�笋-�J�)okD�V�g��j(Z�3�2o�/[��qͭіҴ=H�}+��%H%W=�0ۦ��u8�,�j�JF���Mm���MYx6�4�ܽw"x�A��3C0��dC�Ř$ڶ�hܪ�au9��fD��P��V��4��h�lo1�]���U��0mm
��e*�N�^��]��6vOI�u�7Zˡ7�����+bհ˂��Yf����e����j	��z�Cٝ�wB�6�sn/l�����e�˝K;���5X*)Y�dl2�F��d
�i�"�SII�)	�������.=�lc6۳� �\;r�j��up��7B��Ö��E�s�໤8!W��&�ν�(()xА������>��uW
��J1"��WX2v���Q}P�B�!�+ Nb�jV7��A`���#2fB��, �,tTi���hX�cE!Y\1�$&�!(�,@��b�5��;Bh���(s��5��J���e^̧�	�qp��/P5�pˢE�oT:��i����s^�/��uWi�ͺ�[��Q=u�ԕd̢���`4��KAf�D�b��]e`��z�u;��	��Umug&F�N2U�f�[QY�=k^�آ��X2wD��IBѲ�Mc�.��1w.wѬ�.q��єqܝմ��3��kQ����tTз��iT�
eq�XNW�ѱ�=�:�&�)qܭ\���U�Qw{��X�嫧ǡ����{��=�G=�q#����Gk�s��%�UM�Y�YqЃ4�Uڃ0L�
q�Ņ;w�
��a��S�6Y��R_KS~}�[�vs\�M3v�9,llܱ��4<�����,�29�¡x7O#L�v����|�ui�XtS�y;^ocMt�A틌AU�]����f��������'V�r�d�M��
��0.ַ�&�y�Ҕ0f�d�e;�����t�.$�YZ��*�R�4��e�MALۼ��Xj�1Ų½�P�@��N�n ��a��G���t���Ī�#!ha����B*a��eK��o*-m<�I�Fն�7�������	!"��@�uh���ר�<u��t��:E������8���պ����N,�:G\G�un<b޸ `!B@X�шC.f�P*�X�@fG7j%l�i�4�Y�/з6Յ�$$���� PRD�6�ddy�EDELQ[0�"-���:A��9A�i�Y�Q%5111�(��*���QU��A��w��RI0�<<=>0��5��E�_!�LL��+3���5n�l�2�����<��:N�f쉦`Յ3��YD�j��N1U��h���۴�EK^�i�����l݆a�ũ��ʢ�0����0�na��#"j��2)�R���h�$�wWQO4���<Fȓ!ʪ*Kz�U�bo1���*��*���4a��a�bK��$��"��*��Enr$�%IIv�BDI�a�<9���٠����h�#wp�7���1c�<\k(����0$���O��$%WmW�M4�ᆇa�uS^�A�G9�TEQEUUS3IUI�%�QTEUSET�L�`c=�Q�-�Qu�[���h��!�&�9��ՋWCfա�4�Ǖ�Ԯ�|��r[]�+qY1�%�w:LT9��J�j�t�լ�ښ�|;-�a�5��
�(@C0ƍ0لNoZ�����|S)`��@��7+1��_�7� �X0;�g�`�����<�+�Gv =n*�r�6ExДOK����B�Y�&�dϙq����lן�ym��$ Y��,	���N��l��H�s����o)s^��>�dV��$���Ҡ(��S?��-��h������\��}$KP���{����^��5-����H����OP۾eg����>+A���E����B8	�m��ݢ�%�7]�W��}ݽuNP&rG{=p��I��a�,4���9����ǚ��Uک�d�ג::9�P�[��\hM�ϣM���E]k�D� ��c�i� ����� ��
Q$eca�H|5��(D3��Ҷ����00D������}ް+&1{9��HNߴW����v3g�)�W�a�e��ɿ{��۫�[����� ����$��B�(l(��p�tk�Y���W~�F��&����r!�Վ�ﻭ�����ð�]�U왗/_Vi�z����h!�B
�`!p���-	�n�G��n�]l��2�3����V�)��A��`��*ڔ`nKֹ���� ]Ν}$����ώ�T"տe��P�� 1�z��1%>��lf��g�sk~��{��A��!q�DhBF�ŵ=�!��d
�6i��v�c���;. Tދ�+bwmѡ�Q�:��|�}��}l�=�xyz�r�uz6}�Ĝ�5+�*��̩�X��+erA�j �]J���W2����ȧ�féb���;j�W���j���^�Q��#�8t��h�m��W&�W��hk�����cYr#�*^%�3B���#v����2`��s�΁�I��d(��Qޠ(^��.(�J�٥�����a�t�5#�|K[���k�]B���t�_yǹ�J��9�+�f����\q
��m��$�B9>��� rY��]`���սj�^x�W@��g�3�޾�ppq��������K��ۡ��9�]��UA}��U�3Y�V�ځmS�.��i��xf3���6oeZա�y���r0�T�6�tW��ָ�yt����x9r��f�:VZO�ԪCG*��������.%|
LV�<[���䝖�<�����g��`����  '�����q��J���h'ӌ>�:`�v� ��C��T�J��i���0.y��-��(ͬўՑ�k���l�c$���۲��Q��j������A��5� P�m�� zg�n�L��C5�i7&|i�S]u{E�88p,K�~fM�,�lU��
���S'���$��}Eo����#ϻsx��vxx3��$���x�H�n�ڜ�Jt:���� ��'���V�a��(N�T�Y�zb,��Y�:�'2AM������V��
�u-�<�|���0�I����q7��@[�t"�#���(+�SQ4�L�w#y������ݼ��=ZV�*@;�ʌ,��ԫ�'S��N^��Oo��US��)���ly�vHI빱%�7�h�A� ����k�FNX��� �Uح��G{�G%�R�l��^c��RX�JhUenÝ����}�{Us�믤W�r��D������u���ٲ�u͓�!;�R	۵7���ɶ��5:����,S���ٓQ�uu��4ӓ(�� �0\��Nҙ�����]ʟ͠���\���s�c�Kp2�����r%Qz�k���v�fu��AR��\�z!���_aܮ�����aS�S�^\�����o>���1��Ֆ��C�<�)�����w��/O �Uc5�����aX�/�3���-���Pg'��fvg��T��_T�����}8��{ �7�H<RY��ۑ|R��v����ov����_f� x��D� ��h@�T	��ԢvFR�!�l<�E�[c�c:+\H��_-of���2h���}��r^7�_Q�+���|]�Е"1���B+�i͎Tfp��ޤ������:z:�
�h��c���t�x��Z��ݝ[ ��{/Z�x�s�MoE�=N�/�Sz �yx�*�<����)|�=T�:'��݅Q:����5�oRw�ma�++���M�=��!>�D����p���z[�&A��"����&=����Uݶw�����mE�n*~�^Q�EGqgXŬ�]93J}���i�.�mf%�{������cŚ�qmun�--�D�!>jA���x��ڣRF^h�oﾻ` p��G	����� �rf��N47���q R�."�P�+J�;F]�jD�XV �G�����p�yR�' K.�]��ݝcs��R���p�]��г<tB�N�H��c��cT��"iA�-S���{���W �Y]׏<����XT"�N����n}��dGsN��#Oqh8�,�Q���wH��&l�.����l�m�Y��F�x+G��^�����������-|�D�-Ǎ�����i�KdUB^��n��.�ɷ��[�<wJ���!;A?F
���3V�N=�ܸ�v�`Z ͞��Ĭ�M���2��.�˺���gk�I�uFs����J��y�ڲ�ȍFnT �\@���um��8�Z%ڮ:������������1<D0��"�h��`�Tkil�����B��ܴ,�*ʱwGҊ;a�����b�(�ji�UM+mڹw�U>�M��=~��`ܡb�9k��[œ�p�͔�W(n�"(6�>�om;LKr�j��l�{�C�ښ���/B���B��� � �ù0�I@�wq�7����f<�̙�WH2��]�a�D6�Tv!B뉑n>�7���뇑�`�:4��"���j}��2_��:����1]5qD<HOv��w�W�n�/A%����Oy՞���/�f4�)�I�Y��^S7���2v���M�\�N*Z�)b��9�z_"Cۆ�w�+�Y2�L �vС����aM�K��}ʌnhv�Y�8�|n'W�P�ʇ��,{}���U}?>�*\�]ߦ�|�h�)���x5yw�/_z~UcLb�s��t7��P6��3��-���5:�`�IV�xZ%�X)WNrhv��jZ��Voқ�ȩ��͚����/I�^.R4��b�WVWM'�v�2r����l|2�+r���:����#���<��6��KVޔm���������.!��"�nW:��2Z���pU�fwT����m���WE���C�Ee�nsU^�=7y�S�hX��Aݫ���⮇p�Y:�)<��yy�|�Y���o��+D����Q�B��^Q�%ͥ1���x�C�������J��<�9���o{�[P��$�IX���R�=�W�z�^n��c��K��ߧ�#���`;��q+���[U��p�q��]P�3̱v����*ӨY����n�޴_1h�Rzbf�m8��_�Ѻ��7�P��`�v=�z@�a�����ڄă�.͋���1zL�\���o�;:�-+���A�Q}�����b:���ộ3KrGibfu��7\Q��Y�f�e\k����p�Ƙ�{+.�QDt�{$N��Lپ7q3����0��=h�J]�#��c�Ww����ᝐ���"A>�C'� X���R֞B�q�I��@ތ�ه���Q�W�+��4���̦��$OMD])C�(�v�[1܇^/8�����R1S�8���趹��2+'�׳�(|�LN���uN��T���eX�.4B�i���QB2�o"�.�T�%HUU	����lSN[�Q�ѱP��X# ��2��*��s9�}+Iw̫ǖ��D�VlMvӻ���d�s���I�2�͔�������C�����h�<���������)͂wJ��+ֲ ��p��������_�ڵ�1���^�����1��7K�K"����\1�o�cN`�=͵SYm7�P�"����?L���7��k 0!n�!�,����<en�q]\w^Vњ�W�ugE?x�ל�>�d/�d���(���'R��ٰ�]�Z�]��� o��u��e�s�����zM��v���q��b	��~>@!i��\���EV������Cz
�ww�1vm�����cc��*�z !��E�R8�ڴ����N7�˼9�3�US�I��ʮ�J�5�A�m��c���g~o���?s�X�k��#D�WV�-ئ���8`���6�
��ls����!B+�(g�s��l��C57&�O�+2.�=k@�?f�x��V�~��H5�-����&۴�x�m@{�ú�;3G]	�I���z�CK|=+ϞuX7.:`��Q��83��z �b	o;����}f��t,�curv�٭=�3���ܒ�%e��f2I�ESk]?���{lo%��5��Dj8�]t0PRA��&�|��U�����[��h��0ŏ�j%����9�;�A�*��X6~�P��P�m�+<5��u��$n$'�湮DV���H3H�nΆ�	����o��� 	�/:�4�6a{A���wl���n]GP[�l�v�7���F���gg��Vm.P�;X�J���Xzi��g�`�>��ZJX�Æ��c6-֫��4ZvgΦ�����TǨ���j������l�{m�uy&!��M�F�~{�s��{�ݲ�f�/Z����y�զ2}�J4 sV��T1C�6�eWM���2<��%��C���� � �$y{@���
�(�s ӑe�6��o$7�ahr��V��|���?
�`1Z�(�z��o�͏���k�=��o����9��{��|�c�7�f������d�J^��Ɩ����	��������S�����	�0-
�?�VZ"���˪�c̔]R���m:�I6H֋�pS6u[�B��*5^=���Cv��HڿT�vL�dH���
@CX�W֯�V"�����F�=3M�����^d=M�|%��+v�%88`��]����.}l�Y*������	���ݰq��ykj*/vE��j#��z���QyA�v�ջm�ð��z �o{�<�����	�Ί�]^��5d�H�Triݝ���  �Tv07� P�1E�eܨ|9���a����]�(~ˣǪ�BN�2\��e����@W�I'��yw�@��wy	��ыN�ڥr��o��&�,#{ 7��Z�d]]o(b����.�����hUcNoQ`j9�Ra�d�2 nuu�k����7�y"�� ���cN���fE�N��bHM�����������6�NmyZ���FoM0�c�l��� VM&��,�"A�y�&���Ĵ��FḎ��K�Z��+i��.�o�����};n����=|9ʫδ������|Ϸ�����:be���|�,{j��m�,ۭU/�k�w�W^䭁G '�W�Qwr0Nfs
]���yk�۴طV�)��'[wsV��a�7z�e+�aUt�T�/Fb���oZik�^�:P
����y- ��٩�Lv�[���m��{E�ۉٳ�J ݮ7�}7/5 ���M�9a�-�+��X8��oNr[]s�����(ە�\��;:%}�ɒ�X��:ц�R8oAt4�%S�&�j�T)T2�*͆h���u��
��{��C��^F:^_���/#a����� �Ӹ�����\ŻY�k�Zgl���#��5zޫ^�C:�:mj�{��f�6n7��Nj6D?��$��5�:M����_di���)k�ۻv����s�%P���f㔋e\���SW���1e������)�8.Mt�ڶ���$����[x��i���iF����X���ocv%M��y5��:��ީ0�X�*"o>n�'Tͷr��p�u՚�z�}�BɦW����숴����m�E�����ֳ�	�J��:m�e㸲7��9Y�Ww#Ʃe���'�Ig;^���d�H-�G��a���"�tr"��![3�O0��3B���^�.�R�hZ̬�Lc����QNMӸ�5*���-ⷵ݀������ �G^z�����q��uָ�^#�:��*$uq��:�|x���k_��>J��z��;i��z[�<u�^�m�7-L��ic�	
���l�o^��<_�x�g^��{��qc0����#�����Ǽy�Ƀ�iY+bX8�`�k^���f+$��l���q�S��[Ī�J
���c���޳��f-r.q�{
4+���CY[�2�GV5�u&�^D����g,�M��W�"p��qZ4�^Z�k#��b{s�ji���o\����V�&�����j�Z��S�VmG��#����y]K��x�y�B%��V�M2oܛ�9//"�%��J�a˹����Uc�	n��!�x�m�w�+�*܆~�$V�X�o5'�����+=&�]�����Y�ޥ�/u���
f��W����[�ڛ�Lv�wnLt�fqwLn�)+�Ws3}/�-�ݗ�|�w�)h�l=�N���.�QU|t�܈◻����d�H�b����>��]F�\�[�j�E%�"��:��.r`�x����	(�ٷb�·�f�\�9W9��nni)�X�
iTc�͓hL2�]RTQ��ː��Z�l§f�Z�Z/U���4���d�ښ��Ez:����Xa>��YX0��w��i�R�Ӟ
��C[5���	g�����X�]_V\��br���n����Vb!���<u�k����1��Ϸ��R	R\DT�EՌ��LASL4E��E�����E$�$�+��.Nt���ٸ���*"��("*�C�2h�%�*b
�����������i�M:xzi�:�oh�����"�H���6c�j�k
��h��D��*���M4����L/{�g*�"&�j�Y���%S2LD9;�y�k
n1ɒI"EI$�4�ӧ���p6EW9��DE&�""����0ʨb���0಍�]0�ç��r�I""I$֋	(�"*�����)�I$I�a����f�"���"h�}f0����d���,�&�I��rH�&�i�����s����I4M!E%y�R��a�ݔ�)%$d��R$SN�4����<���$�*j)���i��������"������c5T�AA@D�R�U�ȉJ�**��|I���ןeu��j��[��B{�1��ݕw3���kY�6ܡ�=�գ�*TfX��и7��1�@}���=�v���g���{'/k���*�o4�k�y�m󾏩n����������r��$���-��U����fL���f!�M�����Ϩ��=�'C��.0�;��ǅ��F�N[�جd�Y�u���7�� �Z���u��=���u��nk�h���_qfot�3c<��߹?2u7-��oRx�E�%�Hᇩ���]�/R=��nA��G.��O�(g;�Xj¶�� ��Z�ѐ��\�Z��r��z��y�w����@ȿ��$6�f�F���v��k�N��/5]�s�G־��O�>`d[��m�	�>��2p�FS�S�mU]�Ұ1��X<����]&_et����<`��ށ��oc��q�O֛[�=wh�\ ��{;~W��*��&fUI%g�a��+��MHw
9A^���A��wv^�dU����wM7a
�x�;�ٙA��9��O���o,�f��&�����b�$#�{���;r��4�m�u����g���ɇ�����7��؜֕�n?��|����R,`˶�ޠ-0K����]�U�1��`:����}����L����5tE`7��f[aE�}�߫��ܳ��� �=͠ǐ~m�1�RcP�9���H��_P���k���:���g�����n�ri�'��d�޹�U j�����Q�Bn[!`��2�D�H�u7M��a{��&|�U98{0���Y�� V�(��"��f<��7,�Q�WG�:���4�l��^�oz~*)-�2g�Ԭ�)尕?	��b��@`5�܊��y�T���=^,V���5�7�Snf���>���ɘ(FD���; ��jqK��.������ξj0�[Rة���f��x�zYD]{�>�p$���u��g֬�fW���/ q�#���s��^�(�1~.��)K$�d�n$��1z��4�IR�)�li�[�Y��	�"u��ݷ�YiSTn�,�j՘!�������z��V'�릊_�3'��~( ��%u�,EfA�����7yna�f;ЯB�L�G_l}�}=�ٳ�Bi5laf�����rq=����E
c�c(A�����t�f	��p!e� ޹�^~��hPC|[H�Cy�7~��-Da�"�S�ue�pJI�pG��7��F��y�n��u��*gy�������.��P8�z��1`�i^�G+����� �@��X~?"�%2`/ l&q�/^A����7�7%�������O��y>�8Vr�Z��d�cz�9�`ԁ����{�'++X�7Hh�v�ف3*�xo`���ib�Y,6�Z޷g�-���Ua�7���ߢt�a_H��[^7^��d�ڹ&f}�&z�u�^?���"w���+�	�h���;y���vX�R�u[�MWgiv��
bg����3��w�� ��Ɲ�o�@�<�ý׾����gļ�s2�
��r�Y����#`� �o�l�7ܹ��z�neD1�g�Q�o�� F�`�O������,�&!�ǎ噺�&����K1,�܁�6�r�II�x������y�f��w-a���k�<�t1�l����|�@!�ʻHZ"��W�V<�8cR��tm�-����r���5�]jS�M��Y���޼�x�^B�ms���f�q��7�"���b�>��~5��JP�cO�xa��z	T��@�:��\�%V��`58}�$�G�}�;�B��6\�w�:��د3*CK{�d{moy -t�����ⅸ����T��u��j��7��uD?�s��"�X:���r X�F�������;�I�r{�JβߢM�i��1C���;Әޖ�F J͚��wJ��;e���9�I���,�Kv2�w)p�;�3�]^��)�&���v���0�/j����|܆��d���f�C��z{Y�*� 0�ģsz�߾�� :u4C6�?���@�?D�6��|M 2�����Z�+[��o�mM�qzP3��0y�9�h��2c�aZ��7h�<+�WϞƒ�|�B�>}WNf���h_p�}�D�pg�]�C��o&��B�O��<�ؒÚ�8Z�F�V�r��s�
r�8K�U��]˗���%j��%&�ڱI�[;/g�=��2�u!�<�> ����*�����V}��K-u۪�	��!��E���s8�|�fӳ�%�ٮ���̧���48�w:��|!9�V�s��&��S�p�o��`�w�F Fduఋ�e�k��+�j ��T�6+�̼�BQ�5@��0��a�ԍ{k�b�o�G?��-���P��1��U� ���L�Y��"3�T�Jaa��:����(Jl�����m��>{h������x�#��u���FVw�am�9h�b	:D�}�Ov����x>�6��ǡ��S���7^TЦ�ĥd����cU�Y��%�(�Շ_��c�+v���]�ȟ:^�kX�l[��������:�,�<��I������h���˜�f���}y>�|��6����]��C5@	�͡�W���i����b�wx�;r�l6MϚ@�	ֺ��\���Y�y�m�-�M���r�W-:I��9��ЭF_c`�a!���k���S��,&�xT��?G��/V�W��`ռ�ȷ�-ٰޮ��ukTpM7j�sxJ��I�%$rP7oN]���3��`p'�]���^�����,����Y�[�ŞJ�陷:~(n�7�ܘs
�򪖧�-U�]|ܪ����x~>�ׇ�9슿�H[��wn�~#�'��ሰ�0��r�p�'��z�7��,���TY*�`�}�1��������i�t�@��JY������`|��o�ݠ�@��[����E�_����Ƣ�6n��1��8�mLm\�5
�o*��s����'�CD��s5�%1��Ts5����B�_K߼�$Vk�$-�#�y��[�g{����x����ߌ\��#��Z��i�Nؚ^�|�p�iLc������dd��-�?hhE��YK�f�^�LF��uoZ�y>�Q��Vw"G��W��3N�P�>���I�O'�� �%w,Մ�T��M�US��:�R+���ޘ|[��篕
\_�`�ʹ�A�}��nM��U,���.�j��]��:m9;X���omlUU�3���z�a[L�s�g,Gvlf���]�[|��j�N�h`��Uk$���#��j��k�Fb�7B ���U��:z�Y���qZ�����>S���l!�ò�;�S�lj�7e��pqs�lF����j��+�른 0�h"B@�� D��\d%*I�(����nϾ��(!`�00 ��C8B��vc��9S���\_[���� J�z>�7g��C+����-��5b�Y>� ]�=[����J���	�4�10Ű���<~���;��yj����z(PX�ʔ��#R�1��6�˺�rO�����K��>��d��,z�7�^�힠��sk�,��!�w�R�U���`%�{,j�I��� �g�e�;�ǲ[�3!�Q��&�(Dw<������*}DLi oD��(8��˭���ۈ>�e�4 ��^�CV9��C�u���e�bP��������$�t"�x3��g%�u@O���t�;�|�f���	Y]���#�zf�k-���"�%A���u���Ps��C�
�^�U��̙��y��/�ٰ#�L1^y���s��bwf/F|�mJ�ߒ��g�or�åsZŪF����\�h-����Ӂ���wJ� =�!�*�{#��}ݧ�����׿�\4��b���3A?f�I{��N�JAѭ옹�{ݱP����k	A'�m��[�Nl��T�T�̍�{DV�f��EjdW������q?m��U3�0��ht��	� ?y g�����qg�0`2hFg)͵�ԑ���f�·�z�{�a�آ&��dID�q՚^y}q�ߪ��f=SKTե0��2:�.i筬p���O	�u�́{Z��#�8tu�� �oq�xF+;���5��������{����=מ)��P� ,�q�)�_r���/��Uor���*��Z�@�ڠR��*�!ukϸ��T?�΁�2�q:g�h�3�ˇ��^�C�ijŎQ�������dsi�F�մ�r��`X����4y�X8f[��<�� �U�#?1
U�b�X��ݎ� ����������
��{���4n�_m�h�(?�>�� �í.�(پ�'�Z-��܍�6EAE�uw�..�<��e!Z�klY�M�QO1�3�YU��7�MA�ٔqF⢾�,���э���1epaop���&���T1����G���ĹZz��WPL�tWPٝqX���ᇷ;6R�nm�3ﶚn�F���{��R� n�;�WKC{Q��	��(V�`�� �H%�q��_- �έ������ἴ�=�i���D}���Ί��f���e�&� ��NlOXCz��˨��Oܹ��q��>�!r�g=F�X���7�~�Ӡ=G���bpƸ܎D �9���Pf���ܜ��9�
���F+�p��I�n��9ٌ�>���R�9ㆵb�ðW����m8+޹�ߣ]Myƴ�œ���3��������/�@����[�U-�9n��K=�O ��`)���W�-���[�R/�
�6�>�FZ��37k�R��06~�ڲ�ܥVVO��� �}}��3m^L��l��ou�~�������@�^��9=@Z'@G��ʿw,�Cɯ���U�~R�Yt��A��B��wL�ٱ���Hz��":��[\$�*���}�K��wۅ���[숀#��I0i�,�7��ة�����ܰ�7l�wTZ�rq�]m9f��S;��fd�D�s9u���q/y��>��^�ޘ<\���v�	oHu����=���[�C�+��ޥڂܹ'3l�zΓ�i�un �R��.�����y��ՍEZ���i]1�u��B���o��(܃����������n2).��w1J�� ��[���ȃ�D�؀�XTS���Æ�����ܩ9��O�}kY���Z�~��~�݋[z�,0�_�>Ѐ>�/�[�U�.@<�[��r�g�y� ���ɦx���1�*}n�Ǔ=.ЇqT�/��U�m��o�:c��»ێ5a�[�^vz`������ٜV�ӈFp!�H�c�uСެ��NmL����`UėAp�<	[�����kM���"4�|�E�H���A�n�̀�t}(�y� {���Mp�BB��yY������� �"*������?��������(U���Lt��)�Ĝ���!�,��EUUr�e)D�)UASEH�W AR $ERUD�@E
9�G@�R�@@Q)U�J��(��� "�B
�)J�� "�(@JR�	UR�)BC�J�(@J����C��
�	B���RB�)B��QB	
HB� %*��@�U�(@@�H%UP@ER�
�	B�%
�@�E|����h	A�	D�h	T�"@` `J@`U 
 �b b) P4) � �@�)��B@�@�PUK� ━ J)��H�� �E���(��(A�h$��IA����	� 9 J@Jh P_���Nz����DD�@TH%Q�O��g�������?WП,�O�����_���-~��������ӯ����_M��?�?�������G٬�������������~iU����:~���  (���"" �
��������	�0|��?�_�ۀڟ�U�__�O��?��N�>����<�O�{?��|�豯�$R"�`!$�D*L�� �HȌ�	(��(�H����"@H$
�B0��"0�#,������K
�)0�I0H�Ȥ��� �@$ ̂�H% 2�$�# �H�(̋! �³ �,�0$�
�H� �ȱ�����#+�"��3
� �H0�,�H�B4�$(�"ă2-�B��- �
ċB�J-
4 ���(%�
4���ШL�H4�� Ĉ� ċ��*4J,���#@��B�"ċJ	B4(ăJ�"4#B�"Ѝ(% -*�@�H�"� � ҨR 4��(	J�B4*�H��H�P@0�(@)T�PX��H��H�H "UH�%�$R�J`�H�TJA)� �	�A�I�@f@`�$ �@�IadR��P��I����_@��)EHR@*�T�
�����~K�M����4�����N�'��?q�?�"*��q�����~�8ϱ�������z��= ���O�O�����>��UEz�������j}d�Z}���M�d��>jk��*��$����v����4�v?����\7��hM��TV�?J����~�TW�NƄ��{�����Mt�4��zH������pDU��o���EQ_��%�r�%/ԇ֟�����'ZO�>���.��ﴇ���TW���
`�>�ϴt/l?̜��rw��>!�{_'�!�x~�9	6��E�_���a�?jb�`�_����1AY&SY+>@ ��ـ`P��3'� bC;�l<��*A�RP�%JQT%UIJ%J��%H��ERJ�P-����U"�@�H��RT�P�*
����JH�JUH��P}��Mj��)"��%kR�hh�%J�T����A$%D��T��(4U)*��U)"�픑�h�! ��$�
��"�@��R�����D��D�"���T�HUR"�*P*�RUEE �T���"�UQ(��  �.;,�Н���¤�5��T3k����U0aWg]��j,�S]U��s��R�+�SR�ۮ��v�r�e�ʭ�w1v��mn�n�[�Z���J��j���th��|   �>��
��lt-��G�T�$H�ɭbF��
6�E�����4�'W6Yv۷N���mfڷl�Z�;u6�Ekn�pwt�vn��miv�wSw������JX�ih4J� ��H�  g�yR:d��ʕmˮ�JM�*F����K�n�N[�u��m���f�l뻮�nv����ݴk�F�Ԯ�E.Q��R�jmt
�'o�T�EH�(��R�]>  ��}m8�R�N��`J��M��j�n�ʪU]�tbV�J5�w:6�H�u��eV�è:�@�T(�$*P!I
Ex  J�h̑UI���`v�h����5m��V�F�M�j�дE]3[�7A��c`�΍4�#���:��Е�"���%%O  �'mV���l��çG:t+af��T�h�ڬ��v�4wJ�ՍJ�iG�X�  �)���UDQI	Q:��  �  �Z� ��
4�X  +f� &��� ��� �Rа�4��(��` �T((�R�E(T�o  7�  Ơ ` �i6��(@T5�  6��i�;�  �4 �iL V�#, JM	$Q�	�  74��8��B�)` �+  4F�( -;�@ :�����5m���L����  ,�!Uv��QDbAG�  ( �pp  ��` Hɀ� 6u� :4#  �c��l \� ��X Mc,R�� �~Bc*��� "�ф��"b B*�枠�   �~%)P�  ��OFU)P  eH�M��@ ��ǇH��������be�����{#]�鳰ќ�=(j��_UU}�}_}�%��P�w� ��61��q��m�� �?� lcl� m�s���ɦY(��R�Ym]�$��>��J�yS`W�.�á�@f���M-
h9�	ݍ���4e�1�[E:��-5zBzS��
����$'Zi�4j��.ЩL��9�ꩶ���Zz܌8�:TJwe��Ye�E曺�WqD` X�1����/j§��T&:ڕ�"t��CV��We��v���h�ނeY�-�(�Xm��(S�k-�K*��dɋ/f�=�ݹOUj�Q�P&�f�n���7 xnl�r�Kt�n;��-����b�!�a8�vH���^�N�V�@�� �v�����j-��%^��U�8�KN(f���W�6�i��?3�:�7�Gh/]��Q0��D�[�K���Qh�X�+5�:J�^�틤�V,�H��Ǜ�ߓ��%��Fa��H}�����\d$�0���"�4��Iۻ���`��!Zf����*�U�d�)�m�ۇR ,wB�2��̥R��و*ȣ��m��%jc���^��۲��G��S�(�b��okV�@��3N��%K�7\�l��)�R��2�v���� Ur��淯e���D�o�bk����n�а��8f�Vf�0��ݩZӃ4P�5�p�&��b���XL�޵v�����9�J]����� �$��ͭsd;Q�Ӳ��1-ͤ6���yNLa4�0��l@�W�Z��t[7wQ��(n�rJ�/0�X�^�w�*B�`��F�&��жQчf��: 4�ؕ��m02�:�ɻ�	��rEn��d����า�|Lx��f�۸^��R;#�.�yn�dV��SwD�;ېb[�^Eh�C#�1dq���L�W�.��Ľ;�U��K]��,����{n�
ʋ[�ܵ�����6�Jgu�%xX����ScB�ڱ��Ul�[�^�*H�F�Ѫz�Sf!7q�P�A�z���]�ot=�Ŋ��S/�P����Z�5�CE+ɫhfH	wJ�D�)Ul�I{h�n�Gb�*R3Y���S� �Fl���W�5��v}��Ѯ��J�8�EՏ��nTmf���̐Q��@�t{��wA���*�BЕ.źT��{�x��"#�{Ct�@����SnFI���Qgv�tד�Ė�ֆTƃ��
0}��%B+�T���6�Cw.��CG��q�����
��-���J�of�n�(�Y���K�I�$�� ����V"T���V�@5��d��3�kq����[[L(中<�%��Xvn]���amZ�P�0IWF�-T�m���nl'T���0-z�)�]��l;ڲUv�
ȃ�ח�6س�b� ��q�����I���ּ':&�/V�M�k!�H�IY��;4	��mөF�3u$��+2SH(�.��ilJ���¿��.�]�'+UnI9R髨����t���h5���%���%a%�c[©��9�hXj��B���l�Zem]B�ml�T�n��Z5�)���J��`�Dmє��їm�� or���Q��yZ���m�HTr�6n�2��l#(9v���ZC5J�.�4�X��hnhzsM�.�2�F����GV�5yuy�[:��[�6����vˉ^ay�vؚ��6�YHGCF�4^�;[���4e9R��e�4Su���qXu�Lى���8����Xա1cVIcU�K$�4��M�X�^]����SΦ����ԩѲ�[��[��[g2Z��0���u���	��4�ϰ�Y���#�"V&ޡ{�ҚV=Z�ͬ݊F�\>Y��e]⧺��@����3/x��ݳ��S*qJ��I;�)Q��x�1��:v�Tӯ.��x&���R �
�:5�W*�2�#	ƪ���g�n
��φ*ݚ���b�:�^�.a8&�LrCf�V凑����KE���J[J���vڋe�t��6�"8�&�^��VaW���iX�G6��D��)���0���]	m��O�ͫ�LXb<5)�HL��plqfU�r�nx���(�bͪJ��u.�8��k72�3iGJloA�gbg
[Z�E
���n�;!�m꿲��b��1X��Z^�Cv=�%;y[x��ާ/r:p�5H�ڲ.�ƹ�ٲ�	u����Qh;����\q���Y1 $Ю��,݅c�w�V�e�6�-�@���4�ʳq��C�5��=��TM�`���%�a�X��tm
�]bueU���Zh����j��{vˋ2�(Vk���Y��J)iT�"h�m�{6ӶM���t�Сv���V���o ��/X�*���Ty����,Z��H0ҶES��T�����ɗ���NaKih��A�MD��,��hŽ��,��{�L���i��X&ٴ��!0n�<�AV(��:A(�wM�djR۹@nJn�j�V�e�7��%�V��m+� ]�CEh9��Dg�:�oZ�A�L^����U�����2/5n�n�K�F�ܗ��vЈ�� L�͏q\vU��:5�����l$��oǪ���{��Y,ST��h�&%A�MD�£��,��C��m��e9LJ�.S���ڐe�צ��Za\����U��5R��tN<�J�%�@2;�A!.(�FM^=W����x���]-x�)�Z��(�*,����V�9��@CujĔKV�3�F�X���̏nc�
e(]=������Ѩ���БV�L�B�եK��]3ZaTfۤ�ǘv�(�I��E�.1��V���.��ۢM�]c�d6<d���R�)�V �x+S{db�)�7W�嗺���6ḙ��QNc�v�KZ6��8��Z���xQw[�Xc�/v��Mcz���LL��	�8~�����!���Tq��M���QM�4Y�O)ۭ��]Z�n�޳���ǺV;�+8�������ha{��FZ����V�鰪Pem�%�t�F�����-be)(嬽3)�(�J=�hj��v�Vʂ쵿�;ϐ�B�P�Baj+&���t�q���ud`��ˍ�E���q�m�R�oFˣ�*��EJǰ��c��^1wz�����iS�0;�f+��H"n�I��2��lرsjM1�c
��
 �j�*[YZ�XEF��1`^Q��Q�SoZ�(�P�;yY[�&���2�ˉ�^�d�ҽݦ��yt�ͼ4�N^�[���τ)-F���f��BK�,���1�f�yW
ۆ����mjB�𚛥2�֬�dm�u�\�eGj1Z��g]�� <�d
z�ʐvHj46"6���y�.ɫ�L�J�H�e����cy�����$	�tj�7���9	-۷�U쩢]�1d�Vm��D�T��@���r+�D�eݔ�S��ܭ�f5��v�w&#�^6��[B� ���Em`+UAn������KT�O�f�
�x�Q!6�S�Kd"�t2捘�ݢ��ՌRж�pMӕ���k�DB�ڒ��ǡ6%\	�+2�wwoj8�8�l;�H�DW1��*eV�&���Iْ|���ۺ�]m�,�Ӎ�Sp��wZ���]�Z�:
�����A'��a%f%�3Z�Ͳ4]�hۻ-�d�*X�J(��d����4*�ʽbe��ժLY� e��27T,��m8��V�؝��XZ�˴.�V�/8��*l�L�6�S,J��,�J-ӧ��f��+�v1ӌ�A#2�e䏄ċ��[�͊�'d��!�;+*��j��i�{����lS4;���CX��&M��L�Klc�K(�n��]�8ԫ!t���d�)Mл�B�5��#����5Va��Q^��:���Z�h;N�%��	�Y�)�Jsec��̡aU��6~ץ��b��l��b��4]���U��6�S��Zw�XvF�"�i�Ga�k�H�T'YyZX�SZ�܄��-)₵={!�l��2��h�����E�F*�#%JN�e��4챥V�YE �u*'5 �I��7^���h\T���{�J����6�^Y
[1QcRb:L�ۆ��8/�2^ ��I������r�q�� �6�QU��/�1İE
��еܫY�����J�d�j�R�"5��� ͸t,��#�+�Cʖ���(Do�8��Y��ǉ��]�0ټ�x �riR-;�����V��v��تYp1��t񷊢0\��튅�
���x�fH�T�CH�VfS_EL�y]ld�f^�񳂴 ���qK�[
�ڰ�]L��L��:����J�m�Ӥ3Vn66ҧ-غ���D蠴�
]�Ӹj�3"Y�Gt��&`�)L��L�PcAU�z�Y�̲���@T4=	�wA����n��Ɩ,�v�P{�����lŴeٖݶV]��$�Lx.8�є^�^��t�+J�v�:F��h�X7�>�F�埙�`Ք�r�n������Ц��N4�+kVbP�yJo6��{0�T�n��5	��+Cģ�'
eݖq:��z6Ɲ��ښ��Ue�N;�L]�W�b��Q�����&4,vn�i�63�.�m��D��x� ��e6��Wq](C�V�C2 >�͊eL1�J�1V���pV�5����+uV��{��B1X���R�MXaVM�Q�u�-�d�,Ն�i�N�n�3J8[��s��j֛1�g5EB�S��:M�bi� B�f�,��Q�八*(*����8u=ʷ;و�fd��V*u��FVJ7�p�J�V����CAc]��T�@Uk�a �鲰g�3�a�ԍ�7�(7Fb�Z��B{M���EG�is��i�*MS"52)�L�!V�y��tZ�5
R�d,= Ԩ%˻���wMR{,�����c{Y���ܨ���9u�E�
܅D@�(&r��$\Ez*8N�����Ycc��WYL�����դ���f�H�,yYr�ZӣKi,�M�r��Y�s��V
W`���kP�r�l�j(ˬ��X�
��Z�Ie��������@~�\�T�ر�L�9�#��ј-�	ë]t�DAQ��Y�v�#E,Ǹ�v�t����!T�-LQf�O�Yq۸�-�����t�Z��Ԩ��ź����K���ע)v�
�����Օ�s0e�T��Q͐�KF���f�hj�Ɍ�n
���M F:�p���쫹qS/t#��b��k�JtC�;���,i��#�y��/�V�i8������
�-[U{`V�L2]Zݦ#1�yZ(ȣ��0܎�U�`E�YM�,!�s
�+H+)�Y�`dfb�'�:GtY_$5�5�FꩻF��`J;���^�.3�֬ͬQ36��4kN4PVoQT�-��R�nڛ���yDQKONM����v@�e���Ҭ�܇&�p$�J�p��W�ݶ�[E[�[�s�ܺxϝ]f�����Hp�b��PQ'^=iZ��*�u+����	l�`����Gr:4&�Ф�q����+71�v�c��6�A�����s�r�ж�,�"R��ͬ-k���Cd�$�#eh2��6-#>A�mh�oK�j��6(�b 0�j���Fki���r�\�ݩ��{I��I`�w��Q�%�B�Liw+)h5���f9��!R��<���Ō�����M��S�A�a�%M7���u�ZVRG>:�ی�ũ��7X�^6��T��^Kn!s#JJ���:�ˬ��É<fSdl��e�[��Í�q��
ݦ7a6T�DTj%Q��B������R�Ij��6�ŌTq��t��&�UȬ�Ӧd`���#Z2��˧N�{���S);Ch�(�]���p����IQx���
���HBu���6#��n^�Vt*Y*"���,^\�$��w�EW�Q�
��Z�ū�)�.����ӒA�l�cm�j�fiݥ��]d��+ۦ�kt�l���	&&���4+B�m�f���n�%���ڒ�]f�F�6�V,˵q�'V�gIH���{�ʱ��k��, ��W1�	�Ͳ����ƒJ��U�����l���,J��a�bҎ��Hi��	�Z2'����V#��b�iP�I���m�a(F囸�N(��[f�4�������Ehv�xۭ9L'A�kd�����~�^*�L#m=ֶ2�5Z����n�d�m�6��e�t��c�0��f���vZ��r�Z��{�����C���OR{��xjR��V%e�v��	�Ǫ�A��Q�2=b��)��d]�d���S6^
�6�-HeL�+{L�۹Z�԰�)�ոS�T0�ղ��f��Zb�5�U7e��2��)��R��wSDТ�V���c8]m�71�,i�Gkbi�����	�_̍A0�\�or]�`���0�Z�R[����n����JՊ�ˤV-ݚRj���%+آ�p�kX�6�� �<�ëͽ�:
�6T`����d�.�Mڽ9*�*Tԥ��^��	��,����Y�#(��	�4�Ŕ�a� �=4�oenv��{X�^�� �r� �0���2�t=f�Ġ�m���U��!��+>T1�ʄ��J��I��F;C	�H�	� ��܊ݕJ5��U��Z���%f��1�0<��6�$���t���ҥ���U�M�l��Zf!��������@�[Mb��TuV��]`�vڏl��K���{�-p$���wZɽ�!��n�ҳNQܺ� OR`�L���2���r�`;h��0���8��M��oM�oF�`|�r�W�!��F��-����-"�!s�`�Q�W�XR�8�Sx�jj�P���{�$pncN�����E1[�n�[��KTMd�-�`V�Y�WU���Vև�4He]�Մ��ZLfd[��Z�]�a�ø��fք��s&n��[�ٝ��:�bN��x<ݚ��n�#��\4�9n��^t6��i
ˮ�۠���#��2>\��۹�{��1�zs���K����(u9�h.e��K��/��#|h��s��j+0��Y����pih�/�VFmcC���ۮ]W�N^��#ך�r�.B�EH�0���Bw��wT���+�o�˵�B���ň�+K3�5\���
�hu]��{��L�n(��z�j�N����5ZkЕn=K���4�����ݱ�gA��X��E����a�;<�(,���J_cC��}ۻ�*%��C]Z:�v���1e��A��qp7��Jﰾwյh���ut���wi��Օ�C�p�<�=nٵ*eC�z��:CN�\���ަ���&��5����4��C)p�;Cq�X����:W'(��V�.h���Q�u;DL1[y4;�_uu^�d���*{Wۯ��:�fz�B��jW'�W42#@�������X
pˁ@�O:�,椎�l�LՒ�n]Z�Z�_7�] ��끜�y�{ݗ�\��K P;dE���|o;�﹪�f����k�ci@H��1��h9�◸-��w]N\qI;U��s�_c��eJ�a��b;P����t��ֳr�� P:$��ќm�kk'���m�&�)h��W�j����x��U��t�y$��RX7�gTb��yI/����:A�tmgeG�q�(nv6vv��-ڊZ�4�t,����r��	�I�[Z7�Ф�`:q���U��D<}�¼��o˅oZf]��y=�+@�+�{W�`��Y��"2�Q�&Ae��4=��Ή��	s;�R��]!ɍur�����ǖ}x��9��m�n�����Zٶ&�/�V�
+�*�cn��o;x�l
��(N�v�˵)��(V���{p�4�\v���U\�G;M���V����]r|kk0�v��,�X�i�D��"ؑiޱ��j:׬ݻz��xd��c��V �L5�\V��΋��K5fu!�ã�۸y�27maӁ�v�ɫjV���*�|������h�ˬT�)�أ�8�W�i��R��܄kFAףW-q���e��0dI+YM<1�I�y��oC.�n�`9n3�%�����:�mc�N��ۙg������[���xr�X����b5H�!�/�U��`�{�v�k&�W�v�YtT!T��Ub�&����Zx5Cm�ݜa��!�pX���d&��²�.27*(U1K{���n"Y�.�4�IW��ѧ/�lq��@��W�p�:嗓���ͅ��ĔF�ňL&�v)�8��j%9�d�ì����P`[u�{*�d�8EU�]�E.� �%u��Z;�yq���%ec�t�+Q�&�ݲ]"�u���5� �n�;��
��gV�Ch�V� �nk�o^�����*�G�8�����$����c�K [v��l�l}�Ư�= J�x���q�
Y��	���uK��}X^�([X;k�*�YD��
����8=��6����qx�08��7z]�x]�7Z�Bksz�P��S���z����K:M���b+�,�#��
>"^������Z��l产5��Eǣ�M^n�aD�Jcs2���{m.tz_e�~�\ܢ���6�*�u3�}�tXi��J�x��z/:���o5u�.�ެ��VT�d�Q|�dhAXxu=Z�;}k.%5��>��º�)b�q�K�'5<��j#�{�Q��hf�	��htњ����7����f\Vb.��,"�Í*�c1tsK���E:�gF7U-�W�s+�	��ԗc�6��ڴ��G��T�t�O�>�6ҽ��êY�c���7�$�t7���W���>�l�	N�o���N�b#��vWh��G�oh�(ᔕ�$��!%Y��ۍ�};��;�c����Z���e<X�}�um�\�B�E���u��C�˻W,�8,,�Gr�ks.�����$Voc)|��ܔ��������K����ӗ�qct��s�eBLy��u��5o�Ń��.&�bá��yݣb��W[i
�}W r��mvΨ����K�0ң3��A�kU`�p<��mn�/�1u�'�w"��{i�lw�i�:��N��Z.8+�o�T)Q66��VD�{_b�񽶺�v�kzS�tuv\CC��g.��
���p�/��v+��r�/��,�V۲$��y���c�WۜG�p����̘��;��˥�V*r>��������wx�=�p�T&g�����R�uC�8+n�G�M�����p@M�w9�x��e}�jCyϖ���۫SiT����^=J�o��nk�GH���@+P�ƢE
�5� w�dťTT�����>��܄���@&$��ŭ��qb}a>�������I-Iml�!W�S���2�us���܎3X�r���vF�YN�殳�F��:�F-WS���sp�B�����C4j�$����m|��-�S�Ύ�M�Ӣ�9Lqؤ���ZqԾ��]c��4���$���s�)��Oz��]H��m}&A|w���S���3��`�C�(����1)�K���8��]b��]u�l�j(�}�W<#) ����]]�m0�=Ss�6;���MW�W	��ƕw@�f�g��Ʋ�{(�����}�p��q���^�C{�<�{�g��RUs�@Ȼ U�Y�շ�t�Q��t���!,e7��Ԁ�I:��{�v3����v�\_]�[�eiN�ox�/ųd*�$;�_k��02�ar�V��0�d���Y;�]̻b,�5�l��]����͜���8)I#�N���/Py}X�s�����u��D��݃�9����Y���F�tk��%�xKJ��+��sY�u���k�P�9�K�Kf�Bb���Y�#�4��o!��oxqme�F��N�[@cM�r,&m��0rCǕu��#��,f�%ז�gN6�$���
�QtR	>l���O.9�7+�8I�v���j �ʸ�oUk�uh�m�s���t3\����� m�h��/7��2�I��.�eN�yD��*�u �Y������m䲸R��^o�;��흜c��`��V��	� aR��.�k�U�M�Fd�&,��G%F&�`e]�Y��b�ƭs�rtsQ&����١Y�VPc������{�*:���y����;v�ap'�<�������{R��d�󌉻��-����E�є�G.��
�G+~4�,�4	������Q�k����9��_s%������E����$P�����3���� ��+(o%��;h/��]�S���TwyV��
{�Y���F+N�׽����df���9޳J��C��Y[�7�:������C��-��G��L���|�Z��ZYǕ��q�:"�.��9x��㓖WL��ö�+���*�2#YX&XǮ�w1��a�)�u�N��)P�d�M;?ho%�	Q]c�|���-�ۦ�6
w5hW�L�(T����H0�J��B���T�*�E�F��l`�[eN�SF�U�"1#Q�MN�zVe��19S�Ĳњ�O��c���(���8�h��;6�:Wr���MC�a���Vf�M����ݴrG���α}�M�-bmp&�l�z#[6��Ϛ����jc+���9�Z/�Ҧ�/G[H��#���̔{x)Ŝ/W	|~�'%����օ��ewa`�Z��Ď���ߊG(��&�@^�{&+4�v�]��\��hR��Ҵ�e!�CKFbRu�-��cu�`�t�~=cNR5�H9���L=r(1��;�E��GG�E��C�tGU�=�#ܠ�,=}X�j푍L+Oyj�:L�c�����G��l*���B֖�gR"K����/����d]�NU���G=�۷��5�ak�}Qd]�j�-�;���vf��L�-T�n�ݡ�q�B5�:=�t��r�C���q���J3x��eһ*�ϛ�͚���j]F��yH�.՘�[w&ݖ��xu
��_ �k�:gvu�G�rvh���!��ol��H�"���cywB��#��(��"���]|��V�!�v�'k�C3I�S��txd�Q	9tj�F�WY:���=��)wBa�evf�L�RB�t�Ep0��/z�f��r�'M`��n�ǩg�[��;Aw*��f}��b;M���W���LV�WD2dIk}dw1���2M��!	�ѿ�Ӥä�vMũn�m�̃"ka6��yZ��r��`+�+
�h;X�WbT;�;1F@wͺ*��D�dhZ�ۃo�l�1���� >��̿u]��`�P�A��bz��*V�5+T�J��%��׫����皧]q5�	�kym2ȿ���{(X�o"�b�q�2��}��kX;�s*�犴J+1F��j�k��O�3ق.O�YM�b*��fiܧ��V��]��;�+�IҊׯy�(F+����vޠxG��@�ຸ��d}K�N�u�s��
;3���yG�C�ʚ�<Y�<W�B�v�H�;�ux{t,�1����}�-v����v2]�cR}�0.���j�k�,�]%�����Ƴ\R|not���|��J��#V�+�!7��q�rj�w�S1P�Jk�4#���hsq�v�I�0��Ҥ\&�>����o]�M�
�����2KAa��7�B-gܫ$|U��hQK�=�6�y4w�۽j�Z��e�9
`UGmib��!_�	�k�59��VY�e��\�]	��]�u	C�*· "�r��2���^>�Fir��b
um����8��f[�<"��Z��"X��R0�E#�NU��R@��(!Jb*T]h��]�i��=�[ۺhW[]�S)���hʼ�R��8�������ChوU�g������[�of���b,�ev����5��UE�]��%.��@����u���3˩7շ�#Q�HbY�fAv�F�ne��`�H�\�%D�V�fl�mwRa1���Gr��Ʈ�b�<{�R^�
i�m��F�]��c��ԧ;�wܰҸ��.��Cp����>7e:��Ba�k2�Z�e�Z��6���G���N!NIK	R�e�wv���� �&Wg#Ķ*��5tʗ�oع^�:��B������ۈ��=���A�kZo��"�����¼����+U�!N�Zw)�
���[=�0�6�������J�͕Ȑ�rhM���.���E[�sr�U���z����_k�e�d�S��rʵ{)J��1\Vemև7faf�0[��$��bn�[��/�'e���������4�]�hV{ Y��ͬ:��ZtN	,�/�к`ڼ�����m%WN��GZ+r�����tZn=V(nq�ƅ�-�!�y��޼C���-��"�y#c�(�{�v)��|����#��g�;}�w��ެ�^�{�NE�z�Sv�j���,��V{�;1�nR�j����gV��/�l-g�&���J�,5�����9��2j�p�l�]s�G{�9y�&�r����;j�>q*Fi�yj,tpoo%�63YÝKz��:�bٛ+��ג��p��]$i�ә���ZF�u�Ӷ{�V���H��k4h^��L^�n����vn�\] �ب��ptj�ͧ�ʕӯSۀ��k�f�\�����V�r�io,ѽ��r�0���̱�j
�[�}�i�t��O���ެ�� (�.es�q��\���z%�*p)yWA[q���+K̫φ��e�WW��l2�aڄK�X�v���+D��ԇEʻ�˷k�Coق)O��ҧǪ6�α5�ܒ�s䤢\��M-]����[��z�oMɦ�^�����U>�}��=�Ɏ�:*�t�X�P�o^EI�(m �zp��Ď;�hx�uҍ�ͽ]2����S8�U��+�Wx�_i}z'L�S����*�ဴ�Ȯˑ�ls����Q�@V�ʩvn1�:0��n�<��j2�Ս����,��U����dE�J���9[M.�=�B��Н����w��[��V(��cŀ���w�����ҫ�0iŏ��9��݄��G�u���o����B0���mP����(�̷Y\�]ՒX��}�vqR���9�sP�VۃF��[e��R7�1ͩ���n��Ϗ">@�̤Ewg�aa�����o�l�:����Ǉ����p�Q7H}>����[��r�J�,������J6=�����<Gp,ݘ��Ci�#r��۽z9�Y����$\w�sK�%O�.m�{��i�Mf�Nܮwm;�8��8�Y|��|}D�����23a�m��=�����&���W]ԧi�6�(��bg��lJ��$|��g,�Δ��feG}�Ow��q����Nv�&�膚N��T=u�S9:�VI�jU���!_gJ���b��OiMѸ	M�̔���Yv�Bih�Ӛ�Y�|���q��y=z�1��5�����*]��^J2�^���X�+Lfu�T���M䨮�k'�U�M���,At+)���Zt1}
����ɫj�U�kB�q�γk��DI趃��\�S��<�2�w���nN��t�K�{�(bJݽѝ/b{�����i�W���i��ݜ��K5��j�;e�9�]b�:2��N��2#68�Ef�v�����}��(|�9�̭�
�L=�\���g��4��Η���ցA�ˈP�=��SH��u#Lb�r�\5u7���B��*믩��n�I�����LIx>��Is�״�W`���u;u>wVY,�M�R}o����'7+Q����WYR�G��rI�i�.�w{�o�V.�7V��-s����3��i�����&�^\�oK���:whJ8�\�1
�l|i�ح�����_�<9ߝ����� 6����m�������ɏu�Up��x���괇a��P��;����tA��ȷ��%}s'���r/e��hs��t��R�UgeZ[�ֺ@��u��퍧����Y�m.�n�1]zݰȬ�	�fˇs���\�����zΥ��lE�픛$o(m�f�6�ɗ���g�/2Z���]֦$0�㵁^�]��GS{������Wm݁.�
o0�[.���>���\IC��C�+�5[���P���/�)S�um�e��B��xM^u�،ll����)���q��
}�E�q�F��M��E��H�wp�Ss���nI,��ʋ��Y����;��Y8҂M��y�j�۷��Uy͎��ث!�j����skj�>���_Dzewֶ;0֬���$gӶ�n�h������`«�����Emɣ�!�:���ψ����{j����0����uZl��d륧� �㙫N;Ë���W0���� �X�)�Je�����.��W���H$�
�/e[�H^������hXy�:�����V-xh'�JoS8"j����\�f�Q�׽Vt��9�&;������"�_Nj�>�7y�Ғ︞&i����n��Y�]j�x1�f@�l����
��eĘۘ�Ԧ�쁞2��;��t�Fn���Z��Q�
=z]	yV�0�
@�,j��s��7���n�Y��(��лg�o��]��h�:��<m�y����-��qܻ@�|�f�V�7
߄so�ᑹ�;;u$�v�u=��xMb�6��� �t�mn�(�n�1,�7�L�r�U����N�t�@�4j��'խ޼�ډI���y�]�R��,Sh���[�4�ݚ���:����"����L{A�k�i��PU��$\��gA��\�I����x�5CS�g�]k���#4*J]Q�T�{�ɯ��Y�J5��o��a�N�)�؅֤����蚎a�nm�D�+E;��}�mI��H4�͍F�T*�ͱŞ���(l�i>�����{���ʸ�M��$E0��<&���q<����b�d}�n,�ӍC�^fN�h�Vl���O��>�o��D��u���4�)ݦ�Һ��
��V�6�t;�q(���� �ʥK�N��r�0��]kB�ue,\�� \۲�#�͗df��=��a��II�T+I�`N���a�5l���tx�u���;�$�V!2��ɄIq����m;�V�Xȶe���rl|�@�,e��H��-�u)��4Q������L<�}��J�w�LcNb��B���阕��u���0:�'q�F�4���!&�N��e�F��k`�x/2R�ΎRw[s*/��Xw����eӡ�� �ZR�u�o
D�pcjD��ׂ*�T�*o	�l^)��D+7�-�w�\|�ps���ݮ}K�� 7q�*���:��u�T�ut&�Z���Ǝwo��U��4
�T �Ĳl妵�y9mNb&-Y��:�����łp�|Up�&���5� ٮ�dp���,ud�;��k�����:k`��+���3�;ʋ΍��nR���I�"� YT �0m�f��P]j�B;���kv�}
�V5.T�K6��m:�>��l��U����s�h^S滌���J�ړ���紣��3���__SP[=<+�'�t�f����y:�T3M��}�V9g�s�Gk��]�dMn�o�n�d�:�y��)�vKٹ�������n�c6'��IF;�2�=���0^c�-�*:b�펥o!�ԕi[�!�_W[rŅ�k=�`�t�J&���:,oC))8�{���)\J�\0����Wp޺9|���&"���v���_u,���%�dN9]WWX�����Bn_9A�9Kɋ��:������&V��Țf���ʷ��?�����uB���trmʝ��5�Hz����uǨ�̾��թ�Z��WX�NӉ�(�j:�7�4QB�
u,\U��X�JwEg1���K������j��ǉ��N�)Qu�+��/lh�٩e��!��ѭ��v���Ц�]! ��7��\���ݣ���%]�O��<ǒ�[���l"^��!�XJ�w�܃����8��2��E&��&sWs�A�"�޿��O-ԳY��^Bu���EL��s�*�x���R�����t�,u6�5���d���GM
!BV�X�b��L��7[Y�V=vA�6�N��=��_w.-��e��}��r��kycRQ��nb��c��w�nv�j��Ǹ:��ƍ�e��k�Yv�kf��`A�3]�j�p�qY�/�v�B�**wq�:�$���}V���/�.�7���{O�j��fq�f>��nTtl�����X�_Z��pz�����^��	S�,�n���*�U!X�J��w]bn����c��E*YsX���������)�/"�ȁ���Ǡ��FnT�4�e������+aU ��a4�23��3i嚔w�:�5�ͫ	�(�lv���p#F��+�$5�a���ɪ�T
��uy�c[���2` �(ώ�]�.�_5� �';Ew0�r���CEeeZ�V�N՘8�nVՠH�廵ƍς9�wD������ Ի:�<ދ9�N�FUƖ��퓥��gA�)Z�&�f��r|�KzqܣSo���Nݭz]GV��3WPGY��j<儞g`�	�h;��,q�	�8��h�������u����-�8�F"톕�	K�[��c9��e��tWn�C˧�K���a��F�ךG���'5	A���ۤ��]�&�oAaW)hP�o�v_���Ƃˀe��7\����
҂�7;�6�COn"��y�n�·.����k0��U�\ђ���}��&Q�+=;7��-L�@���Yҳ:؉�ӝ�:}4	\��F.�,���
���V�r�U�c%���y[��U�{�pig�gj�Z�!��c7R�:���	��y�3�:̀ 9Ծ�Ѣyk �j�<�c[��:pO�qx���\�
�2�v��]�o��� `
y���%��]uݎ8��X���e�i!�p�Bw�w��;�]5mqJ`�u|�s=�JP�l<�F�v���5v��Uc����9��L�u�a���].���B��f��z�p�Z7v�ٳ�/�O�F<BYC�qAؕ��	�7�N	��ps�!1��C���=�Yb����4�n��F�}��K���IG�ܚ�}{D/�E�_!��ԕ���\�����9��.�v�ְla><��.�_
\ݫ/x.�Wn��IfLkdV�(m������h��.Һ�.�s�Z6mp�q��\��O`�I�R:���-��NA&
v��u�� ��
KD���J$�C0ɭ�y�����[�x�K|˃M�a&��x�8���v�͛�8�nj�,�����bU�Y���-y�w�!���hV�u���J\|J�R%W�̉�?[x+��Ѹ�w�[��*�3v�\5�ڤ1���v����n�%��&bw�Ι�s,V��2����蹀�p�)��ͤ�����;�hSZյ��d��.����[�Ũ���.(��z����|���vQ[eu
v���%�������wm䊸�<���uܢ�[��c%���)�ʍNͱ���D�x�7�*��FdG'�YП89v��JНkb�����<�1��>�,݅A�,gD�S�U�Y��r��b	@�Z�c����\iN8,ˣ	o�G^ ,Λ�҄,�A�ٸ�M�9e����q�ȉQZ��]X��M|�Ą�{Lǖ������Y�9Z��ER�3�_l��ٕ�1�T�K���Yv�����L���S-mЮ�I�o`�6�����<V�ݪS��h�BĔ$G�m6���F�$�*�غ�p.fݮ/�9Xj�o�<����K<[�H�p���!&[[N�u�͚'�lZE;�(�ϐ�@.��Ӽn�1���s���ƌ�`�������E��jӭU���N�뤤Σgi�PW5��Ie'�n�����oXT$}e��7\�O3P�q����m�aӸ�*&�����h�"�b��yN5

�����n�Y��Ylh����W\��(�sn��H�K�j<�B��t��vl�F�vxL���A�id�3 ���*��۲���ۺ��A���jwf�B��H�2�]�B���a���K���r��ukkqt�v޺����][�'v�F�	qv�6��Y�![H_9��ݹ��j�!ژ�6ikv�Z�.�v����� ��!��2��z�w.����\��[ʳ��	e��WP�%���ݍ�+��[ǭ�|U'�u��{A��ت�\y�8����Ts5j�%dd�w9G��y]�����l`ߞi+��q��H���Rc����;7o��ZO�|"+���P���4D�ng��Xț˺ڼ���b��e��=���MnY�g3}�&-��%�'PV'yJ�u!x4fVfsT�đm�+���Em�}�j"3���L���S6\�+M�>���$�����;�[��%�VŜ6��p�|��Ðɗu��Ev_D)`U`>ϰ؛-����t�b��F�A E3D��PV3�x��
�Ԛ���{emԱ�uⓍ�nlvh��x%���,oN%�Ǉ;��o�+���y�[�'EuӶf.n���䂄�zBR����_ٸc��O�7z��֢�`�]�! ��(5�;�;�m�,��b	���4l���6E����q5�Ի�Q�Ch�SXIqU����Ib}�h��7w�4�r�ÍU�����HI�B���Vr�'�U�����0W���roo��F�N�5Z�GV^�wγ��պ��&�h�CS1�Ԃ}�-��+H�;m�ɀ�n�S���P�0`p�wX�v	��m�����6�<k^���\'hW)U��ϒ�
�5�ʫ&i����)�9�]�Y�ξ{F�R�[�W�#
�5Ğ���po��OzSP��Yc�%���)�W�݇Zt�fs,�h��wn�_�r����{�����N�G��Mv�|18x���*��7�0�T�Y;�c��ęՒ��Z��''�Qh�8F�݊��>-^���љ.���	��h�����j�i�V/j^�u�ʶ�;zУ���@����]*#%�8����S��Q�/2�N%;]rb3�;&�K�D��_ec�%��c�#���H&+4��z�ҁ������UЛ�2���Ȇ��^��K1������(�un#|���i���]7�XP�+�V���z������cxv�#9�ł�d��\&5e���p�ˬ�f�g$�NVv�ZoO'*�N�T L�Ѷ�;�n�����c_���)����5�:�F1W9��<�bۓ-���R�t��J��\4�^e�{:��+T1�M�]��� ����O8f��ZK"F��}��a�tt�$*d�'lƖ�\z���R�=n�gPO2Z�ή���N<H;�=�˭s!J���;b�K�=�l�5�lc!�M���+"Dv��cy�|(���9����&�6��辺�Ntѧ�t2���Ɏ)w6�ɀ�9��/�@������W֣u;��.ے��J6�����I�+�wr!��9�"�ږ:�Ղ�Y�V>�:|�������.�f���+H�ܛ��r6��m5y�l9���c�v2��W�V�KX���_W�:]/�<��6���3k���� �[�K��ƧyٲB'$��XQ���j���SYU�v财���"٥�uJ<[�X�蛷K���4 |1=v�1��6�2����F�p�V�7�Mi��8Y�aɒ�.�z�^?��h3��w�-6K��wS1�/�.�2��{����yk������C�G���-�B��Y��&ֻ[*������~��W�l��ؠ5h$�o�ߝa�
n�2s��X��u�\��jZ�#u &!���anfwvR[/���j���b8��)}�e�m#!⢦#á��چ���q��{7o�ݙ�5%A���u@�t����mo��=�F�+҂-��n�G<(Es�6�㗩Z�޼'1��;�
�8�$n�H�N�y�y�[���7��G
p�%�ړ�X�T�]����M;x���)* ��]D�f�.��$c';�6���g7r���aE�����͊y���*�"	�ߥa��(5`gd�s�`��2t��nr�3�Rr���b���� v�q\�0Uн �͚wR�P
Elq���tEvua�N��h�y+���E��E�j7�	�H�)9�����/sz�Q+x�_eK=A�1�Ӹu�L��ۧ$��S`\�����D�����(���@�JJk6O4�wwY��)գ�l|F����kV��ۘ���/(�S����˦�=oj�z^e���#H�#�GDlnW�嘨�C*�t��2�M]}r�2�*���n	�N�,p�=K)iNX�O@�M���t�+��V��t��g��\�A�;yw;(�)S�Yb�¾����ɰ0t-;̦���L�qt�wzz�4R��ִeF������_Z��X;�&���
��w��Ԝ�'����n^8L�i
B��xj%�QfY��,�mC�p:�OV(v|%�gJ/n��#lk�W6܀8w9vel�!޵����E(�1�3�Hv�щ�j��:���z�u���I�On�o_ͼ��E�G����L\Fm���͙�S��n���j�=���j6,��1mZ����i�d�ok�m��Χ��D��e#ֻ�����/��N�VT��-⡟NO)J�!.��C�;9>Tt�k�(�>!;H�ٗ��	@�xs=��s�x�Ru2��G�zw��U_}_W�|��}5R{�W�5Y���05t{�����q��u�2z�7D3X	'�X�e1���LG�pgq�4�Rx�����z�n�u�*|�| f��j�H�<d�{F��q�+�I���e���`����_hK\�sڎ�	}���X��50��@b��sC^dOu�u�W*u0^��ɽ�z���\��@��MY�
0s��z�z��o&f���6��r�^�7k���r��eh��˕�Lpnԫ0>�8�f�6��Gw��[�*�4�}W՜�G��>�񊮈��[�`�o��g������>=��*:[YYkvm:K�F�`&Mh�D_^�cQCc:�⃒�b�9�7�=�¨g@��a8
˭u�N���3��R�S�8e�5oU��ѕ��B�1G�:��U��IhM�꩕�M����R#b����m
����YyŘ4��l���yw��>mV�}��ٺ�St�9R�W`�vQ���C�k9��������W�7ud}Ξ�>�)I����Jڼt+�EV���u�z�|�;�����%��Pj�|6�g��gL��z�a!�sVlY7+Z�+ٙ,XYǞk���A�	�7�ƪ9�"C�{b��˕g���[���pa��}�
݅�W��+	Wh�ޠ��X��LJ�݄R���9��2�sy]�n����d�24��-���B���B"(����J�(��#�KJ�*������9AR:���*�$b���q�5�U\�L�X\�*9r"���#Z]�UY��e�.F"ɧB�����DUrBJ
���Y��R�*�Q�Y�D�*�I����9��EF��.�DU%t(�J	p�3�QQ£�IE��p��""�Ȋ�PV�TAH.s!d�J:K*9�;��h&W9�.\��Qj�i���(�i
!i�DE\�UD�A+Y�j\�9i���$AEDUs�"�;��+�v��ʯ�G.UU;��EȊ(�Q����\���D"*.EL�<�ܬ���˜��vQ8��.(��BȮPG*��i�\�(������X�"(E]\x�Uȉ1�"� ��""	6���*(����9eI�sYE 	 W��}w����)4=�(>� u�F���K���}G0����q�q褖�V�Swz���I⩇����J�d-:�����̝�YWT٭��˸��(}��A|u�o*]c\6�t���ȭ����<N'�=���D�@R�p	�,����v�O]�vm�|�1�Po*���+=��'�9��$q/g{f�wq�yZ�� �?2���V01�ܷ�?���p]��q�%;�w�ܔ��}�`#���r��Y@���d��	�C4Ǽz� �����&ީ��]ͭ���E8t균,}����0'r�ܫ*�/_�1��^_qZ�cE`����T��=f����j��.Y�ɾ�tNΚ�:�Z����+>�r�C^pL��=�ڤ��\�l���,�X���6+Ӗ�\ ���z��o����Ö�3x{����y���������}���hL�pZ՛��PR�`�ߋ0�0�Q�S��Wr�����ީ*V�msלYB���~���+��?1^�R>��o�z �Ret���/��uN��te�ޞG�����U_yQ�ͯc�}��
3�n�qm�F���wckv�T�0G��͑���j�Ё�,db�S
]�X}�V�Vt1&Xv1���e�� z�0�ʘ9NC��w���v�M�a��=�u+It�U���U�D�fa�j�jq]�X�S��4m��b�Qt#kz��h�$�'	d
��_l�_:�Ҍ��r��v�}�:nG!̣��{������B4�ů)�L�+<�� 'k�T�]ƝO(8O���������J�=�Wm?}�G��/�n�˼�sv�WS�v�{3,���v8��Xg�����}��i�6裝��վ�������ݮڲ`	mxKڳ(|��x�����d�sq���c��RU�<��-BL���;����9����O�ƃ����*5�G�1��bǧ�O�v*�����G�+N���z9����fc}��M�7{ވ9���P�����ҴB��l�~ʗ��y��Vz��øe�U���ʧ%�x�j�zx��[�~d	U�*ѓ�)��E�;��6,�yI���}��]@aN��|��<�P��<j}�������AzɊ�FR6�k����w��w[�Oy��]����Xk�3S�ɰ�\FAષ>s0�z=�egK%�j�k�N��TU�����Ά�����m��P�S ^>����,�`̣p�B��qb�G���\#�G	5���e(c�L M�W�y@q��s���0rv!��k�P3���k)}��f����'��n��8c��,1�^�I��K��BȒ�=��K��b�������b5ǽ]˙���ޫ%B1���z�njʑҼi��3n���<����{�D,�ޤpӣ�ٜ�v���<SU����,�L�<G��Fgf�m�=�Ώ�\!�Q/3�4�,��J�t���$*�eU��U�T�<��uͮ�x���=_j����}.eh�������v�u2<Cu�#\�x��;R��*��f��U�he�=v�y]���]���!��_J���`��	ŕ��&l3Y�-��{�V����?O�S%]��5T>�]�pz히nx�^�����/����]oG�<�#Z�&+��;�{���Er������	�`?���xV��E�ӱ�ҫ�Vxo�x�ē��CwƦ����>0$�i���}yR��Wўf����.w����n?��*f���s|�-��^�Tn�r�&�G"�8Z�;hZ#��@�9>~lS<��)��_���k0��tW�WF�*�t��gz:R���-W<�'FI�u
(Cz��|�+/C��V$ʖ�j��dT�8g����ۚg�����ӯS����I�Oȁ���3�1n�*XlX�[��*nL':m�w���αu˺Wv]b��-8�m�s��	�2��OZ%����;�\~u�����u̳�<�`�r�&=��v�(�y��U��ȹ�-To��/��WR�
69;��|�ko&�k�}��n@v�]u �+�絗�)�m��V
�Wm�V��0ܿ=:��s��=\^��6��^�GhMm.]�MW�_h�j�2%����vg6�syPO_MV�fD�O5)_Fw�nh�T�r[6C�����Fm-����%�����Xr���g��ݟt�R��9������: �ʫ¯��So���=f6���X��o���HOO|�W�����<�y�UW�kl��<��&S�mYDI묥��5A0+&o��O�C�K��GW��<�m>����������y�_u�,5��k��څ�/N�D�_L$7�?�|<\��g^j'�:c���U�^�/����8�!����<��S�g�9z��=V=�I;��F�*}n�#�ق�Xu��W�/�
�y�>��u��##�aה�So2sn���*|�\=��D1�r��}SZ��F�u���I��k����j�H�\�^�����t=�f�����>^��.���[*��}(��Z�&�3��"�r�3�P_^n���+̫8ژ�s��yzeP�i�wL1:QX��{F���w�g�ʎyt:,G:�>9&�a�R|�3���ʞ����ve��9�ϝἋ��N�qv�Mx�������JQV���'���.����܎�	���w���g�q嗜�*�R��9C���� �_m1*b���}׹N�|�(�1[�^�ٖw-����/v������0�"|���P�3�y�CϏd�GHFܸD�ǖL�P�6�{�Z�Y�F#��z��>���#}��A�Tmu�Y�Ϲ��ps���4w���`��PyX�N&��k��8�[�;�b��x+�~�����&�Y�'�Ǡp[~�8x!�n9^���I~��<�^Y�nfv�~�L���.��|���ֱ��V��
^ ��J��xm��y]���Az����[�+DT��"K��'�Y=VC=�	W�+���3^��c�*���W����=V�غ���K�f�Ʃ#j�@F� \/G�T�ύ`!������;	�*��]�@�V��i����ɇ>���P��#g7�����0l4F�ח��K����L�Y�E,�J�7C�u��c5c&���B����{}*����P��W�
^�CX'�2=G��Bm?��F�G�\xmV�Y���D�wM�%}�=�g����<7ȿZ����ѣi
>֜�ښ9P�mz6CW��
�y�+�ruX}B��jѐK�m�zI�c/�_��<b�$x�9�!
�U:u�V�|1�c*��ER7s��9��&,�N�c�ݭ{W?e�6���
J�Ä����k;��A��f�7K�����������>	S7!$^�&��jU舻���3�.��Op���T ����ͺ�+nf�:��"-�V�|��ug�o�#��z���&�=�_un=�=Z���& �`���-�)�vv�ux=ܢπ�h�\�B��ݮt��r�~��{'�2W��h�{7��%9OiN��ғ��ܧ^�x�uup�{U���չ�W�N�Z6L�N�[�ʪ_}��y��#�A�q�V���u�z|#�e��R���>�#�����K��پn�h��3|�Ͻc �����b�M����@��r;�yW����cڸ;�{��<Yɑ��H9���_g�����#"�`?�r�R�v�����3x-�h�l�{t�ؼ5JYqP��;t��$A�/Ju�J���+~B�sþʹs���U�߽yZ��k,7mޕk�&g�l����)^��N��H���*�����8v�~\���{M��7^w;��aK�6Z��
�{y���ϊ��U9R�ڲw��'�L�����(!j��_uS�e��4=�2���k�	��Xh(��"E�3Ew�ߦa!����B1Wg��,��y��ޏ�9��������u6����n�
z�\f|��_E�hkuK��|�F���ĥ�\7rNm�;8��[�%nat��Zj��,���.���� )�$9�L�/s�P�=I�������V=ka��c����W��h1J�'�W{W�b�ͷ�3��M*��F'���/5Czn^_��YF�j�uL��e���(y݄`~�N�ݏOW�+ׂ>�;�e���ۨ��ąx��1Q�8��+M=2x���D��p�f�) i�w�>~L�;YO�ok��*�Դ��6����+��+Ѹ�6nT1�<��7�k޾W)]ѹ1�-��t��m�  {�G3�ٕ\�r�J�s6���
Q&�v���U�٨��0n��+⺋�F�
5�~9:��׸<a�D���W���^bE�ǝB��ـ�������z�c{�����������bc�~��·�<�[].�︗>V0���jT����R��^'���^u�.2��V���?0��f��%�R�o7}�pb�\����*Ү%�}x��:<ٽ��@d�x��qy�}��vE��,S���1!�Zk��_)\�Wd���O��-�-.�Vz:�Yδ.�7���e�9`>]p�~�*Tl�&m��3���!���Uō �֚�]C�a�|vk�*�&���[�A�`U�V�Q���Hr���ū�vr�u����c���ùG�����K$M�\�W�Fk��gJޕ�"7�e��Ng�`����z�h6#*�`^���s{���{%!*�����4;�>\��}#B5�����pi�Z��שh��z<;2J�e��q?���TtH��Dm��w�U7�⮇q���qy!WG�����ąlJ.�]�qd�Y�_d�7�1����1�8+&���q9�G��|p�GG_�?��r:��yT8Ԝ�]���K6~ȅ�*���z}F�j�w��+��U�%)�{�c���y�J3��8�p"��^��4��:A�/����6���/eϹ�c^裝�yޒW����Q�'Aכ;�/��e��~T��+���'�}�(E�έڀ���@+��w)�gl
�r�zM����(H�ꒌj�sM��M��4����+��+�2=�>�mJr��Lr�݅���l����`�3agò�\7�Q�n]0��"�a�O�(<ⷊ�������������[0���}?��e�ᮯ��G�z�P )]z�Y^�}o�*\t�۴k��A4��9�G�G=z��2��~�}�U%OK;�׳V�mT:UUg�Ѡ�n�Z�n����rn�F�ب��+g�9J�1������S�a����s+�L7��-Z��q�)`��oeo1�.���Ŕi���e�0,���p��Π�C��:� #z2��|�%�v��Sy~�F�"NO�x�O�
X¥殌]��d�;�3=O�N\d�=]�1U�׏��N�Ӏ��c9�}������M��_��.g�s~�ݡ�Q��s�Ũ^��M�ק}_nd�텣/�Zy����R�px�\����&�c��r	��J}���qQ���.wk��n�, �<8�3 T��1��E�=��k�N�w���n
�sk��v�}��z�����K??	��㽨�C<��ص�dv��׻�b��W�+���U���B¡�;�y��I��ҡ�=r雤m�U�Ͻ� c����cw�j���V�G��A�=�^�C�J/~�0����ؽ��|���Q�^\9�~��H���K<eQ��v�H�	H��a=��|:��<.rP����S�8�B��F�gV�|�'�=�,�ާ��`�\=vOGk�x�7iT!K��"���k���Wz�<������X(� �w� ��~�	E
ᮼW��"=�5�/�=��at.�� �-:��O=#��x�ƽ�͆W]��D_�ϕ�d�TMZ\M��F���<�4�A��:VT&�t-��2]	8gU�N�d��{]K1P���g@]��=w�O`����ܢ*Qvw�oy��1 A���yg�@ÒV��-P���a����x�G�lvf��w6S��omu����ƕu"�y�u4��wb�D��)*A�&uzd�F^ ���=�
5���/�o��|�����}���.�T����֌��P�����P�[ަp��x=~8��f��o��z
~�u���3[�fw)ŕ���pz�df��W�,d�ܞ�kÀ`�����3g���I�����W%&�����?x[��J�>�xxJ���#'��<@��YhS gXW��>[-u��C�Y�7��cd
����p���b��=��=�X� ��󎶦j���g��ϣ|kL���1q���$y7�N9�!�V����k?i��\ᓷ�Ќ��.�t-�:_�7-�9�����5�x`���ٔG���X;t�,�뵷���[v�8=vNȣ��oO����agM��(+5	O#�s��t�W>�:>;+��|g;|(�u��g��?t�R:8�s��LqQ�l�r�eK�g~�57���@��<�����0�����=�� :����h��v�K��S =;��q��������ժX%��z���Ӗ����I� ��d�@
�l]�C��w�M�1�W��d=9V����J�&C�F�kgY�Y��dv�ξ�ؐ�;ҝ��k(e,8�R�4M��'s��ԇ
`̢s�'0W+���W���oM�j�mٙ6 z���d���G-�ԃ��>��ǸI�����N����7�}�Gٴ�ʼZ^��ů8-�qk�@�� �)��aog%���sn�<��X�`��q»uN��V�JA3o;v�J4�p��l��W��L��d�Ӻ;(��[:)xa����q-��Y��ؾ0(O��v,��{�p�{)�ίeG.�u�L.̻IC��7��av� ��#(Np�\���T�v��ZDEo6�UN�.	�����A��nj�Gs��쳀�巍p�i�Vnqͦ�Pc�5*��)n�?���]ڐxS3�f6��ir��-�[����Syɍ�jT������ȅ�v ���&Pb�-V�q��acڒ�ݩ K���O)T������=�ÝB�c���2��d�7���b��u��	�+���Y�P���Y�d�z���'u�0,�J ��6��l�V)��֗v5.7���](���c���P`m^7�Mu�`�{����Y��˺G(�՞���E�� n�ָw�t��{�k&��Sw�a�6�=y �RJv�Er�k�f�dm;�tu=��R�����H���k��'&!�с1nt���.����Lw*\��Q��������ޭ=�ˊ�wu�K�����w�Nj���H�#��i�/5�Y�,7�6T.'�q�ޣSn<���ŧr��	�r�-�+Sۙ�7�m�n�Z�_(҃��=����k+�#�_s��Yi��3L��L;���ڱ
�:e��R<���-o[\�Yp�SI�C4ɪv�/��|��#�>|�Dw�^՞�����\=���h��8�3LB��x���̚{�1�Wq��Η���&y9iիc�U��S���۔��؝o�ե0wn�x;J��6[4�2�'�.Ħ��0m���ܰ�QUْ�@$p��t�1`b�c<��1zsv
�q���0nh������7�"��NM�T�V&��c�V���n^V�+vL�����1t����*N�\M��9&�$�i�.��7�6*!�u���0VngHeuEfuC�pE���꘣��:�+���U�d�W&P��:��ݢ˺�����7#��:�g�����QcxVc!ڑ#�~�
�E��R.��ҵ.A�_s��*6��;P���G<Cjrڽ���]�;H*��ed�'�h�8��i(�;V]�\4��T�I��guhIy@���Թu�������/\�@�t�yD��P��YSz�s@p�Cbb-�Y�p@W(.��Ǧ��|�>\���+�Q	'~��^��]瑻���I���(��#��/&j�[y�2��w6ü�Mh�l)-Zr���h<�J�����_Qj�/�;�^ʶ��圧1O>�V<s�k5�*s����<�e�\��8Qȣ���+�A�*+�ʈ��APE8US&G"��QG#���)5H���j�r.�*6eDQD)�����S
�<@�.$Eȹr����9�N2�*C$�Ua�r#��#�qZ\�� �V�Qp�G-�nI"3*aT^���)����(�ȝ:YТ��9��B��#�Ȉ�U���UPv\�)�eDGu�9'YG��Br!r�G=u�pUxʂ�NEUE�(�A^�zqa�Ш���ī�U�Ȉ�")2/Ig�\p�����G"(��
n�d\�/"�%DPEܥ,�Uˑ�	˄ETQ(��C����"���8Ug" ��%VV�TAw)�dI%D� �������HΙ��w��r�*�!�Y��U��¹q����i)X�,S��E�����V�bsm��C����ۨ:��k��s�>����~L.�����u����v�U;<�6D޿����z�t� ,���?���:I��<O���HHo����z�_8��?���ڻ�i�B.:���p�}" �?xG��;���{�ߟ��~zx��x�T��sI�Bw��g������;N��\ǯOi�ߓ���'~x���
������?1߼��ۂ|O���>'���8�Bw�?;�x��Ǥ©�t�����w�?�Ļ�%��u��P��@F!ъ |�ɸ��u�S��P���o�ݠq'}v���ϝ�n��~��O�Bw���7hqS����˷P����r�W�����m�w�����>�{��0Y.��b�]���#��D}�0D���7����7�'i�\v'����N����S�v�����6�NݧN����v��N�7�st��i4�ܔ$��>�q<z��n�~OS���-)�M�������V8�(}#���O�'��^+����:�}C��𭸇�����������;�������&���&���;����O�!�{|�t�$����:�޻�8�$���G�μE#�=���^�_��E�@g�'�zs�����C���Wx�@��9���t���F�$<M{Hv}��ޡ>;w��wC�k��������L.�~��t�o^*n����v��} n�®���8���W�7zm��>�|�֐�v��x�C��!븇���|>'�©���Hx�!���|C�.��n!����7�$���Y@���\]s�hoP����}����
�'�=��~}�7�m�tB��t�]}C��"!�#G�8�LX����Կ��F:W��u�;���{q�x�8�x��s���z�Ǐ�>'��aWv���o�I�������  :�@�?}G�#î�_��<����>���?ɸ��H{��z��]�4�|���v��'���ϙ��ӿ8�8���}ｦw�ӏ���t�v��]�?��������q���0t����|��a�'�~[@g���#�@3_�כ�j�x:jݣ�^� ����8��"F C�����I;wG�wn� O���v��J��>o���<C�azC��u�+��������M?S�<�{�
t��������n!;��o�[��
��si9j�ݢR�ip�ّ��s�b��*N�\����c�wn]�k8J#��u5ԮīZEv�c�n�K/u����:W��t�;V�Ok�!���Y�d�}hJ�(n	@�쉢;1�p��:��T۪k6/�tg�=��1�B�R���k[{p��JOLḮ���̿u,�N_�	֟�� �C:��=&��?;t�o�����a}q�x~O���:������=N���"�W O�@�����!�'�;��8��q���{���Aw������PO�<��Փp�7�}��}G�������q6�C�wc��A�>\L~C뿐�}�����c�}���;~wC�?}}>���4}���E5�:�姸��G�@���B>b ����8e���8���|=���ĝ�v|���7?$�8㸇�ӏ�ˤ:M�	�O\y�;C�i7����p㷬������"�1��H������<�';�^�ڡ��ܯ;�����<>��f��3&��9�^�i��_�`S�n��������0�����L/h'�Q�>����,z���~C��<N&���p�l�#���� Ml/s��&k�3{��>� }�>#�}��B#�O�������H}Msߝ�7�'{��:۾�p����������:w�i$ߞ+��`�0�'��8�&��Y�?���?�C���+�'��of.�fQ~�?Y�}�aw�y�wh~O�q����q ���n{��I����|����;�s�'$ߓ��N8�~�q��)���!��=����X��" �`~㗔���d��7ysK���c�#�H}DJ;;�7�����x�#�?�����|:��i�O�����t���o�I������q@�~�ς "��yOg�?C�n ~K��z�wH~M;����z��ۯ�~Ǻ�Ҵgoz��DH���"�p���$�o����o��ݦv��O��;��M�	���}N��	ަ�������GI��y�G�n{m��t����@�G���3�G�� 
i����G����^��7�yo�#�(DH�� �{s��P�]�q���2� ~I���un�F�L=ߐ��wI�y�������<�t��$<C�C�bM���x���$}��#�� ����Q�Ǖ�z��s�#�|Dx8Y�>�#���~u�����Y���b{C������|���!��{�}C��wc�t���q���A}wH}>�hD}�
�v<h��"�׳�NJײa����e����0crʳ3v�գ��f[�d����7^,�(M����59��G��
AՓ��P���8/�{.#��d���w�Q�/�τ����9��жE��[��K����]��;��g\p��D~��Aq>�[~�&��S����N�����z�Q�\w��N�C���S�]=�$=q������>�i�ߟ}zM�t�v�>ۊ��I���9������׭9��+�<~ Y�"�����O���;���@�}���]�5��ލ���	�</�z۴>&�Ӿ"�����}{ôRO��^>n��
oP��<�����!�.��������L�m(W����"�|�b��0˾�_����'�	\���t�wi��7�?�t�����$��ߺ��۸��q>y�t��*��c�������C�����x�ɡ���j/ԭM�>�w�����?�������ӁM�>];�k�����۪���7�n;󴓎�����@��q����:L,�`:}s B0��ݟq��?a�Ϩ�d1">��ڢm��c�~��+����{K���n:C�x����m�Aw���~�$	$���t��;qԟ�A뎕�w{�~C������`��Hz����v�pN�����n�����Gބ�>��h��?|1�͊���f���ίm�a�?�0}DG������C">������ߓ�㏧^�+��&�un� ;Nx�����wg���N��7|�ާNӥw�;>�I�BL�A�ͨc�>���|}�/z��OZSk9�oy���H�8�~~����0�!�]�?~�j�S}B{�������}��JnLXG���{u
�$o��cQ�6'�mz.��ۣ�ަDnz�Ӕ6峦k������G����ֆP�9�{׌gK��E��+�vۿ��w��|����=Ԅ�H���y�+n���nQr\�^�\�F�3�:{�ތ�ɽ-1�&������>y�=�]�nmG�LǖL�k�tC��_�+Ҙj�Z����/lY�X�pxIsT*敠��va5.h�o=p�y<�ΫVX���PN��n���.�Pv�e�}X�o��O�Er���d�$.��*��t;h	z��N�P�;��P,K����o;-gm4��o������*���mC�^^�ٵ���Y�%���*����U�:%w��S��~䮡�
��;��������,J��x鰰w]d�`���g����)��u��>�!��l�YB �lM��{2`�]�t��Ʃ��r���WN¤�^a�&�.��W
�c����\rly�i)��T�"��$�:��N�4�&+�h}�3>x������{���o+�7�2��Y�5��[�͛�yP��e� Lj�Tf�����umGw�HWB~��r�v�_�^\��)?���s����N�����y�
U{�ᾊ��v���[�{�S}��w3 s�xRBmW�~�e;|��^9�T��^8�w�����Q��N�� �}�]����Y�Y��ρF�`N��m�}x����.�f�9�V���	S�{�m,G~v��=?�r�l��s� �b��D��g�����'�yd��֐0a~�AS�忼���U9n0�g����k?mK�����=�"�IM�B������<y��-N�^�����@�jU��\}�:�kgvC��Y+"}�_�����C:v{w�N.xz��K�����&�t��ڒʫa\���Q�����N���Y�چ��H��^[Zv��q]�о���Q� _5��U/l;��������n����2�.�c�Ι�뫃��YeU#�[��xR�㚳_�k��.���u�����,�oN;�%f�����9�Z��<�A�+�7	�^X�pmY�S����3X����Y/i�*ҭ�d��Q���\-��i�Њ�S���/
���a��z��dy?b魫ˮ��װ�t��3V �Sվ*}k�ӞPp�۟c�s�w:��F,��⎘'"��.���������.����[�U��U��GX8N��]u(7S�	ռ��|R�<��F�¹R����Ɲ���Q�1r���6Oq�	t\�s=ɩS}}i��\*6�r3*��9Y)��@>Uą[�|xa�\/T�=1��U���ח�{�Wq�/M���/}��mhu�w�����ϻ�s���ʻ�>�*a1.��o7�'�a}{�WF���|��V�L����y���a����5(zx�k����̑礷ޝK��K��`��;��^3���YFP���*���e�r̡����u:^-d��xhk7�u�����Ù���ŃO�j%��\���յg%�B�>�+q}��z�N�ݚ^�P���1����۫!;�{�1��+F*,Dt�PΖ;i+b�v��_1��d���%fJ�}RY�N�4!Kv�z�;�qf��z��3���> S�������o���@{�+Y�\��n���ِ�e������Q�_����d�:�@�}���7�ZN{���G������ہ��C^aSO~(T�x<̔V�/=����]a]��U"L��]v!;�*@�
Ϥ�@��D�0l���ʛEk5��;Y;��@�s�^g���r�@�T�`�0�͸T����q�xY�4�+kJ�-7ҟ����U8�l�|�0�T�e�e�Z��[T���Ξ^g�����^Ͻ���U���֮>�J��3���hd[�ib4�O�+Yϼ��i{O^�+׏��ڻ��^����g��z�]���v$W����\|�G�
�<��X��<%ZU��}��u�:��4���z����v����cݡ3o�{�k�Y@�.ƹun���g��0O-�-.�ً�z��5:�<�^ǝ�&�x2w�.ӟ\K��ꮩơ�,�K�]_oO(���O�35$|�o��4nD�����M�Ұ{�>Η�o��"������ⲢGX���@xؖ�M�W�E�`Q�C�tMG�K����&�<�\.�Gv����U�7�ݼ�d�YG���&�.�C����n����05V*Cϑ�N�i�C;f�8v^�i@`��R�m�h�Ӱ��V�gR58�v�m�erb�M���p2@F���,r8�v�X���}��|3=br'�d~ׄa�ҳ�\������'W�9��V���@Oe�=�و�n��"�j�Q��S��Q�vN����p�|ym��+�Un,��=U(���g��,=�ci��t������s��򥢰�MG��|��ϴP�C|�:�z��*�x�f̎��f�W/��<][�ť��ϖmW�2Z�E�/@�e��LEốb��3>u�a͓	��w�vR�}.# yu+���Kwp5�.������������q���k��K��UJI�w�4��H�7�wU�b6����^�2xƩ��z�Nϓ�ڕ�G�a�5�ν*�<��y�3�(X�U�[0�� MX��vdȗ��&����:�x�,^�P��;ԍ��R����ߞ`]��]E���7�罖�=}t4]�67r(�ތ��5�;�E��_<$g]*�B���/������ ����������󰢯���)j��H]���G�J�0~�e+��v�W6���)J$>vY[��,�A�ᙓ(�a䱙�ݕ�q�2���ٱ�����j&�5���ʰ�i�0�tW��7����82E�q�I�;M,��iGd,όr,��n�5yh��(xc�b#�jhл�[:��@��)eƧ�\� �Z@�
�ې�#�V�0ڝ`~��ꯨvt�"T�-*�WIu�w�[�W=�_����>ѽ��o�?W��Fe��Q�S;hS�;ҽ���	K��>w�}Pm�# �s��-��ɐ���|�o(�R���yľ�2���3%ʞ앾�r!��3�u>�E%��k�mW"��\#6���os�,	�)(�Wӵ�ا-w�x��C/�U`8�G
p��| �[�t��ի�e�W=�^RY����T�3��*<�S+;�Q�`VJ^lIIt0O��*�s�+�pf���W��4��Wc�����]�N,���E��Ҙ�͞&:��%q�ͬ�������x*�V�9�U�Em��NA���VdB�_W��q#�z��r�;UD���ر��v�P�*��f��|�H����붡!��Ժ�"p/�w�<b���	�V@�"8m|���碽D*e#��2sb�J�h\ߝ��u�D�+���T��	��V@�[�^�~eJ�ύ`�R�Gv|�b�y�6??v5�<��W���]g�L�}k�C>�V׺fi��O���[>��K�v��z��9��	�N��d����XW��(��{��Z�x{Y��ۿs�Sm����5��s����v�W[�n�qKg�5���i�&&*�8�l���f�B���w��5Ӗ�Ɠ�z۲�:�|�߹��������K����&ğ{2�/P"#����Q,z.͋u�
Vy`)�2ln�!W�M侵ɍv<��^7y��8��nK]�"�R�;ȁ����{Y�*[L��j��Eh�d�^:$�O����у�ͫ);L���;�ئ|��y^��C#��e�����B�>�M�8�x��xvX����X�H� �����A����l�k����ڤ}Z�]����9�C����
o]�0��*C�[�����h��Y(g<�_\�Lo{:ݟG�\ގhv+V$��W~�
�>#}ىWe`
���g�g��a��q(+5��EҸƈ�1{��x��a"yw������S7a|x��F�+S[�8�O	�ZU����x��FWmy˝Z��br�}:G���~������},0��|T��t3��Y�����E��kT���՛:4�5�	Q�D!@W�`����U��v嚬�{G���
���W�R�:mfr݉NJ�q�'B$�
F�����ua<kl�ob�ɋ��m�}C��E0 �^D]�a�ʱ��{\�b:�ݣ2�EmzY�(�}�o�/<)/ybQl�]�L�L���GY��x�JyH��s	%��Q\��{���79}غ��ف�ۙD괅[�tpqꛓ��Ec}N5>�x�<l�W$�;�#�	�fb�U_}�}[^՝�Y9z}�?hVeG_�0��S���4C�Ƈ#�F}�x�uj�p�C��.����v��ŭ�쎒��v�MV����ևZ�x�+@n�{"���ʭ���R}=w��mg{td�W�7]���`��_bw6���;���;G�F�Ꞁ���(��{��J�̚˾^���� �oQ����\��u�ue��÷XYFP�yT��,K�ඇf�����wЮÔ']��Ǘ����cf���p�u���
�K+�>��fF�i\5��x��˛U���a�'ؼ<Nϼ���-:������Ɯ9�k�2������7zm��by\�GM�9��\8�`ܨp7�!:���g���Ȉ���O��ٕ\�}���������v�m�v�m ��m0Vs�leC�GÞB8�jj�~���e���&�ݻ��mo���h�H~�����c�Y��![��=o�̬#�hqw�i^��o�o�Ip������DIS��v���Z�8:�_���=jB����:����m�&�F�@!6r����fݗKlrث�/y��%<�$��{�I�^�kE���̤���Z��.�,�w����*�[E���������y�w�[�Ɇ��U#M�w��a�*�����T٫�e�c��-�P���n�ې��k2WE/S����uL<ۣN'����Ӻ�D�꼺ĵ������gC�f�7�WV��>���e+G]J[J��ɹp�K���xk*���Ϸkٗ}�$�brI��ChlT}��3���%U�RqB�We�Yw]���I(ӥ�,���gD��"��1�d:1��D@i�N����G��:͖�0�H<��f'\WIVh[��r2�VX�z��|l�W��1r�L�"��G���B�u��wY&�ج�@����ip*kr�]u�a�7q����mn�sp*��&lS[E>���ʹ��d�T��da�%ৗ���c��^���ͷl���:�sx�Ɓ��]H֣{��շ[W�9tFV��<��]6% [���nm���t)$�M�n㕤�w���	ǵh7S��������F�s�Q桺��y.�Z�ۂ���@���T�-V���a
i�Q��N�t�Fr;>��Ri1P�u%��l=R�9�]SI0���n��<,�In}g%!R�]���&���cd�س�`��&d�)���n��W�EWu �tlqj�83����uS0��V�%R��ԯ�����{���I�,�dE�"&�s�9��$��W]u/e1�.���K3@.�e$�*�����n�_Cθʚ�p��oZ�S�pgsˬӴ��u�֥��̻(;�C"^��W��cPB��;.���A����]��֋�a���o�Suc+1���y�+W&)>���]2S�5�5-�9��KEY6� �M�5��T�2_�&V�[\3�8�8���"�u_*�-����hâG}\�3�֭x�\"��8;(�C���9<�M-(�t�;��WnK��h��-� �cu�(������'�V8i\o 7͎͏z�Y
ˣ�S�]�ڇgR�w�%v�D��R��Xk-�6����bڋc�O�iIf�.4�ױVb�RMWf�t��gk���='K�e��AlǗ�E�RE����b͛��㊬��a�3:�J,��$��1�e��9��U��0Ӻ4>��D�t����E#Ⰿ�:����X������n'R��q,ҫF�S��c65ZV�	<�۝u���m�"�tX�F%���zע�+D��`�Wt�-���ew=��&�i+Ֆ^P�Cymd�]y)�#����/�Z���n��^�w�����8�z��d��;��fQx�򢬑5¸Q�xl�{��{�b�6���T��D�'YS�o��V綩��zw�u���(�Q�ɔ�9��JQH��F ���;�Q�mZ۔�'N��Y�]�r��7���Żf-5�5�(5F�cO�bщ���toU�l�B��P��?��dD��\	ADDE�q%r*��0
���#X�ԕ�$�\�D:y�Ȫ*����4\�9r�����l�ꑨUA�$*�D�T��*(�HTD�V	� ��qĕʊ�W �N%r�
�ѡ�/I�s��G
�ǜ�Q�Ò��t��v���U� ��W�vAD�r*"���;�9\��
"�r�:TUDU�]����X]�M"=VQ�PP��@�%p�dDʹC.E��TU\��Ă��<J��D�UMWI9:�L�i�(q4���� ���1�N2�W\�:zI��s�EDA\�W.:�s��,r� ��D&Qv��AEr�L"�#��*�Y!�aL�l* � �Q�v'j#�+�@���cꊣ�!�uw�� XMR9��3�-R\T����,�}��d�L�g:����#�O2TNq�ws�[�c�k�C�꯾���3�K��]�N��m��nY���	�b��ڒ��a�iWᾺ�qح��{u����-^̱�v�r1��������w�|���Wd���O��<���b�b��N�sw��3���ك� ��=�w���,瀾�t��[�/��Qj�W�oY�i��9=�q��|�N����n}��;���$�Ib>;!���6P�F�s��3)1a��cř^�8g<�L�b�
��v}�jn�����,q��[O�W���W���g�B�{w1Z��+M�s�_�0�؇
����C2�徣�_ǝ�����Z^��F7xL��'t��}VN�<2],��*���P�{��'skW��+(B!�=�BG/��.��[�i�y3�Ō{��B���z}J�OBUkgڶ���ˬxO��Z.��+xvTlpBv�����/��!�Á�&GS0��EIY]�W�uh����'X�A3ù=KL������E}��[wH\f�a "ǹU �;*���a�)~�����T2�j*�Q������	�ֻ��ʵ#�W��Y�ϛ��q����3ac��;��WB�����e���ZX��B�Ff<n��V�H t�K��y�W뙆���m�'�t"7rV��P:m�-�:�7x�5�Vs7¶mp{�E�� �7�5�`�������oT��ɴ�~��\+�,w���6�ږ"μN��CN�S!	&��c9)B�<��ﳻ���n�&�h�,��=x��QXvg��g��<��O��ד��x��>�6�k��v��hҪ�$e���
��. EQ;<%_�0����,��d����+�t�+-�b�a�'��s��\�i�9�:���J�AZ뛣��g��_��� +��U���A�1_�r^x��nx����!��LG}���	��ѷY̾Q����R�lu���-�$jc��st�]ں�,�[��P��z�%�C�ɐ����Z�ǜ#���D�zqIE_����_���u��<�"h��Q�s�c�7�����ל�Ay2��r�uұ�V(}]s����dS����K��h����w�C�0o?7A��Ծ:B":0��m�TTs&��Gtw�,��������Y�C6��`�w�x+<7jc���awO����vK�]��=ku��o��U?yx��,/q�Gjƅ�E�B/���u�>�X�&��RDc�f\�C��]孚gt��IB�uq�S�5����(�}}����"��m�a�T���9�����={�K�����t�+��G'Y-T7]��-n�`�]À�W�����3�{r�ե/+�Kɸ�3
4������]��׃�������#�Ɇ.�"�u�Ǟ#���M��\O�΁�@gK���]���t�*T�]�R���������%��C��|l2/��ßr���w�Cĝn/��NՐ�C_t�>�ԗ?EV���p�mKa��5��U�b�ĩXA���o<%� �p��	5��wB��HV�t����o�t8ˬ,��瞿aO�\0���r�a:�Sƞ���3|ޘ�z�C�`�kN���k6ɢ�'��-[��X�,T�����Y〬��*�~��3�uW���
�EGs��Z{�S:��*�oU��2o�>�����!��x�j�'p�ͶL���H�����ُFW�I�mQ2oo�+�ixϕVH�#�C#=��#�ސ�������G9�QtGgC��Ϙ}���=��,Id�\�|0�N�AS��7{��[�1�V��d���[�;>k����N���(GX0y׍V �x���f_��nႡg�Ώ2����J�ǔ��[�w����ybz��w��5�2+Ӧ�������|6���ɋ�'�M�����n�xJ���9�ݣm�{��������w�m��7��&�
�(﯊�~��x/R�%X��z�n����Pm)��jY�Л�m.,{���]l�$V�&��O�dgS�5`��d�V���oOR���:ݷ��8�^>v�4�)z�W�}�}�֭�����s�(�����o�Jqm������̩~,��ü6�����E��E�PʥW�x�ǉ�_��Jx#��y����},0z��O�w�,3ǘ�Uo�!�ƿ` �Mvs�p�=���ޥ>v	V��T���W��	v���{�t��k	��X���o�lm��ll��`L�Ǔ;���|h�����&Ih0K������xRRZ
�{}��Gp��r�eٝ��!���?�'�Q�L���N�����2=dt��J�z�o��_��	o���4!�`�=_[��*�aP��M�^=�g����,n���6L��b���/tceۢ��"�akxԪX�C��������ek���U�3�"cgP3j��o����k"�v��@��*ѓ♮�n�s��c�����oS'�&K~��W�v&�3v_q����AK���>�&�H��򐺎��3�@+J��V&ֺ�WgRPm9�ǼrvPީ|�����X�w��
��UB��}_Mb�:n�U9q+nM=��'��0z�p�x�&�m�6}9IZ����Ѵ,���]nP]�|��涸�����/�x�S���,!`��q��ő^�^��쫬o��7�)B%��FnF/���:����1�s�sC4s��:qb/+�o,\R��'ջ�N��n5����_}��%lW]-
��E�Y�97��	�(�Q�UΤ���Ӕo�S�ì�1�����4��oV��S�-4g<w��� ��߆�
V�
��	�J<��E�|E+>f�=l�S4��h�ћ��\��>[J�	�4Dq;=d�nrkޖ���=�Ш�\�Ui������P���Z��	�T�aDIO�W�]�'�䩎�W�����ԅc���=���V����YZ߸F{��U�����K�Z ��L�g��N���9���3��g���B1u������F[wxZ���>9��#���Ղ�gQ�]���ec�'��}��VH��i�{qٴ�'m��n��l��5����흌��ϫ�[���[�-��!wc5��bG%v>y���]>�M�Ÿ�v���K�7�D.6�������;l�4jƏ�}"�h�n�Bd &�\��Q��m��<4��@\���=xS���	E�po�ҕ����:�<3�Ywⵁ��ņp+���'�||)�* �<�JK�.���y�ݿ(����MeKEN�uΦ��.5���cǔ�i�X��,-��ռ]��kU`#��Vګk�{C��<A��w��.�nX�����+�����ʌ�/�&�Xg�MghW:������)����<AnX��)�7n�61$:Ω6u��E���^��3��> Uf �<ߺ]*V� �;�I�����X]�UyR�Y��}���w�6ʸ�c�g�*g�<��慈��WG��3��D�WZ7���}�m�+���xO��~V�{\цW���X���V���6��8��a�t�,���&r��@Ңlt�l�.�v�^��#���:Y�A��'t���taXr��/2�]�^u	#N}.��V?;OR���YV��ћz3���F���&�����������-�Q���^5򙯅ک����j���=�L}��̧�]���:<�Ǭ�j
�'�o�ն�x=h���,�v}ݹ6\
�1�>�ΰ��hͦ�a�~�3ޘ��c6kx��O�L���vxK�����ġ�,!j�7qu���x�u�&}��t��n��u�ާC�#Oj�n�"��s�x��j{5�������F����oȨ�Co&�B�����z:�ɣX4�9�?7�=R�gv&)��[ձw��g�1�H\l��	��*�G���T�����}ݵ"6����sOw�'��.�����w{��Cf4��g�](T�!�ng_�3q�@���B�Z��N�k�����j�L�]o{p���>��l�
*�̽�&5�agʲ��&I���[�Z5�RO�>=E4y˶�G;c�O�`�$<�^e_K7g�۴k���ˮ��k������_U}� {,yls�%��eM��/*t�#�Nu�v���o�a��P�=J�W�:�X�-Sylߺ�5�Gy�EѲ;,uʭ�����֏
ϡ�:<�V��#���\X�<-�$�Vs|�L�3�xWO���</.�3�yK͈O2���T�p���������s3��'wE�༱_93�n񈒕"{���Xr�
���BB��3��8u��#����v��)9���q�*��}
���1e͌�.����W}[�#��GZ^3װ��}���^��h~3���ٝ��-H��~/���(�[}oz���g*����}e�ChpN�v��^��:�Ϻh��?�WsH���z�7��%�M�4j�NX�����|xr�&�Dt�'+�}�;m�mҭ�D�lϒ�B������]B�{�)C�<s���*_3�.g��w���`�Ӊ�0o�)�Z�+X��$Ϙ���N?.�X��NK�|��k8�sl��HYYnϞ��e���7��W_4bx�}���������sܒ��c�{���wm����KE�n�r@��M��Euֻx8!�,SLji�_?=�����ì�`-Y�� �ވ��׺��@�5;��$��+:LC����ꪪ�����~r����Zj!��u'�!�V�=I���ߎ(���,��Ӱ�Gg�7����'�±�U���s��5VMGy��h���g!���4��^����dZB�]S��<���N��_C�}���_zWK&x���E�y�0�L�m�{ǏT(��V}����J��vJX�}FqDy��JL��	��ӵM��wӝ}�p55V}���s#��wG�%akA�X�nW��{{�ғ���6�{���p����k{(����+ۘCQ��<T#S�������>���xTߕ�S}�e���f��$��/^1�'>M5kz�x*n��v9��'�ە-�_NB�5��0��|f{�s��w�5� ��Z^�|�ip7�Oz�w��M�4d^�(����E�z�M�깼kЗ|_���d�;�تz|6P��(}��9^�N,�nkz������f��K�.Wt�ٙ�6��P*��[�|�h�zS"�a���'ɐk��k��/�=	�R� ��eK���61Mh����3�ˠѶ����.�|���vAG�����+��f+���������O�_{��m�#���f�Bѫ|�8���}e�[2߃�x�/㦞����u����QY�ky�S�Cے�Ƽ�y�������bܧ��G�C��Od�
d��vw.6}L�~�zp�f��3h{џ���%�ydGy.��ux�����F��{�4��;'Z�1f�S�,6"E맍H'(���p�9����O��g�^��P�v������C{���j]�&W7��0x9���g��^�-߽-`P)��ǗO@���5ff��A_�v4���឵�;���@�ݶr�.߈^ߗR�~*�P�|�K"V�B�JuՍ�-5�$~̝9��%}�y+���3���t�9�Va��r���S�=Ӗ�Ulo$��<��G���%u�U���}{��J�����{B������ܝ�k�ɽ!�vO��4�n�=�bRjw�:���j%;yoK�vp�2��%wC����`��a'Ǩw�VD�^���W�o��súދr��)�\�C ��+��"evp�mj�9sv����]j��᪖E���t�Ve���e��r�:I�mB�Teen���tG$��*]���4�qp���_}U_ ��ېk��3������<�k�zg.�ո"R_�0wTE.�)�S�&�k1x�Z�#�������;�	�jz:wcӱ�iV'����,�m��_gl����ĕ�:zaG��\���0}-N����[2[O7E��c.��V����s&�U�Lv����Y���«{<{�\��vM^�צ;�U��y�'m��i�~sCϢU��Gf���=�9�Em碇R��fm����7}��6ރ���⡽���CyiW�m$�`�d>G8ߴ��T��o+�.�C��	�wjxHt�t�����U�5; ���������N�(�Zr�1��3\h� }m��1(k�#�5
�}�������;��W�.�au����.��>�ɕb��1�'�眆��u���F�i�Y�M��/kϼ�baL��;��:����F�=(���t]-�#q	L�fH�3�:����L�:��3�$5�1���b1�%2�"a4���n�Z���=��5�,�2�{�
}N��mJ��Ҧ05J�\	B��;+�6��j��,y�Ch�e�1��Z5������d�,��rG4�WuԒ��e`s���$�Q[��e̮���ĹrX�O��fk�ڜn�NM��-ֽM����$7��	2U���bN�Y`]�����'\�	kV �Τz�.��SA���-�;�)��a3C�Bi�A�I�Y����1�ƄWn��*E�ʻ�6��mx�� �p���e��<hoC϶��̽!��d9[L[��\��A9�ML�rV�ʗn���!�M͏����K�W'a��<�`dEݢ�vW`�S��(�01���w>��o"���� ��[X�v�Ρ����h���
��a'e�br:�[��\�}�7}�گh������n�+R킲��1�ݝg7p#ɋ5��	r��u8S滎���Vլ��Ѽdǽxr��a�c4��z��S�R��T�s���h�m"{5�m��w�Wq��^jJ���sts�BwR�u�y����H�nN�`ORٯ�/��:�lvu�|F,.غQs��֗P�b�Gf̦��]�(]�Vٿk}�W���AX��?35�`�Z5��C��jޝ�r�м�lJK�C�7GK���ڱ��v�;�l�2�6�����Mݧ���[��^���}�Y�En�cr�X�>��&�lD�X�T�t�J�a����]�a�o �΃}LlԮ*�闲숥�]7�Z���U�5��&�Z�x��Y�̝1;�~�x�[���(ǣ�5��<�V��-p��%]�.��wnk�gp�1���jh"ŀ+��t���ח�M �S9�@{�qlً^j_4���2l'����Κ��5�%u+}��2I qP
�,;��4�]��-q֞{i$sN�i�R����N&q��%��,�(��û�*n]�����td��0�^dwN�>�����\����P��y���]D�����&� �y��}�w/�"����1*��ķۑ�O6c���n�3�r8��������k��E�$Y���*��ֻ�P�3�sq�v!$�%��]���ۦ�֛�u��Z
�s
�G�Ԙ3;i��&�KO��W3�5�D���G��Mӛr۸`�r[TGo��|�N��<�FTg������t�	2�q65.�����v���6 ���-�K�|��y��u�QY[}�-Ea_M�P��C�p�3/6�`�U�G�ʔ�7؝֍��L����E��#+���4uwڍh�����r"����8���5�,NQ��#fd�R�S�Mҋe�0��sH7�9wQWFK]1��͋n0�wμ���<��<?�|�APQQ�u�9w)ET]���.~R���D��PQr ��T
����U���9Ur���TL�Xr�rt��r����p�QWg�!\��ʠ��Q)ӎ7%Tp92�p�Qd,��0��a(.:�\V��QPr�p�ª���S�J�G�G#!g
)�rFQ^#

���D]�x��Q.�&�hQ2��Ja8ؒp�Q"�Pj�G
�';='9�PR��"�l�i\�.UP�iʢ��E���QQh,��#��UY�* �EE����et�V!Qx�&�(�UG�dJ�R�TfG�,<��*�1!s�	Z��p���UUUUTEg����/(Gq	��u�ο�}��:����&+�w�sS�Υ�:�����˾-M�	@"�us���gn�2R�ɜB��n�oJ�Jld�/�������*X�nw���_���4y%�]n�3ݢ��������`��=�))�g�Qn_��?:��}��V�	�g#|�%p�m�3��47/*Y���3/ӗTN�
z_�̼��Z��=��o��b����W�������ӧc)�z����:{i��/lrr�.�kq}}ɮ.|3� �K��{���)�Ơ��x���75���zg)�m^�V?ۓ�(�wN��o�T{����+���O\LEn�Wݵ��C{u5�d��r�GS����'�T�{3��?!S�ԧ�+<�ϥ�	���eS�IfIx�xU�۾J��{���{�_jZ:��u�ʥ�(ǀ��}��Y�<��|�ㆢ�]W��Ϟ�ش�Q�w4�'=����,8g`T�^��7z��\Flӹ��/<�����_���n$o�?_�Aޕ�hs���p	Y�w�[����V=ӯG�̺��uO�U���!�	0g1����~N�?7���������%�ze!(�E�5}�E��O���w�˛v��p�ն^T��w��h��֎K��h�Y�j��Z⺻k�!��o{�F�l*�y��N�{��+/�V���~��t��^ksp���Y�k�hʭE7��]��Cz`b�g<��o#�<���G���E\����y;�'�zm_ɣV��|T��!
�򬝭����W���R�
vUu�I���/$�)���5&@��%
ًv�<��Y�޳�}�ϥ5�wy�1[;U���o��|P#"��L�q[�V=�)G�u+��*\tP{\=�(P����#�V�0s73�oG�h��[��5�jzLLy���X���^�_9���46��;���2s��j*Vec�r�>�i�{5��Sۘqxڍz�;�O�2tr�E�O~������؝WW��'G|�P&��=S�c�Ry����y��u	r��ͬ���tQQ�c�Z��W���F��N�~��!hW��E����{q��b�JnY5�;�e�N�nl���ɸ)����3���ǂ�@W�L?4���I��ڽ��Y�t�m5^��D��ܜ|ef�ne5s�S$��=�f��]d����'�R��D	�KOv$ef�6*�	����Uͫtv9|[u�* ���/�8tJ�Xr��Q
4�]c���YU��ޮ�[/&�k��]�T!ϐ�,u�g��Z��}����I��w�~ݑ����4�@s$�W�M�'�����^�8��<��=�ig?[o���I�����O[���aԱV
z���ǝ��;4t�jǳ`�k)����������)G���-|"ׂ/W^:�����<׽^{�K+�����O3�G���ߢUک��BɵPw�N̨���������m��*���`fv	Y�U�΋˼پ9����2x���,D�כ�}Րm!v�8t�c��[w�"y�|�|�{0K�)��09n>�풮�̩�k�8'{�v��t�X�f
��5�|�$�Ԯ��uڧ+��#<���b�Q7`vd����\�@�}��4z�]CǍ���[>S�ކv���}�iF�F�K�Ov��ٯ�U��^.�T�	�{�הo�(!��^�3��&�aX�+���=��7��zTE�|݊k;s���Uߍ��'�ܧ�[ynϲ�TO�NwwS�8�G\�A�D.���z��"�T�Z�E��A�a[�e�5�77`a�Hxgpr�F���������E�y6������]�d-,R^�J�S�����?}_W�W���=�y{���$=�6ӡ�*�l�O=J`L'�Q`�a?m�<�
H/SC2�|�?b��������7�7�w���cg�����P�x_ڄJ�NM�J�n���|�,c�r�I��?r��{�4�;�u/���X��,��wSyl��U�v�ޚ��wE��VMLիkg�����G����׾7�g��1*�&+˪,�m�����ݯ�ܿ�vTi�Wݸ�i@���R����z��6~οe<�����O>7s���Ҥ/�j�2_R�pRd4]��!�ѱfz�w>�O����E����~S�u�)���<�ٗ�����3���3]<vم�1��h��=�_$���U��sb�Ş�6�8=k;�����=~�ԡI��!Ń��_[�uj�I1�eȭ݆�˟��]���X���}�9���/������jLUY�V�.f��H[�����߳�N������:*���c8_� �»P�"X�d���:���%g�d}�������v^�8F82ʦ���%�u7�rb�ʔ�c��\�qu�u�M�<��_ׄ�zk��4Û�bX�-��53��)fN[w\�I�]������E�6�opgk�w��}��|����'3�ƪ�5�������fW�~|+��k3YX%�q?7|�֧�7�).+���'/�.�0'�+���OO_�ɽLd�}����*�ď{�����^(�����&|��%x��W�;����V���w�Z�^����6�T6�W'Cg���yZ��S>�(=8;�c^hR�o�r�?4�"��f�ϔT����QP�u����
	��u����4��p*K�s�M����w��=�noݷ��z���;w�Ge�ڛ���y�x�X̼��]�-��G*�^wd�w�����ع{<�G�f^���&��Yް�o�{���t�ږl�O�g5Lo�.z�M���V�M9�>�_h���z��}����靲��?��= ��<�oU��F�����}���C����G�<�V56����<�Y��S�v'� v�uL�|6�,��wn��r;.�rq�Qm����9��$�$�r�gj�4J����ͻRh�}|��ٵ�ދ�=��\�6V@��uac3�K�a�.��v�5�wpV�����+�/@�~��:����\�:�S��\�r���t7��7Ɨ����X7�_t�$��v�M/�N�[�����x
:��xg��JO;��վx�ћ7r�T�'Ŵ��;u���{��"U���u/���	��n�^X�f{-�⫔g��H���2T�xpڊ����g'x�<vlu�}!kEz�Z��\6s�� �E���e��0s�v��;U^Ԗ�/Z��O�օί��u�����k�%�|�R�c>����sz�oY��
�y_��n���l�N��r��T��,�ܝ����������cp�k�IEb훎�N��]fR����Bq;�*R�{Rמ	S��p�G2�E��^O���kPg.�跤���N��
���ۤ��w�ۨ��t���2� Ɋ��Ӏ+�{�10�}�+�X���^��y��jݙ�~���@�)�+X�ggR�e>��ِ�"b�gV
�w<U�3<)�\��t��.b����aޞ�.d�R��
r�cGbO�j�ݛ�j�;D�*�΃6�3��XY��{h��u��\���K���e��E���O_=hwT8�ZXHĀMT�7a����ﲎ'���s��B%p�z�^��j,l1�rMwdw�o�r��E�M�:�fz�o�+�h�Wxљ��i�X��~��lqNY<U^�훼���^���ͅ�=_t�q�����J�����J>oR��5��J�8�cPyk^}��+��o Q�ƥOx�}���R��o�ي߁�M��wL���ϻ���[� �S}�T���&��
�*����;}�#�+n�>��u੻�뤟Ղ[���s&w�s��r8y
�,��VM�/|ӝ��>� �i��Z�_k�GO�D�ֳ��{�OyP�aj�o��{��7�)��h,�e���we��8��TS40����*w�6��5o�������z���U���L\���z��y�L�%fv�]�K�z���w����߆�ueŌ�f�K�vm�x�K�?4�����9�.NMΉobVT���y0}�tp[�1�I�̏q �h��a�Љ�Y,�}h�w6sX�Ӣ޽Y���4����_|>f�Dk�5˽�˕��fu|���;��C�Uu�r˼��[��=e�Z�������z=���V�����s�-O�l�]~C�%�r��q$�jQ��W��EM��m.�O�UK�>x�@�=~�t���1:�wLSN6]�iȁ�[}Z��ֻ��Ǧ�
�1@_OAs����厥�k
��|��"=J ��������$.�>k�v�����
�!椯9�*P��-y=�o��-��Q#޸={���py������8.��a������3:s��N/;؄��6�;�:���X�`���7�uюU{��g��2���d,��d����~�o|��3|�r�'\����&�g�wE�^?�0��g۰19`���s$������f�oaӳaﾾ�`��9������}ӻӱ��W�=x�J"͊��-sh,*X�u�q/k�w�Pr=�`�^��P_EW���lMV�}1�����S�WǦ�+������t����I�a�A��w��g#�k�Tю�j��ğ��}X�]2�� ��������}a �v�Y��� ��𙎵Yq�c�s�����-��� Q�+�
y��K��w���@�.c9\�����[�ݖ��+���x��� �^��B�3��Uo�Gqdn{^�z�T����1G����p�>�P�]e�#b��.鷭V���w�<�y�/�?_���9�x=�8f��}o%f8�WVU?-J���bQ�&��毲�!��{3Z������	��F|%�g��Td?/g�;��i�Л~��\���?��e.V2�{>��,o�w����e��#q`Ř@��uf�[���_@�W��`�7�U��༧�y ��W�b�ܒ;ӡOM޽��N}�~l����U���#6{~^׃��&���]⛧�]V���ɽq��<~�E�8�/��-��ͥ�!�B����p�؋SS'��]�=x6��������tվ��]N��(��h}�8�tg�
��9����ۭ^Tu�{�g7(5�6��PyӮ�!f�ןf�W��i���׃�T�ֻ7��+�s©��f����V�>����f
!NJ�}CE+֋�0�M�����y����Ċ�@�Jѓ��^%;5*}gYxubLvS���ՎT5��x��wY�|>�Wke>�wc�/���0zy��Y�/:r������=]Y�<�Ә(b[�K9�	��\�� /}��z����:{i��=#�X'YW˜𨺳r�ع����v�ؙ��;���ҭ�Y���Q�5Of(�����5�Y��x��۽[�y�O��I�{�ٹ/��O{��y�)݅~��М�;y8ǁ�پJ��I�)�Po
��]b��k�B�y�6̊�h�MM5k7�3�
��Z;��W]5�)�h�8��;{w� ���|���y��}��/;u�F�M<�{���n�o�h�q�S7��-��}Z^���X���\K��X�e�������~�o����L��sk�*�dl�ޛؽze�*������wC��W.ȇ��ʃ`�R����Y��b�/h�>��6��|��>c)4jӓ�7ǚRf=7��o։-�(������[:�����{��ɽR��Z=�/�*�6�;%*;e�:�X�!�ىvc����`&r;.	����>=�W���z������� A�e����ٗz��x:�x����\�E[�H%�cc�Ʈ� 3)�e./hm^��(���T+��T��yb�d9|���}5���J#���Sj�1��	����5���P��9ֲ�;N�;Z������{xN���S*:5��ĺ�ٺ�I74���'���@�B�-7�=�M�QY�:�*���)�і�F���܋���Vn^�A�\��.����f�@|s�{�:����S��7{�=zԫ�`�{�Fv� 5bw.���%ЙJ��mF�WP�GyntÕ����!Xv�ݮ��{*�)n��7ۨc6ФG@����[y�nP�ƫ���$,��q�N#���S.,���NT��IN6���s����wTC~��ҁ7�C��A[t�gc֬:�*�aI7��FQ�-�AdD{�ތZ�`�v��z0N��魎�I��z�R5vC�Rt��M��_h��`�ii-Wv��|�YB����h�R�嘬h6�z��&������1Q��[���z4b�Y��48��1�S���4fǰ�5��`6D5$T��{R�֫�[��@M`e`j.Z�֎ܜ����W"�QV����UY�2�r���H��t��졷�&�sm���1��+�iJ]�V��\���e��F�-�lf�ӄ��:�@O�G(�� ;H3�] �������U��s�U��)����� b�wq�.?��۱�@�OD7G#x:��l��Ri9���[�A�Ϛ����u�dkSU�͎d}ff��\���Yac:d|Ѿб`�e�'�l���^}��s�v�R�j� ���ԎI���0��+ӭ
�}K-qNp��&��X�1�B��Vn���$��r`��Euf�8�v� nޭ�X/1����Y�nC�C���s���*�9K>�%�׳�,�]M��
Ӽ�xC�j�R�2�p/m�{��o:1�t�V����Z�mY�Q8��Ba��oi�\T]We�8�I���
�M�7n��7�d���u�8�Ժj��Ȕ)Sŝ��3Wr� &� ;I+3V�"��v���!f���7^cJm�tpᘄ&��µ�M��G��Y��\��euXE�mXa����7�ohs�,0I�b��.滪u��y�1_l����y�a�u�5��\�Z���R1�w`�!��3���V�c�h�;�K�����R�H�����D�bʑs�`�l2���Z#c�y�hݼ�|
��#kउ��C�ż�*F�]
��!�a�R<en>.���Hku�ֺ�"���|�����������+-ьm*�!�_PE
5i�[M�[&�\:�-�H�^
�Du,�W"�����ث�J!��	��}��G{ʦ�gm3@��WP�3��-Y�䅻;�)@vW8�ى�ݝ=�ˎ�z>����b�}�t�"˅DDQP���3�Y�"�L���DQUY),�*�xȃ�ˉ\J�\�
�$Օ/QdU�:��S8p���;@�W
��+�ʪe\(��UC�9T"�Ar�\��.A�qӔʠ��.�L�����dE\�UM����J��"�献\�����U2�p9��TAEh��l����\(��U�*I(,�9%	�P�(�Z�I�-�T\�U�#$$���:U�yP�iK)�T�I�vS%i�AZ�����DTRt�˲��1�r�(N� �U�Nr�:UB���5�J$�Tɖ��ʠ��Fe�"娊B���7y#�Is�Y��w6��%���jc4'h=������@j�v��%|�u�5��e6#���G1-NH��&�UW�_d����{z�_�U��xm_J��&_���~E%�W��y���9Oq��R1��P{�Kqu4���U���jY/b٧���������;�'�~�3�*O/Q�޹�ܞ�$v��l�-n���9�ѳC�Ǉ��VA�[�ӳɅ0�X�cx)��g���z�Ow��Vy�8���/<��z���=���ǭ<�)�1�6����.��<U`�}4dա��W���S������C��sƲ���!v��X�j{�Ǜ�ݝ|��Xz?b��w{^�nc�޴ڝ���o�7^�B�w������u��=��,��������o�L��rnS�<�X{��3>u�﯐^�V�;����ĜwhO��+��zy�s�lƚ���ߏz�Ds/�Eۥ�]^��-�'T�[���>�o�{
���y���=ҫ�-z>S���A/*[�y���~�m�����<���4�.�ɜ�Z�
}b��{
ǻo1e���(��)���R.�]�:כ�*\�t�*�[�3(3�r�c�8Vjd�$�UԜ��.�-�Q�[f��@徻"9�h91�T��>.��g:�F�M,nw���>��6��6��~(����r�T��^��9c��Ga��Z�|�a��Ks�z�ϔ^�Νa��z�7�W���Dg?�_�F��??yBϔO�~���%QN��9�R��_`��6�U�W���3�2���2y=)���ʱ�e�@�9�V|'���"�NUV�Ip\�i�f��G|^��{�A�,�����2�Y��	��O ���U���u�j�X(�K������;f��I��Opl�V�ٓv=�8z4��7Wo��.v���t���c�g���-<V�9��X����ݨ<5�ۄ���Ͳ1L�2+��59��[PrU���ue:�{;���T���Q��>����1�������x7�"�*���V�b(��T7�W�}d9�x+8��&�[����N�qS���w7���<����f��δ`�cv��K;b�~��"�iu���\��4�S.�6�\Y�n�\gAt�[�8��q�6-yR�%}�lYޥZ��,�*A�;��1䮳B)W$�{�-�F&��x�*&.���Z�ն�� ��dW�fL+��+s��Wﾯ�	���/KNߋ]���6fs�-䝂���G��|�w���#���ٙ4���cg�OB�^���TYZ�+��9]B�]��Kh��5P+�zg��]�B���S����4�j�LB�O����x}��>�m�.���Ρ�
�弩�>Ҧ���dX��Ok��<�V�v���t��ngh�b�eUɽ��Ƨݥw��1Ka��=�h��ϥ��Q�c��Y�f��RM�r���y�b�ׂ/U�O��5�ue�V~]�� ��#��P�J3�l'�}2�߷�o�w��>�S�Ku��%�$=��Dg���@�z��k2����n��_C9W!�����-��U���=_t�Wl�g���tW��E�XQK�j�nS϶,�pN�wjK��C9��/k��n�ѡ��z��܌�o�'�ዕ��w��7פy��P�=��K偒p-��glY���|�׏�׮�a����D��E�-^��1�R�:]�W<Z����[v<m��B�	y�xF�M<e>.��C���l,�V
�e��;�_(��w�R����z�F�zg2
Qr��)z�]��3��p�xm�$nj�ux��'���)���+]��2����C��0��I{Jū�X]��C
��V����=�YiH�oޟM��oj�!��@�?U��=Qh��(�(�/��`5
߼���]B�< ������5O�򏈛<�dz����>���|�5�i"ړ�Y��>��W�V(eO�����>����T�v��Ǜc7)Zg/�6��H1��kM~��'�y��y泟9hd[���\o[Ч�˽or����o�kF%W{}Vw�-^����b仪fz��&�$O�%a�w{����w��������_!�c�d�����dＺ�M�;ڣ�ca�M/$ޤ^��������e��I���E��T���j�Q�:�sܖ��Rwx1�I��ۗ�o�`��&Wl�5�lm��m$v�t.�7I\��ݻ7��ꂳ7���X2~��x��a��㢫
XU�]+�Ӿ�\��D���D�N`���8�N����p�W7�f�gO
O*JM.96=Di�W-]�V�+7�AH��ݒ>�p_d�x��-�Q�u�`Ό�jj�6�Js��'|gLt��N��#��r4�fW�*�;7���w���s3�����j�m��� v%{�<5J>���eKW(�r�����}b��"�^�a��ɰw�7����uW8c��5�����y�γ;Λ�񗜪�	��/����.��9�'�^0e糦�^���z*��C����.���O�զ�w ��~��o�tr)^�{]z�
˴���[k�=<���ـS՟]���y�)V�Kʗ�.|��g��麥��}��.������ͯ|�g�����T��>�̛��Q��>x�`]����I��.�/�(5ü��I��4������1ǝ�.��5{ਭ��z���ف0�l
�:���%g9�pܬ|f;�'Nf�O�c<{���1_��,�PF�e�qv�����k[^����u�!���z���kOjys>��#}�rW����������ȥZ�j/^ջ	��N�d�α7z��}؁�Lޝ����r{�����R�{��U���S=ʈN~Ϻ�ď����-�S���E�Ϩ�)��:�C��9�����㒵X�|/��������w���؝:w r�=A�3����7N���߀[���输�
}���=<�w2 k�#��iAu�-�y&��oSnOg�#�s�L��ɹO������3>�{�S��p]�i�靯ɏe��:ϼ�`�����=3�>�*9Ct�.�Ÿn¾��7����C���F`��ϥ�>��n�2��T��'�����^�ݯ;���ژQ��>���yw�k}�{�����̣x.�ud]n~�����?Y���*5���s5�Eg?W�����2��%���I]3;��]�{̨�H�)����5Ҍi���g��V+:,�:`�����*n��}>;�]���:�s�;B	��G�� 3����}y��ў�x�G�yOd�V�����<m���;�:q��x�zxE�<����(�N��[�̒��x$��I�^rvd]E�N��{�R�nm=8��W
!�m�J)�x�SH���57���Y�x�5b�ev2Ѥ���n����\��:����:�G8Ѯ�hu����dĳ�c���Sy��s�Q�Uf�V][��R �l�����V9���cw35Q���' +���z2Ft���%L���e�nx��N����^`��Sؖy	ͭauɼ�_�'�Z�&��0�=af̝7G'��͒�*uZ[��r��	
:>ū�y��s[d��n�WxJ^:��s���n���A���I��JG:������>���g�0���Jl�S�o�v��=��H��=�p{;�z���D�;s��Ϸ�wz��7ӧ�s~ų��Y'����{���J>��`�������^�g�����/{�N�5Ӓ�W)�]y��뒎�4�����Ֆ/��x�=\���{k7Ӷ�����T�M�~���^����̏ڻ��=�+�o�a�ub�_��Vv�&ҽ��<-Z�z��m�6	�]&����e�c���y"/beP��#��
�R�����%O'�ދ�g�'�4�(/�{�z���
|�-����g����V��k 6��<�^�ꖇ@��,�H��u�s+�XƝ�5�g1�$�p���'��b��%q�?S.������|ӌ����:N /�v�Tb�NN�T�P��+��Ml��WQn�g˹�itk:���6�,5m�s��O�
�x/OM��Sy��/ d�݅W-<��,�b��j��6:o4�Vm���d����5�7����3�rP9���4KГ�OO�☘����B|���Uo��fEH&��֯��/:��n�u]�<�~���ֶ�v�	F���.�w�I<R�F�	���{I�h�^�'{F��nY�T����ؽp;�_���-���������{�9��8��}.J�p��9������٫�!���XU��`:�;��g��n�zW��+3��*�U�-��Q����:}�?��&� ���Ã#��7ʥ#ϝN���uޥ�����ԥ.w�lU���[sz{=�	�z\���S���7αAI#�������A����f^s�-d[�[E�I�L�[ys[v�;'i�_{��A�ѷ
�&�����}ej�ݱ��
�Kƚ6��c�j�]�Y�6�n�g,˻�������5 �JfM{4��)V�6�κ ucY�Y*��.k����ag[�:�qm^�.�j�b�H>ˉ�r�CHv�{:V;-��I����qfX�Z��nw8[��.��(�УY;����-��"1��֟�r\���7����ogW3�EY[6�Ӵ�-z�t�x^��s�(+���|���掤^��yh쵔�=\}���M�o�FwF�q��W��Uj�F��|���M*Ù'��R�����=�;�
�d}��ӯJ~�;��}c��gv4�@�f;����^�{�v��{IM�/`}(�o���@���&�$j�Ѿt��i�����|��Nͥ�q��Cq�#1�T6m�����{ۗ�uA�<2F+o9^u9EA˅Q�'���-�}�39R	����Ѩ.�l�_�͗�`�7k���Иxt�t��3���F�]���=�/��R9�X����E����;����1ۧhT���1�}�K�ڻ�]��7�v�Ý��ӌՄ��1u�18w��:/d�wvs>K>�� w�I��������.��h���jm�|r�p�T�t[zr����̬�՜̞�=6]nA��á�6����6,<��\.��p��j�Y�-r�&\�x��Hm��m�-D���_`*�O$�+�9����Y�e/���}UXL���\�tf���NiX�w��˱�]�"�F���7R��?q��uv+�V���_V�vw�i��]U�(��A�޴N��5�AY}g+B����wZ�͡�F��r��%p��!5��L�1�6��x�.{eܮ�Et�ƬG��]ȷ�op�����ij�Ul]�.���'�y����z�t��S��o�E�v}Oܳ��&�n��oblǣI��=��Wa���bc�����s�4��r�5���k�=ᕩ��6D}�{;�$�3[�Si>t�~�9��=<�s�9D|��#�n4�=ez��nE�	hcWK�\:���[C�fΞ�K�k}����~�,���j��j�G�Z�3��w����7c�H�Һ��|���o�������eN�Ւ\�s*4���3�z���Lj��ὗ1f{g��z�����;�Ŀb����T�Q:sp���ܬ��/��-�ۀF��t��p㻤>'r2ss`����ǔ�yS�FV�v�9����UҶSӛ8P��bb�f����F�u:�%�w�����9��tC�输�����m�q��V�*l�Ȣs�m�'�����rl��Lq�t�x��kym�]u�I��qD�R���g=|�	���$�w��C�u�r�f�厨k�H��)PK���
�a���x�/;�͕vjqs��Ʒ9��"TKk����*��i���U��Z���o%�5��^�j�Hn���t��Awo8���#�N�U.�l�h��յ���;�s/k���Ma�T/1ڥcF�o㋇�#��}���/eVk*N��U`��c9��wp�ݰ�O�J7ٴ����k)�ߵ��#9��	N�^�t<-'�:U��񼾵p�^�<�^[j0�qN:ތVfӡ7R���)[����[�7-�0}Į�b�"<,<�1J�hg=�fM�Y�O$��Q��̭��`i��Fm�"9���œ�P����K�u�nc1V�oR���B�Wu�Tw1]��[��ho������l�Q�<3y�td������PZ�u���;�~�(9���i|�4�j�,�V����%�ȋڱYF�]������às�S�W��mV� ��&���������~�l-]�}+>�n�SE���JM2/fX:�
C�Z$��%��]B�_>=��8^���W�%b�Π�b��굝�����bE��.�Wh�y	e�9_9�yǑ��*�fP�tl��'GC�k�mެ�x��+�̮��͝L�V*�5�R?c�ޝ�[vyS�D�[fZK�CC%�t���0�!��Y����P�:Kb���[[���sʱ�V�9��g�ÒeYW����e�+V+�˯Nv�=2��6s��s7�):e@�]����8�G�����o�څZK�W3Ĳ잧�X�r�����5�w�1�5Rܺ�`�ӽ�Ygx0i�^�O{r@��fT]��O��׈�ǯE�&�ib�q\�/����۰eкR�41��9��(�u\��E��s�٫�*zΛ�	����Y�B�7u��nm�Rh�9����Y<�d�n=�k����9!�L�a�,.�tO��oYb���vZ�*$H����(�T�h�~��i����=4X=ٶ�J�O��{3 	��Pb�>j�7b��خ���*i�vI�X�I�[���zE|�j����xEܼ��RF�B��N;��c+rj̙�ɨ��e� ,͉�%�n��Mr���hpVD�M�}F�P��/�Y3N۫������:�3$��g�D0'ݨ�7Ѥ�MϮ�N��K�[}:�Ł�Z(9�*%׃7j}�h����xg|�=x0t�5�:������Z0�k
,��q�H�T'.�(���SL�W*�PBe
��H�*��ʹq��9�8���i2�iˑQZ
�˖^,s���J�%Yr���(�.Gj(EgMB ��$*�hP��ꌫ���H����t�G`�i��r%D�
N
cI�q�Ü�^F�DY�9gJ�$Ê���IEq�I�2f�S,����]��(�����#�Zg(�.�r�:�C��qZJRt�B�;J��T�$D@PRT$U�t�ː�b9��r��aU�X]�]�v"eU�Bt�Q�)$�&�
i��$B�C�̬�8]���t�� �P$�]&r/}[j�s�4�R��'���d���%CY���6_����2�ʼ��qQ�哮j�]����}U�{n4s��5���M{���Y��9�PX�:eG��^�􎡷��ϱ�A[� ��7s��}��_Y{+���^A�y(`�3��g��9�}~��T��x��D��ڰ����u���C��5T�\�S�����c�Vתy�l\@k>����\�O��ّu58t���=���2}]����]��{�Y���^Lr�Sb��~TR�1����y�W�����y���Tx�o�ܞ$v�������:qG��W�~����} o�����v�A������>��U�*܍�TP��ώ.ԝ���I��N[��S�{� �m5�+�ҽ��,��N��x�g�X|�.t����GOw�P�OO��nfs�-c�޵&�엗��խ���K�|��S�7ﾊ{�_=���R�O���s�7��p����Y����S�&U�OD���j_+@e�u�9^�2>�z�TGwb��v���f؛+/r���Y#�xA���Z�85P�z=��>W�Q�n2�з��j��50Ŷ��[:�6�*$�9ٟJ�e��&$�Z�b
o���{y��1����&��y�k���_�9���ǭ���|l"xZ��{��Q�#f�[����L���G�����O����v��uNe�����k����h����1K~��|.Z�y�z�t�rݼq˽{��\�/��M����L��=N7�w'�޶���L��4;����8{�����}�
�]N����\7�yU���2��P ���{c�_OQ͜63��]���|g��ǹ�OW{��p�N����"�M0K�X_� e�,A���|]�W&��`u�.����(X��6G��6u�Y������_L�N��Us�O��MNP$��򼻕(��Y��ޛY�_,/�Gn	\������z�Բ��?U���o@�3C��T��ݬ��]��^�� �ϗZ�����S*�lV}Prʛgx� ��|�U��R��ĭ����k��Ow��9,&<"�*Ģ�ܥf�)\$+]�21�dV�0���gx��ވ���%��z.�̬���ͳM�_WsjP�)�wf��s�ɠ �f�s��f���.on�ꍽ�G�u���ۺxD��oi�|&bqҚN�����T�!\UYY�;�ڟ{b�1A����uyE��Yw��s>��d����jgud7%�e�[��v��{��g��.�c�i�
��|wy�<��if��Vv��������O� iT�
i���u�>���m5��s�-���˪�5�T懛[]���zSJj�s�oA|*GW�����瞯o��.r�*��e��dx{K>�]�;w�!�qy�O��x(m����g`���l(ԯj��J�/j�S�דso3�_ў[��e|zҫ�f;+��v6;յ=I���x�YU�4��ܓ/�sڞ��������#��Iﺔ��60a��# �u|J�oJ����m��K�	���ySw7�f/�v���h��"�{�{/��:6��^çf��j����^.X��Tz�i�\�(z����BI��F�^�O��P�f<T:o��9�����9������y�[�P��ʃ�q�Y<:�w�x7u6�d�
�05ݽjI��wUN���w=%�V����홶��f�]���So'U�m��RK�����m��$.��*:�DN�rT�����\զ��w�*��]�R���6�gԺO�����5�jqZ[�/�=��ѽYj�{:�����-`g*�����!߱���-�z&˻N�O�������z���L�5+3y�\�a�$����(�y�ufVt���j��<��������	�Uו'j:3Hn�Z��m<��ڶ��<����5&/nE�e�Q7�B�F��;��.oyw~�:��C�M()����K^}�i8�F�@u�ܭG��:H�O�^��)�O�7ݖs�)ӊ�#���{��G�uu/m?R�o���ƜޭE�6cN����U篧���j;��w|*${�ǯ֞R��ȷ�b�z���USލ��Ϣ����M���v�냸t�;��K鯡
��_���Q���Nߋ]6��6e���0�	=�ӌ�륯�S���9���j�+g�I����O��=S���3f��������Zlvf���7���1����ie�(����^�;o���|��ʙ�2k���^w�\�7z�$�������[[�)�XO�]���D�Yk^�U�z�6d�<Uѷ;B�O��U�V��$��N���v�9OqCCHw�.��/���4�S��=��?Q�iV��l�{������>>
��hֺ�\��=�ȷ=@�~7^��W��ţ�el��+�k}�<�2x�Y���݉�62?):咽�s�}��[�(���=��-eL���~�8Nm����^���c[�U���G��q~GbT���K��>�+�Ԡ��zAkj�ƶUt�95K��_�G�)_`NJ��; qU�C����/�h�[��q��j�oMfb�x�n��u���:�r	hU�P�w��c�\�p��^�j|�� ���OM�����u�����ڛ�^= M�M�����ޙt}W(%�#?f"����=|�b�d������Wr
�ͨG{9�U�;Q�)���[��̉����C�,��Z�1����~�Vՙ-��-��̍Zc�d=�O*�{:U��T[��ߎ(|������#�������9;�nK�Sx��Q���)���/��&Ѭ�=#�D�&��N\���m��x�3����|����b��J��j�;`��u�x��o*-�+���y�|�)E�hmN΂��+LGz���i"u<���@��н{`�	�^�a�s�+2�wyt�������<�P%C]�lM��R��K�volM��>L'�Qf�|�V����M�Ӵ�|�-����Ō��yw_�B8��=���6���i�oؑ���BN�O�,�KE���7Ko:#�'	\��;7w:���c�z{z3��B�]�����ò[­q
q}�#{�ݛ�8m��[}�c�������C��N�|�����	�I���n'Y'S
�5j�t���xne�8k�׮�Z���^�r��Mo�w4T�=*�����%<���*���ϳMz�����1ܛY��cq�)�_�S�f�*n�s��ӯ�����B�Gz�$����iwu�{1L&L_�{��n�{����<Ī�Os�M����>}�T�VZ��'޲�|�s���-�Nn����+�����d���AV���*�4�$ְQ��^�S��6�Ȅ��\�փYu�{�F7b�e�Љ3n;]W�l{$ޝE����¿Gp��*�#�4���}�H����A�]jBU�{Hr�m����
@��,{W�+�p�+K��|��Lػ�V.б��C:�쪷�r.�EVS6�,��s^%��3g�ס�=V'���Q���yP��JOH[�e]��E���ã���4���Lzӛ���7�2��JTr�+�?�wV��\�?\{�Z��y'l.K�r�� �f�p���-��t��>�^�Rʁ���SD����4��s�����+I�M�X��Ł���������(&�>��&d�/�.j����^PV�.����z�����y�}N����w��FB-����^>�`�=~5Hߖ��Wv��3{H^ڣ�K�l��Y^xL0�������C���Z{S˙��$]c��[���ό=�k�z�Ov�o	���@��%���{[��9u�����=6��)������&^vwʋ��6�ݷ��
�Onu���˾riy&��^�.�Sp�~�/Bꛄ���Μ��u[���]����쁌�M'�M��-k�	�w}b���,XSa��,�����iV��pj*�ڿ`�v�Y�d������4Aq�\��bQ��ή"��j�\��_�m׶���y����#����tjε�n�oN��RT>���-�	mg_���oCu�߸���j�oo�p���3ϧFt:w�f�o����Q�Qɲ�No_jR�6� 7�U#������eB����!r�t�ru��C�#FN�b�8z�H�Y~Cq���t���1�R��䑫g��C
�vr	\q�����mx��xH��ә5�~���W�\��� �fV��ʒ9�K<6���R�9����a��fܟwQ~��{��ya�_����2�r}�:�����rE��D.6��ܬ�\��{�s q���{KU}����t*l�S�󠜩>�й[�2GA|v��t��	�z�ū����{�i��҆ɯ����+��Q�D�Y���'@��2<����L�j���b��a/%ӗr�^�s��Ue��}Y��^�:��H;N��ꢈ�,��ꂓk���RmE}�~Q+�o���4������'j����j��Á3���Ԩ
�u���<Ή����+'{��!8]sZ��;�f���?m�`禋F��������*3z\����轡���z�����3���]�v0[��Lt�}W����|�g�ܗ��3MgG�Q��,g����ɫ�Y@��d�=�k>�^��{���F{�s��6Ӕ6��z���ݎ�]-����u�a�d�]�]��޹`5�^�>��lo�����nA>����,����U�7k~Y�x���+�wB����%+�~$���z�/ê|�8n�LWS�.�}nsJ~U�>�<nN��J��{�N��{�b��k_���ޤf^#�ǦR7��z6d%{LX����n��X������|�*��]�g����vk�WGe�� ����<ωC�FՄ��jw���8��;������c}*U���Q���^=�^�`��'jZ�@-�O\d
�W@U��3zP\n<�P��w��ص��r�S�uJ>��z��y۴={*Q^�2��̠Ϣ:�\J�����].���}y���畱Oӊr�����5un�~�����caݫ��ʢ��BF�by�:�����(o�ᆯF��vއ|W�UG\�&o�2��>�NN�<��j� W1-��Y�VY�B�2%�w�������6�Xs����Z�Um����ngΧ W��)�$��)~,�� ��kw�W��s'WV�Cy�a1?S��7�X݂��M�F��7��'>�S�;��p�s�U^{�ٱ��0�X�.,'r����f��aiM�nmՈ���I����]�S6\�u�[W�R�u�{���� �d޾�%�i����Ǵ�w��X8E� ��Ѿq��ΙŞͧ��,�gG�ڨ�ux�P]��t�0��ي�RN�[yj����ޫM����A����y�&"���ي5uK�!��W����2vL��ݲ�?�~��~Z�u���=�:�5VWL`�(dlϙ� w���u�-u�Of�wu�h�.����R&��;d͇㙙P��e=7V�90�Ϻ�&�4Acs�޹����ד���ψ}���uX�,��§�\D���K�c2��oޜ��ٞ���t]g����e�	�ʎp��2��:�7��[��߿2��V�2}��Zxz�����=���z���t�û�ǜ�S���p'﫩��R�g��\M��.t�?�;�x�fO�Zޯv1��{;-��g���8��t����<���b2�M�>J�m����z���� ���Sy7l�y����^R�^ET{ƽ�H\zg����R��V*/�Zf��1����Q�/�MVwwW��V^tKx�ҕ&�)�uq�_]B�y��Ϣ6�z������kާ5�9CTo0(I�<[�C7._�^|}w �[��r/�e �o讞�]���_)���B]2��!i鷗κC�Q�����i#p�K=��=����������$$zT�}]t=q*��G��<��3�;���{E��#& �ڨVe���5�XImoN�0�A��O���L�q-+ս���gdP���}J�u���j7]:���7�ޱ�j2^�,V�����ι��*�%�5�pډ.����ngݜG� %D4���Q�����eswfܗ�[26�î��ںt�D֫\+b��kxlg����Xc&�<��]�X+����c��o�Eν�=�\��MGW|3��V<��f��ѧ�@�0�?u�+�)>�3$�����-:Ӡ�}�Q��,30:7hb�N�_T�Ӂ�7���E�э�ӭ�V��莅�i�ߺoː�gJ�JPc��;o7��>u�=��0��!-e��\��;+2�.�fإg��)�e�	��٢��F�,��PL�t�#�$ξ����<���-����N�x�ʼl�x�wF��ov�\��3.��q��_*�A٣J�a�H`=r��gev����,ボ��z��� ��#�d7�t(�ݔ�]����ޚ�@�Ct��`�݅v]�}o��{;�͊\�@�����Z�]����7�Z�D��0��p�v"��P%]t,e7�
��;{i�J���}���ۚ�v9�Hi��E���$溁�_��vF�W#�h�YA���c���Ѝፕ�{��=�D���*U��ٝBə��/][s��B�n�rҽ�&��A�;f͚�Jޅ�Mۨ�� �((u �##|�8m��%:ڈ��*^�1�z{~M��M9O����#�n�- k�[8���ڮ�}8�J��)�,J��R�nۼ;��n�7��z��'F|~��G!v1'u�G2�B+y�cL�]E6D�&20�"�j��l����[��r�=�G�ٚ��X��3�$��J��e�V��]ƺ@^qZmչ[�Ә�%�A�+ם���F^ؤ1ei`�e[[�8�Ϧ�%
�֡�ə����s��!d՘i�Ŗ9K�9zP`�溚-�px��h
��bk�wI@���������5�_�}��?`����,�';c��Ԏ�,-�M�f�Y X�q�L�자�]zR2�{�8�{��J��2��v1u3@=9�i����Wi:�G��4c���l�կVRK���r��3-�K�2�s��ջ/p��q
�=���`�{	uj���}sL�:_P�^�oD�����=-_1���
�����H]�����k�L=�2�۠4'˕aJ]c`(�����l�x�e��b6���}���n>�!��E��@�K�O8���dD�������1�qP�&�S%CVf��fvv��fƒs/��M��a����'E]�a��˙� -<��� �$"���مY7���t'�G�iAV�ON��浤;�I;�9��ܜ�p�u��(ԙBK}�ۧh��oD�����$uv�f���	��\!��ktQh�-���J8�
�ό 	���u�s��R�U���ݲy;���Ԃ�͈"���_g��vg�C�� �G�Ii�)�kT�B]$�©8�����I&M&28ŒE���,T
)2g4��.	r�;����t�ԨQ�eFaA�BaT�4��)�2�f4����]5()P��euCYvke!����Т��
*삲UQ��qT�P��BH.���H)���&F�*�5�����Wbv�G"��.Y6]Z�e�:���HЪbWYsS��%p"�T&q!I9HUt�L�в4"�e����,�6ĩ,˨��*���"�f�"�����e��B����;I	������T���9p0�p��RIS5VD�C��8QkI+���B�����L����T[�������>}��T�dt;2�����܁�E���X�"^��vVZ\��c]c��N�ɫ۩�ލ��~XxO���yH.s�a`�|V����>�eqQ�)�-��ߗO��X����R��6.*HײX��Юg�q��>��F����H�(�v�~��*��k�g\{��s�g�׍�8<�[�/��z�붴1{[W��T�z�N�����g���Ԭ9r�%7�$�#pUJS�H�n+D��-��xS;��L/`���\uZ�F5N{�Vm�B���q5�r��-y܁q�E� �B��D*��Y'������@��Q^���]�'��l�{[�93>�.�+�ӣ6��=��Ut�z3+���37C����.$i�����wp�c����B����;���/�:n���U�����QT}����o������p����\IܛU�q���
�x����@Lm;�/:�z�S���42u��\F��d߮Yk�U7�%�{��o)�,�O��FVi�~ɬ7�9�;*��9�0/4{������O�!7�.o���]�u�����1�?e��}��Z2ady�ټR+��e�&+�y�^����c\�?�� A�,]�bn�]��z3�c��e��s�wPB��kY��kթ�Pha���!r�{^F�@� �CW¯m�9w��,���	�>�ɝؐ�_i�fEu-�Զq�!.����ot8���ܮ��t�]�#��s���3w%�V��΀9E��*��v��B���.媮�{ּ�z��X0���rG��P�=3�|G	CόZ�dGcO�<N��in냏/K��v��꩏3�׺��F���ވ�DR
l {]߀��z�_�yLvȭ�]+�ﷱ+���X#���pܦW�r�ܯu�_�YG��#j��[�� !��F�z1��2�tb꧈���CĦ_F͎���(.Vei��U���(�z�Vj�W����~*}�����]�s�.�e̯*-�#7�H���c�΅�N����p�'nၐ=W^��qW���~�Q�#L�sq'�=��q+�b�J���P��ײP�wM}ʝ�*w�܏�&���X�/�;��G�j�{�5<K�ӒB[>�ɡ�U;8J��L&{vanʖ�>������8��T^ʭy;���eȨ�T���E�/&'��DT�(��)�Ê=��۶��]�z��ԥ��	���tx&\�T��^�� f);� $r�k=>�y@�
��H�}]8�	sH�w������T*�e���r�U9�>�+�~�FE�X��Or]����E���}�957��7WW�u���:�]��(n���u�KS��ޮ9x�jOu|�n�*�ye)ݐ�A���9�n�V~{�����u�o�$' ��.�=B^;�V���{I���X�;����f3=�	�; m�xV�W[�֫0��O���3�A�PY�a�=��=7�2����
�x;�?S�MV���~�w$�Ó���0�=�����A��@	��L^uQD^*d�8{��TC}��߷�{{�y!�\vexs�͕C���56��b���0����v�n��*���dݬ�ԥѸ�HNu�>��YF��5S�zg��nV���GY{Sх�_���z�U��uY����@R�3������q8�kF��F�����Hݤ1�*����g�~����xQ��/�T���F���!e���Mu.R���6���nDs��}�Ĥn%�z
�ܮ��N�-�h����3�_ѳ!-�(%���R���{�3��c���9�ԑpR�).�g�g���n/ñ~%��\�����o�(s��V7ܝ��nK����)Z�5Q����^�c�^TuF��U����e�\t
�W@_fw�J�����Ӽ���:����9x��S��������h�����R��a���9���\�ˉ^���.�^��\q�%�[��\�6�Z�cE�@�n��G軈�2��Gvwk䒬�k�o:/@��eCNfr�:��M.�:�P>��][7�}\�u�c�zk�r�м�9@�����l�;��b1�r����\ejII��{U8m���b��H���6n�9��۲�9�|n;�O�F��~�T1:�E{�BF�2X��dEL��u�������N:��5�-��c�S�h���>��S/I����W��\��UJH�KF����jw{�`���"=��d���,�Y7�Ã��r���;������T�Ͼ�u�/?\e�.Hc�طI���X�wr�ajn�-��1�����7`�y�W%fx��.�s��v�gm��''�~�VQ������K�������EU�<�Va��;'b0�.�X����E�,�l�|n=������0����g>�29���t�o�*k���fT+��LTaXLת*��9�V�EeV�-s��{>x=�<p1�u:���}�§�\���r���g������;�6�=t��+�|�[��_��
�þ�djtx������ύ�d��q<2�mǦ{��N�����;b��Ƒ���Xn3�gM�@O݊�TGe<sЕ6�ѫ���"2#��f��|K�_�آY:�����;�$ZC���]��6�<��� ���L�ǳ�YloO_g���ݍB�me 3/,��b�:�w���U��`��oT���{f���+8:ؗY�}�*�i��I��ͫ^`iqy��Z3��S�B��]���Β���LS5���n6Ѵ���-ھ[1U���[���rl�"�n�8T�Պ�t��آ�������Ā���CT��~��oŎW�!�ub�˭3W7����W���]Gz�Z����Ct���*��3�u`9�+��V��ߏ����~'v-7G�u{{<����/�ݱ���YE�tE+�*�g�]>�`I{��Θ����_��I�V.鶆�K��:���g|y9Zz_�Ȯ��s� r4��]t0���=�=�%�xuQ��r�(h5s�*� �9�q���i���|j�p��]8���{ـ�M5�w~�����vK�z��e����k�d��N��gG늟2�����K�z)ıQz�:�8��̟x��Y1XϠ�A����V�O�Į9���c>>���S���(�ݵ��}�[������=*��
�P�Œ<��cb�����^:�a+��㽇�5[���^m��SE��hh9�t5@M7�r�H���z#��Un�MF��(���'���*������H1�J�����T��*���]w��:3����㫟]���y��9���)=0*YҒ��&�ڡ�����N����+��Y�W�D�?��in!H���<�+ei�1��{<v��w��'��.$�ܜ넫�V+GP+B5K�i����s��p�z�xaշ���ڷ��{�H8��f���q���Lū�����e��Ff���U�:����N(鿖��>j?q�U�_�QҢ����1��vXkU����nF���6<�c���H	��p��R���s�p������2<�ٺi��������5�P���}q՗����J��xX�q��~ΫD����x��!�Ԕt�
�ƃ61f�ο��/����w�n�E�BQۮ���3���1�R.���b)��W:��]�|g2w�緂-�
���(��K�z|�H�G��T}s>sq�o��m��GT�~��6Ы���UOM�f�M+���+��!.���`����&/��u\�몴��՛>���t�Hœ��a��];:ܦP�9zn{�q��(�������ǒ��C���O�m.��.�&k����q�,���^�e���i�'S��zaV���3ܳ��I~���\כ��(��=@n���E������g�#�������_GxKg}h��Z�H��������l=�j��HYB������G�~����x\�T_�צ���;���N���C�"��~y4�MZWڕ�C�@�noU�r��|��V�+�q����-�-n�n��ΰ�)u�_����H�T2��ݱo[y`�ܞ�pu��o��ő*��,[��v�mP�'m�kz)�f�#`D;f�lP�m�v���=vF�����p�9�^�'��#{ӟS�r�ߏ�\r�a3���"{�ͳG՛7���{��+�$�\Bw�ˑjeI΋(_ѓ�.d	��;TE
:�����ٶqT�j�xy����
�*���2�r|�(O���S�.:����su����^n�{ ^�ݼ�qe�_yΣ��P�vY�W����.xhLT����u�>��F�=�}���vlx)�Ϊ�{�¼X�;��M}����P���;��N��fG���]Q��&��+���~p	^*�����UT?_ޯx¿e=7�t�ʆ'�L\f��D�ِ\f�Z�������۔_aśT0\F��#��!���J���ġ�>��.���닁�徐0Ӿ����N�V"=��bx�c�d�����}���V�ֳ\V~�?B*<��
���ۯ�W(�xT��pc�@e��7�S��F���g����_q��Toҁ���V�ꊚ�{=�^�δ�O�-Lb!�2�����.�[��p�Tc�Qӽ��w�\r3�J�ҟ����\�����͍�����,
�Y�A�=.6�;L�+�q�v���N�5}%uS����岰�B�`�;����/���˷��� {�r:d,����׹b۰�7�+켊�����[K��ʗ[ݾ|+�'�ME[&9���;4�I���]q��ӶX�8�����̅�,PϽ�\�ȹL�D���?F{F����8/�7X}��Ȏy�h�O��U\D\��U��n=2�?FՄ��65�;#w�0�N���Vug�k�n�i_�/~,��L���3�v�����
�<�����k�B�47,GL
]1&�8Ļΰ��5�����i�z�t��G)gҀGbL�TD��\�9u������	^�����A�x���2�n�O2t�T=���\U�t�1�G�����@�y~�@�w}��\�w���z2Z5{�
�)��/I��O�X.ʓ����Ja����kf��k.v7��
�#�E��>�w�� �U��;�������S%3�����nvUq�Hώ�9yШo������,�ey.ԡ5t���g��uATZ�(Tk��q��'>s�S�]��V�Lz�}�ky�!{� k^�gD�;uWp��X![���+��Cu	���IӺ�5W�uGݝ�;��������g�r�����A�t�o�k���FfT+�e1�a3�����Z>�O׍�i�-�w��;o+q��s���8��9p�JWt�p�gorobݩ�nc��ي��8�ʋ��9�,V��]�Y��w�Y|zj�<8b�������=hWNvu��G�N�Y���R�5A�&��wT�9����y��U��.'�(���1u�vY���|�R������T��D����W��{�q=UN��*66����kJ�ǎM}x	�i\;��k�F�G��������������N�
�\��ԩ���q��/Ǆ���=��)��.��崙��~���>��1㋺Z��}�˫.\��WX����q�� b��6P+�0n�o��~���zӇ���Qa�)�W�̢�8y������'UT9���Ǧq��9\mHC/]X�y�I���W>H�t�S�4��mw,�1���b�JT��ٴ���k���R��}�bWp4���o�N}�o�m45�u�����cE�����^QGS�%qT�[>��|]T���U�RK9&߷1u=[/��}�P�#Up�Y%���NV��_����QՒBFܪk�9
�W��n6�v.ޯ;�}VE�Ό�yZ�Β1�[
9�v�;��*,f���u�뾻<�}�vë/�8�)�%Q��ʹ��Ll�e`뉖ΎNx�Od���`H"$��柳w���*���O��G��oZָL�3��j����>������G�u/n�,����7��:�wa�[R�v傓#j&�\�u��: �]��+we�{d�$n÷.���Olm��
!�}�b���ӭ]�z���N���
m�������ՕzU�'�JG7.�Z�?|J����c6r�KH�����yǯmu�/A������pD�R�P1�Jw�2=�W�����xS9��L/k��Z�8���lUOw�_e���Mq��e����Zy`TE�;�.#���������B�u�u�j������^���E�0��C�5
��Yf�;x�8;��rf�WE��ꫨ�焘=�P�K�ż�y�V����}Pu�P�3����N(��?���%G2WL��5޸�4��R��F���>�<�s}gð�,߲�[o�������Ңucj�LuT.>;=o,��C�F�2��m�)ʇ�O����5�{����@�~��~��=ę�/7�8ܔ�����#���p��a��a:�mYumq�~�C�v�J�_������;V�]�7�`5y��g��{�xG=�
�G�'���NEW��T\Ϝ˗�+UB
�����FԬގװ:�ɞ���Eӷq�n�z/Ϩq�$%�Uxp<�xڜ�����'P'O����$���o5���^GY&��];�L�mhg\{��;�F��C9r���VN��4��4��^����v�=ԇCᮖ���W��Bu�q�m�\�Ͳ�;i��z��9u'yx�j�{.�深��2�dlL�����<��'Õ9q+�ȫ�63�]n��ټ�e+w�AY�R絭:�MJ��=�A7u�{��O79n�:�p�wN5�C�^;:�*೏i�d�s^(d���[��-�r*l�%��yN���%�ʕ��)PW:��4 �ܺ9 V�ruۅ����rӬ��.,���`)B� �x���ԔC�ieҁ���ue�o��,��PÀ�v��tKf�}�����ۤ�&�҆�Xz�V��'Nh]����歄x�b��2�d�v~���y�X�9�W�/���t�ͥ&����]�q��8iӗaI�nr��=`1������#n���7���R=�0n�f����RgԜ�M����o' ���1���OA0��v��Y�\ ����ޣP*�x��g�q{4ek�M*�2�i�f��;i��ΕՏ/;�Z�`W..=u��:�� 0k�����ǩ9�ԧ,�\��9�%�f7t�"�'<ӎNՙ������jc��Y�c���&[�&����Q�:���,�[b��z<���W%��ܸ�p�P[=Ɛ�޳Ñ�7r^�',o����.q��e��Cb�1|���<6��3)�wj����3Q�2���ˬbu�ľ��Ʋ����%��˦��,�����3�7��3s�GWZ^&r���6"9����v����DSȎݙ����&���oC+-Ê�;��+��s2�� ^�磔+@���(ϓH��p�	�s��E<�r&g�aj�<W��rV��sE���zU��&����e�7�@3�EІN���mʰ.�;��@i٪�eA&	�T������4g��
�hh�h��;���}v���4�J�r�yjKgz�,=E�z�ӍŹZ���*Д��f�1K�.e�@.�U��t킆4�ر, �������Ç6�ud7���9Ժ��3�1}l�]�4Zb�:ɲ+v��ui=�v��ݜ�e��.��4�MkriҭpVLu�S@917�2+���X7:ݱ+0K�>�"����i����jL��(o��$*���-�1�m�	�zl�}�Rq��V�Ѿt�3��I��!��E��/I�}C�6�����\ު�ASg�Rĩ����2@o*ͳ��wQ�	��u尫j��s�WV��7�&�+��!����仰`�[T�����F��1G��v]�i���{��P-ɭ����`���\�E��,�N��h���"�Vo&���0r�,;�}C�G���0�Y������w�l=�w�]~����.��Jȶ^ep�O情���1��{�\�/37���Q ���(#2����j*՗.	]#Za*Qۈ帛�8��	�p�,J�#��a����q�x��V\(���D$$8�8ΑBI�:AF��S
f�)5� �p��@�@*&��q5����BN%�PP�)��(�EgCP�juB�U��L����Fi�p� �T��q]�4���X	ZE�E�����XZ��N;N�XSB�sX�-\.��YpK@�JD,���G"
��\����@EvkID吔q*L�ɪ�����^'�"�&Er�3�U�[\�T0�� �$�"�e��-N\�Te�P�.�A�8��#�y�V$��p��DTH���}z$������f@1)o9n�L���l�[H�]}��e�g�5�컾�K���6�\�(�hS/T�ӻ�ặ�wx�gWVw�_��<b�g���dw\k��pܦP���N����5t�s���d_�۫�lR��+sN��[{�����W&��-���⇉A�M��Pա�iL�=+��ge[�s���Z�{�~��u��h�p�����uT{�.W�Ǚ�)^u��Z.;�u��]{��__�H�]n�y���zߡ}=X.;�q�-�@o"�G�Y1辕�ף*T]n�7� zF������Z-��o����O֮��Nn��5}$od���˕v�|J�]"���e�f�7חȸ�5�c\mm�|\�=i�+y�+�T�s��P���Hb�S�g�b/Ն�Y���-#n G0�	~5���w��W��L�.} v��\��T����\o����ڀ�g����gau�w����VQ���и�N�l/#�T*�e�L\vS��䜀鞠$�#[��n����;V̵D����Tw�2�;���k�uq��q�P�uq|��;t�۫o���}�~���h����n>. ���7���Uz��+0��Kÿj�j2�c�����`��Z�3󊌷ّ4�h�������� �%����^@s�.R ���Σn�D�ߊBc������@�5w@�����Nُ��&���h�w5�V���*7�� �>���lbڮNv�vuթ$�67����m��rU��5W� �����owp��MkRqS�B�}�����v5�94t�ˡ�.^�<>��׍R{�=�L��d�f۽�.������e�����{f|ȸ{LN����)�M����9r��q+h�zr���w�p���Kz�w���1M�iP2��@LW:�#�ʘ�>׹q7�.t��:plD���fV�����{:������:}d����1M��5T�u.r�дv!?m��϶�N�G}�7@��\�!ѹ���i��V�����(x�G}2��l�[����k�yn�sڳ���^�5Y��^�p��u�c���;��.��d\���F�2�?}�a#:�x[�ޫz�}jp�'v������\D�pB�|�y:4�I@,؞������<����<c1�bй�7|���Ƹ�6�6�K�iۤDʔW�����Y;�42��끱�^ڒ�h�Fd=[�NVLoy�p�{�,��/�'��ݻc�vT�$$t����$���;;����w_�nhS�X\W�_�ݨW���r�ģ�t��R2�R����'��I�a��x�����knɊ
��q)Ȍ䐗�j�r����O�rsj��� tpa�R
&6u<�9/'oT]Ϡ�Un��}.c�r�(��ηq_s�7���<Fns�R�=�e��wn�t�I��ur�MwgW��y)�ӝ�˹�5j�5��e���K�Ыn��z�X��?�R��V2/*~w���*{@L���:�Um���zn���|z�4��ٽN�v�����V���☝�^&'�[YF����({�%��ɮ5�=2��~���N�^{=��^1W.:� W�= Z�juQ};꫸Y�&[��Q�aum!��Fw�a�;���o��ݴ#�6Ϗ�i�o�R7
^X��D�~���~9�ʅ{)ɾ����Qsm���Y����|L��qn���t�i�`~*����E��V�����G�O=�a������{���a��gѴ��gMb r��3�+d�q�;�}��)h��+�U���3}ީ���mb�Z���Ɩ;�b��n4�&:���`j��=�r�iF�R���3\�}|/+=�a��~s�,�OO�H�Ε@^Dzk
�;g�$� �������s�h�E�]�W�[�s���fy�����x�Ζ���}}�����U_�zkC�2�Nϰ�Hs6׽>�^���n��5���Yhh��ý��)Rl#�j<D{�p��y��/�/~}�P)禽*�,�b.�+��e�.�:���j��H-�P�L��BT�*�/�-MIK�"��}��ܳ�����<�T�qD웳���i�a����@�O]�f�����ه6[����d�LI �Vu�lc�vq��`�5d�[Ɩ��z�3�^̱���2�[�v�_W�ꐎ��D'���=�}O� �5u�߂�����U�pة��G7=�P�Uv[%����鸉^vǣ�(��[D+/�oH9G������[����5���<�d�s�W�r��7���|��ťǭ�ў)Ө[/�aU_LX���b�ڗT|�tKf�2R�g�R0�����f��JQ{Z̽:/��*q1;��?^f��n�{owOms#޺W3��G<1-�&'�ܪ��+��}���=��ҁ5�y���H���}y�1O�ՠ�$��?f\`�T�����jo&@��	���Ml*�~�T,n�ـ��F
وl��o���xe��L9�M`�>o,	���]TQ�f���!���S��N���W����#�@vs�L*�vl�ܝ ���Y@;�s�tf���WO^�S�λ47G\a������X5��q��3Y/	�QPu�.��Qs	��7�?��m�Q*�����Ӆ��/����ɞ�"݇��z���w���X�{���ΐ��s��Sδ�L�P8P����go���W�;i��\[�μn�wk��oU��\�\KMf�s.,!8���x���t���z�o^� �^K�:�Q�'���r�u;O��^qݽ�����jc��Ţt�m�9�z�l���͛�ZO0�yRoN����ht�sfP'|n%H����O�������o%M��s��w�~���V+��ǯAyy<�*���דc���?�%�gǲ��_z���<��)���vș�k<�� ���IW�Ͼ�OOz9���C����t�ĺ�����zr�U^{w�X�E������5*_����({"5��v+�]m���'�����5��R
|<=��۫����O�Wa����M ��2�3�b�.�F�	\k��pܦV��/��ҽ��OnY��硁ѹ��Vv�׽|��_�ԇO���z�����eq~��Q9\��{����;GoC�1�`&}ۃ��T�8�~˽1ޅ�Ҟ��u�W+���͔���.9up��S�yl�{�hy�m����Np��BS*�u�����qu�]�>�L#�%������V����hi�5�y�ǡ�5|d.�$�n���w}��-�򨼔��z�oEj�w���CF��څs��E΃ܝ��[�\�S*HϹ�e�&'��=�^CE�I?I{�ה`O��TF��3i:k�	�s{�!`N1�l�]��mG4�֪nK8�Cm!πY�Ꟗ"Ϗ��Ϯ4S��5�ܕ=5�4\s�(�J\��l�b�ݶ��3����ɜB3���&���X� �]�J��z�q[kWCwً�q��������q� +9���w9U���L�9��V�1Iݙ �}y<u`#j���U�t0..n���I]=���)zw��zA��]1}.�s�S�?uosG��Ϩ�T��f�ޮ�����d�_C���]7%{/a���ᨼ�����:��C:C�5�q�q�S!D���h{X���uc{>n ���k��D�G���~���-��ON���� �O��zӎ��2������xӰ�YTQ哛�uC��I��q�����g��{&|i�P����qG�w�T᩹��c�lzϙi�GϤ��69�jx�gðܭ�<�<��{7;W*}��-�nw(���q��Λ�*Tr�&"�י�T����ˉ�ys�ᬢ7HKG���UKnw/6h�b��֞ҭ,�S?!�SJ�s|�e<�R��ȆsMD&��]�ȝ���N�ѵ۫z�E�S��}-��+*�=��P�L�>%�XHY��}�̼Tc�8���0н�4:�_�K��ؗ�M}:¹=��nO�S�w�U�x�zg��L��ѵa"�*�w��v������{��l�+,-vo1�>�֪i����dttUN��V���|�Ɩ̤��W	�`YK��i�3�ݓ�}o�n�mNf��s�y��������/��W��}:�����b�8-�_n���E$�q�9a���LaS������Iȅ�r:׫�ӡ\o���қU(�5���@U��z�GR�ȡB�o��M�!���*��;�.;�{��X�׶Ƌ�~v��"z�*��Jn�l�QF�w��1�ӝ�^������s=^��\k�ܨWλ���:Z>��pT?Z�=�:*0���(ޔ���3��)���J9nq�~��+*�\�X����K�Q{��i��_���N��z�^��ٻ^2��Z�:V�&��N�D�7��ﾬ�2�W���S�s���;kC''�3��T�I�2'�oD�Um��u�wo?o�蚷4��q�%�f�6LlR��7�)zw��������ލձ]X�v����yۊ�͗r������=���S%���Uw2|L-�u�k�°���-�u��]U/?l�B��1�6y9�)�ϔ�5�܋U,vlT׃��̨U7�Fdg	�ʷ�g���m��s�.,�&j2�q���3z���΀�>��U��Q�§�,,7s����T�O]�k���y����\zr�oD����Ӹw�5����/���6�Y���\9�Ŵ�VǫL�����j`�ť�Bm.�wRo:njwhG�[������o]��GB�펭">�wDѣ����w6t�/ِӥ)��R�J�){Ҋ�:sEZ\r����V��֡hG�n�^d�gQc9��{�(V[}������qk���ٿt�$*;VF�L[ |�wq��c�:�2�m��d��|r1H�7P�k�/���%m�ݧ��O��^7(e粶�f��s���0��(�;���><��D,��i ?eA=!�ɶr�k�5�w�p��X6�ז��m�1k0R�R����F˾��UZY�ʿ����PᏪ�F\yM�o9~T_���>��Q��y�ϻ���ۛ���z�uq�{��U�>���/�]SW��U�I�,k:K�S�nS+�ݱ����մQ�}���H��,j�^���
��o��9:��� �����jn#�YL�5z�^��6��Y\r5��r�1}U�(�O��pw"��օ���
�G���U#ǥ�G��=�V��{�t-OK�G��;�	Q3Δ������>�q�G+d�g�X�쿩�1���`����<5�,��+g�LZ5L��{��*2�����O����G_�ލ�,�+���>>��Ae��^����o�P~�Ɋ���h��/�r�<�y����]h=�;���By����?��b@w�V�*T��0�;bͯ�v!���E�p�ոm�X��˕	��6zeuܙ)6d�T���g��v6
�R���n���j�?^{��G}c<����_��n��	T%�r�vb�`�XA#!n񊻈m_*��X�{��:��:4Ë�]��M�z�Q�A� NG�wݵ����ax��\o�S}��'�"��r�z��j�>Zվ�	�#�N�����v�2)�Z����� +=BaTGs�f㓠|�(az����:3O@����]u������_^�h�Ut�z3+��/L��(a���Ρ0���e�z�8j9� ύz�[{i�N�\�nk��q��/�ΕJ:vo�0�������\�3Q����p���A\	�½��P��ӖtΉ�����쿷&�Ow�lƸ,��r�m��}��P��ᕞ_����zrQd�"T�*x�~⎐����D�9�D�|+��<5�V~�A��4X�R��DTϻ�^x��oٻjCQ^���yX �n���^f}���y^5�
�G,�Ӿ��X0���:��r\dǥ������O�u���9�fX�rW*�]S���O�c��>^�	.����i�fͬӊ��y�߀����zg��ze�ٮ�2�X}nV����4�gdlz��^���)��ڨ
f�u�AOUx��e�C~����6;2ƽ�MA�Y$UaUFç�ZvF�T��y2��9{��u�kOK�J�yk�\�w^���.�I���.�l�U�%_Mzk�(��8�͆*�F����y\�Ϛ�f.Y��c+]��)X�έN'}`gR��w�KA���˾��e�O5���L�ս�W�u{�ݪ���<cɊvQRΪ������3�zR=~�x��>.Jq'ԍ����f��X��Q� ^�v�{g\?F	M�*�G]��^�*/�qt9O�;�W=;�V��f��lh��;��:Ol�Ԫ��M��xd%6rHճ���#ʫӯwS�^Y�^<��%#��T6k�ݨW��ۓz�p+��`��I�T��΋,u���8O|"��X��9ג޿CVy�H\�=�W��W���{�\o�S.O�u�\'�"�����F�nm��j��o�7\��Ee4��мR��We����t%ϧ��E��V��=�~]ݞy��}@T,���Wګ�Y�¯����p:߶�ʎ�%}��]=`������W��Gt[��A��Mp�PCVMu�~��ۨ���!^�����,c\��oV㑷�{f���޶=	UE�d�*�����>Y632�lϸ�Ľ�x}�{6���~��;�aثKFg�ӽ�?R�ck��鄦|�؅����s�8�
�h��.��3ù�"��,]C^�1n�� �4qg4:Oo2��mhS������a����[XN!}2j�I�
���y�]�-\Y4���N��0�G멸��]͸�!�
X2Se�L�[�=�{`ܱ�a��M����]"$ԕ�3x��&�\x��8�W`�y+x��Z�Xq��I2�vx�>t��ᕹݴLnkn���R����s��ܬ�}�������1�5�E΄����j�ׇ��V�O���`ˤN�w$�[ub���m�庫��&�f�;����q*�����	�T4����1�a�(1�S��`���P�Iۣ'@N��Ֆ��׎���#w���=nTz6mxq��Q�n�6	p�ɩ`t2_U�wO���Eъ�<GJ�#3�C��.HU�wY1tI����0���ٝԈ����{����cH�*b^��W��]ë(g7��'&�1Hv<�Q�sF�j�%�n�f��/:(�>_IhN����
�֓�
�=}sr
�@q'�e>�<�T����K���W��@���N<UK��<K�1:���X�M�=+
�������
�ޕ�����sH1R�PF�6+J�i�QV�9vÎ��(|���5��5V����n���o$��Y{����E
�[�s7�{������qlTc<�([t�L�}T֗w��ΣnݕEu�`K��V��|dS��=x0�y[1�D�� �u:nn�g]��������@	sV2/t�.U����;������U����!v�	�!�����%����B)����"w����K�ϫR�ܫ��;M�2g�=Y�R|�
��N�O��EF��9�[�5{�呹ˠSl���(ӭ�b}�&㋱`�έݛ��WDJ�2�[��{}�Y��.y�u[p���r�\&��f�T�De�OVŦ�Y;���w;q&n�U-S���c
Tl�.�|vd�:��|�N�|�5wø����rCa���ߖDɛmVdk�\;��B�I��q��.�3�y���	r�-ժ�������v���+���RN�9sq�v����fLM�͗��R2�.�*�0�HT�5������Y��J�����l2_`�8���Qu��;�j�n�:��yR����N�i��aΧL�m�T��ŖI�PŔ��b�r�$8��Ŋ�)!�:��OI���r�n��^Ejs(���_JmZK5���.��q����X4����I;@g�.b�͢�ʔ�d���䏹mu.|9���e���MC�^�� E��*$=��;�9[W]z��3��vu濹Kt��(?���,�C����J�ԕ�ի0k��A��`��ӭڥ��Ժ�"q
rPN�}��sj
�M42�Ƒz�~y��EQ��H֒d�.(,*��U�(����őH�%�Vp��s��QUS�ǃ�4����*�$�Ċ��
.JВ��UDD�&R�6��*�TAh��"!g.��h*�j˪�qLUD�B��
+�Ќ�A-#��MPBH�-�qaEWMS��E���%PЫP�Zդ]���s�U�*��9!D,�(5jg.r�E�RX�A�(�PY�J�8ɑ.K�#�TB����Q*���\�	�QXVZ�%sD���*�D�:uYr�0�B��r�-��T*�D�!�P�NU�r֢�J��r���0��d��(�3.D�QL� ��*d�T�B�#��*dQUPV��"�ʚ�p�gB""�DFj4SC�Ar��
LeA%�E]*��u����9ׇ���+n��)��ehLc4e��Ӂ���s���+v,�RN�o6e�Z����_.ʰ"��%Z������=����B���ǧӘTgB��RE{��#�5W1��k�OĬ�)��������v���%��J��PO֞�q�n)���!�ƫ�]+��=nsH�yU9�ze����v�^�l�1�{��.N������W���q�Gľ+	��[XMCd^�v)��n�v.;O�����'��|����n��I�*n!��s�(\zg�����S�$]Ƿ�r<FE���J���5W���4{-����3
w�xr���_�˄�A熃�yz����"j	�|yVA����E��<9�k�B��]�h,vt|���r��}�.�YJk�� 9J��\/�E~�۽�{��C�M����JU{�\j�*9�+	����pS��@?K��#,���۔+R��=�PT/���,���BwN˙�Ub�!���|j�j�����_���ʭ�*���]�� 8~�K�i� h^����j�χ��Ð{�Z��t�{7<�&&�$L�18�����e���g�'"�Ӓ��%q�s���i?k�eg��ax_��51���
�d=����vәj�o�Z%X�t��@V��N��+�����Փ��ј�M��m=U���k,�L���ZB7��6AԠ=Z-X��Bxg<��} �h��Xw��u�C���p�|�d:�m�����0Ҧk0��ꎧNOnp*�.�ް8��ua%v~�:��Zn=��79'�u|��V������?�m�ܕ�xMy����;�?^���뫬׳%����C�(Vs�f㓠z�gЧ(
�~wBn������ݩ@sf���k�W~�7�3�+��qP����Ι,�'@6�]�q�#^	�5�~i��h����I�҃��hg�x]ڱ���<S���r����Zg�����U�zǶq��d�_w�ۯ���u����^���*�c=��U�zpV�#ޔ�R�����=0#[��T^F{G�_p����[�q7�����M��Y�^`HU���a��+�jC�s36�>M��.�wn+ ?��	�c�1z�O���Y���DK��{���G����3�40��s��ۧђ���`u?��!��X�}I��>���,��<;�S��Ïz\`�:��M)�=K��~��5J����x�F�=2�#�ٔ�����R��=�8\�VהQX�C8��;����l����Ӑ;�|l�p+��n<d$�ڽP�Uv���y9znW��WyTȺ~rL�M��fZCF(�(�q�����zC��՝�Ѭ끒��RX��*�YB'�:2�-F��dR������8�זW����F�qS�k���1����9X�x9f{��I��%p�lh˾�P̔�梕��g�[�s)ݮ)�	[oYQ ��^02��:��[���SZ_��v�5�<��Zп�R�8���Zᮽ�l?}
{�R�9oJ��
�<JP��y~�2x��W��3fcIA�	\o�@-�;���4<yW3^�C���)��z��f���.�~���*\C�#j�z(\7L�/}�%�q��o�2��W���	\s'ْ�a�n��~�}���yL �e���A�E� ����4�>��7;�_O�+�a�~��ITLQ�����YpN���0�kX�*;&��RÞSX ��@R�RGU{���W`���e���������B���$��V�į�����s�gc��'M�R��~�+<<���4S���qS�ݗN�ˎ�Y���ܡ������}����(:��
������8��ߣB��'�USwt�V��_k�n8�_���*���?�ٝ��ۓ�_��q�}(N�;H���UN��^����ݷǧ���]f�V�F`^�톿7�_|�k���s)~�b=�*�֒w�O"��@��v[Ѯ�=x����o¸_<5�}.G�\��6e[�]�<O�� �R2/N��T��wi�I�Md���	�\��=}�ϫެȸ�.��PY��|��*>׍vF��o�%cIr^7�6=v���74�bf�MkA-x��J�އ���&$s�k�;S���u�ѽ��r+�@� z+�y��G*z{���H߹��B�O;CJ����ѿ񺕤ʿN%��:����q�SxTF�fX��]1\��u�[��7	��O�;�7'M�Լ��g4ҏO)�㕃^�~��u�;�L☿L�S�L������C)���L�gzz�Q���ٖ�We덼TQ���G��৪����/�%q}�c�'�c{�զ!���my��,�C�4���7��u��q�(��1N�*@Y�w�T\�*�y����yu[����_hy˫���S�h�}�����1������!)�/)@}�R<+�Y@A�4Ǹr�/u��s�a�{Q΢�t�K��q�N����j�Zt��`!)$j��Y�#Y�������{NG�J�~>�{�{&=���+����u��N�hk.�Z�RG���.�r���ѧ�n>e�LO3���%�G�>>��%x��n1P���Q�)�%Ϥ��4[OYB��<��^�]�_�)���)��w"+(��=��"�悇��T*��]1�0t�\�f��C��f�{
��z�OϑX5�g8��K{���s^��J���oS	��Ci�e������R`�u��wgN��᭧�
鯩J�z@W-_%Z��=�uݷ�+��;�6��&S�o��Uqɋl��Ο8���Y��l�]zsO���8w*�
��4��S�T������O�#(��,��3�_�k(l�l]�����;芫�Y���*�,l���u{LbT׃��	����a���� ���o�d7=��e@��]D����U뇞���
��S�؎�㑷�]�m���K���T;�b�"�S'n�ϔ�X|	�.������'S4�j}'�%^N���w�y�����{H�Ld+��!)bt�e�a��W�@�>Ί+v�[?�L�N�]�?b�-��?,��/
��T�T�:�#ܩ���׹q0����gA�.,ןl�{�����B�����V��XU��s�)�A��׺�9t\���Q9w�*�w�p�y�������3��z7��^�JG���S�=��P�L�7��z6d-ay��|s��?x�5y���r���n����C{g�w��R*M��]�W=��g����^W��no7�v��=oj��qZ����h����^ZF��n�{�"T�*�.��@O�w|���Z�gWQ��)|o�<k�B��Wq���_{(`��lx�T��2JR+��Cf��s��F�#�8T3ٛx/iE��kƸ���N�h�[�dJ`ϣ�l�ۂ��!�q�+���C06q|��q΂ E�2"�Q���P����0/�Mu&��u��m	�Zk����J�1�[���{u1T��yݶ{;�>Vt�������T}rە^ʅƢ�*���#��KE��ݿ?1�K}����:�.�U�I�2�F� &si�*hW�5���|j�j�zw��%��^���w�4r�׷�Ӽa��r���xl%�d��[9D{-W���=�= ������݊�衴�u��픹�TÈͥ|T�8j��'Vd�l�|�'��EW���[YF�K��R&/!�ݩ��������r�[�'	�P�i�t�B��9?\	4���Uӓ5P��ea0�ҽ���yw���-�;���\Y�v�6�`��(Tg:6o��yu]�g"��:�4߮Grj�z��[�W�B:s1��v'��vTm��&��f��3Q�t�t�g~���Ӫ��eXZ���ɍ��j�^:��h�Ϗ��4�r�->�����2�+��d�A��� '5�<��>D���7_�R��ۯ���\Bܳ�qΌ��l��C��3ѓ�W�	��R1΄GR�C��M�n3lD�ñ�Q�+fd�L�?Fk?��k�1����|���!���G��� b�
�-���Cc�����M��M$0�r����Zi-K2��٥���5�'�]�:V���{�ifI]Xhx5�$z]�Tw���y��X��q���W�[��E���fj�Y�%3]!z���!ң�_N�O�0����.ޫ��̵��a��ɜk��LخT�jH!M2���o���ww�k�BQ���.�7϶���`���ηI[��?d)�{;���Ǡ���˶�œӼ��]�Ԅ2�Պ�]i�ȷX5�R5���ތB��U>�����z{й�n��8��ǌ��3���U?�ej�����g˺���{��s�m�$����{�)�}H��E;D������_�Y�������`n��)��c/2Z�ɕ�T�y�Kz��x'�����Y���s�o�)y�]ŉ��<6�������ѝ���]/H����-��'*u`vS���	H��f�;���L�6. �f��Ͻ�cQ����1PO���<��Sp�N���	�5�KF�bx-�e��Oǐ�8}j$��
F���/VK�>��T9�(\�n��{�ހ��z$U�F�_1M�&@�x5C�Ou�����θ��Nf�pP�η����f��ٮ#��3�����`TZ� �y�s�>�N��ݼ��gn�e�f���!�NI���>�W�H0��=����VP�߽��~������Ih�a��|��Y?^ey��A����ֱ�}*�7 ��ϑ��rkW�k�Ҩ���T��H jq�=K�
�Yk�n�ސ���_?��H��)vÑ5�W�NwGm�e�[E8u��}�3�$��Uv�>���o�����x=*��)���
N��:�
�z칇�x?Wl�y�B�vl��[��M�u��IEQ��?�ٝ��ۓ�]�p~�k�rP[�P�so������MU�{�iE��#3���Ϲ�ό��� s�_k��_����=f��cţg�/	�?4�9t�������V��� {���ک�����e���;����ⶠٟ{]D��7=����P��~�q��:vq<�i�2��@W)�g9S�ގp������a���W�s����&�7��h���D�V�W�V�r�����ᮀ��ʹYQ�jx��������jS1��v�OX~=��Cxg��w�W���g����t�F�~-���gO�$�%<�D���������s�;��ʔw������u�Qs�"����\_�lwz�^H�˟yC��t>�=o���]P��˖a�tj-R�9dEU����N]��8]��F%�&�t�пVv���|�5W�����-�ǒG�'o���:�T+�!)�.z�}�t<7��ў�`�2�g�n]��Y�wZ�NCqs��]�ջ�&NdAgWEC�yPc4�p�X(U��j��(h�ٶ�vs����7W�Z�7O>-8���n�勻��Z�X��ѷHz��ƅ�Y�b��u�O�[���wͧ�J	YR�\6P:븰w��~��>�p��eBꋭ҅Ĺ�7��k���h�yn�2����At���=�lGh�
3��}j=���K�M�Wo�ı��Bf�B9-�.��'dhW��\���#-Z�'uqع3�~{$?m,\d��;�@1*u����A+Ƶ�C��*��˓�w!.��Y���(
q�.E_+�$_H�5<�lVQ�)�4/�R��B�<8 {/��<U�/

u���*�6�����9A��*����}@s�t@�����T/def���߱NS��I���X���>R�ssD�Q�����}6�h'�ˀMC@OY)���C��՘a���\�%��l^��ά���k)+/:��/2vӪ�>���:\�>]����2���z��4�a{��eV��ٸ�@�,%3�GJ�bx�7%�aDFR�j;uۃ�v{}~�,~,�5�����u����ӫ<��=��oP�m�ʣ4�5���׹Ѫ�s��ۇs�%�e�)�H�;.'�;�T��=5�_�q�^)���yz��"���$� j
��Tf�=��,B&L|C;�����%;^�/��#�t#��D����H˄��ld���	���:�s�އ�KR�Xh��j���C���a��{,�-�L�k���w�r.s�E�CE���v�CڲڣݙY[�����/lM���ߚ��?����7O;ѹ���7'	H�%�`=t�@-ծ��ZY�-/�|���:�e�\B�^GoJ���^���<���ZO_T{�<c���<�|��;��Y@k�Q�LUmh'!k����^���"�e{4=��^�ަ�d[�:�z�!����7Ɋ�mT����vm��Ln�Ε��8P{�}y-����|��{�$nz���t���w*x��q�#�4M�c5Wwb7rϧ@ݟDS��Wp*.y9U�ʅƾ�ʅ|���:Z/A�e�K�b�37з���t�q�[���.�d�ѳ�u�S�TЯ@(k/ђ��׻P�:��;���d��t[�b������>&�W�]4ꔞ�-����}�FU��>���(?j!��?^���yo{�Bs>����L��!9�	�'-M9 \u	\n��{�����]t�O_��w��t|�o�	C��/��b\�8��p,f�T*���*��fr����ɬ�:�׹kD�8�Y&��ղ��GP�+9ѳ|� �Ц�c(�@�n�O� ur�;G~	[ջ�np��#��h�2�N�KWC�DƼ Q��3�*]�YȖ�ʙ ��H����"P��t�)�>�f;��v�hJ9���b��{z�kR�;Q�s�B��ŻM�]���Ы��F��
vY��U�`�y��LI#��1�v<7��Jr&;Z�Cu�j�K��ܽJ���7͝�+�I+iTzI�/�X��_�V�9�'O��X���^q�qҠur�Բ�%y}ӧ�Y�k՗R\�����>	�͈�J�f2��\\E���M�tsg+��v?��9�S��.�E<q�>�1lgd�Ũ�B!���/����_۸�5�Lux�k�0V)b��hɨ������֝�n-�s�"Y��}z�A���Klgf��P妭j�gR|��ټ�S*��3@0r5ٝd����`A�����zIm풔PuC+��vUҜa��(1�
��g�&��b��"�v��T���>��ĭP�֍k1K�	��to������u>6�ن�����D+�F�IT�χ�7�qt!��ڝ��%%�L]gp	[J�A��yY}��;�\�X��wӪ�3�m�ϊ;�\ohoP];4�c��,P�Y�ڸ>xk)�K���w(�P��@6�����m�p���4MF+��)�;eb�S���{��Yr�-��O�ç	��eV�.f�Q�����jƾөw�q�h��ǵ�.���K)��0�C��S�Xt�b5�\/Y��f��B�(��p.�wC��
�}�۝b@8����t�M�����t�r��O��a���������og&�,�ߤ;��`�ݩK�ځuԥ
�w�WD)M��F�Ŋ�"�x�˶l`IڵZ��;��/�������'�O�i鹸x��z�)���k�S����#kl��IŽw	��x��_q�.�|Sm���ۓR��k��	���˗���H{25"͸:&��f�(@�l鐣����d�A�<;��z�Kڽ�|9�o;4u6��-��E���;�/;����D�9s�+�X��4f�S��*���t�����yR��^P���J�ۈ�Z��۩�-R����@��k-(]Jŉt�O��L�tֽ�}p0y�V���w(mYj��Ӝ)9�j�������R��94�g�z��v�wQ�m�6�L����Xۯ53��of��3.������>=�Z�s7r�ߘh�^޾j�x��F����CO����j۰z���Q��̶)]b�`�\�ڶ�9&��^����31�Q��7�8��0*:z�m�ۓF�7���x��X-L�;�����⬙}�LC�K�*�Vu�%�~� v��Xµ4������se�i��QR���]M�:3���1k�:@Y��=�x�J����ao��kǸ�K�\E,o)
O���:�T(Ɇz�
t��[O�Z�x9����Wcny��rM��(�5Λ�5'�9�Rє����Q�5yd�:�_�9^YT6��f�yP|�l"vM���MAJ���m�q(/#ި��:v�]�ck-jIP�1�Ȓٽw8�|o�Ԥ+	��Dr�*r�X�qR��B,��r#$�E��ב�G��NG�<�<\�I�$�t�Q�K�P�L�j�QZ���UQDUS�$x�܂����sJ��G*�"�4�����]�nW*�+��Y�
�$�4�G
�W%Z�$�&�sP��("*��rL"�'9�t.U�q$�3s��,[��*��Uʪ(�Z�8p����+ǜ�����H�Y�A ��ȍKs�w"+f�"��+4�Tr�
��Z'qXQ��d*�Y���Y㋄��+�$T�ԉaI��*��¨�VU�%B�
���R�R�UDW44
'E0�*�EQ��+0��(<y�DI�GbĪ+�#�PAY�,9��QETDE����<`Q�(���J�(�DUG.W"�Ȩ�(�I.��q[(��0�#��r�ך;{kx��/!�x������Ak�����QL��:UX�'fŚ��W�+��}ڷmnmNm���K�k/���i��۹鑷>J���0ߐ�m�x���o�,&j#*5������2�ԝފ�3ڰ�-�s������|O�YLw���*��l�A���(�P��5��S����W@3w�r�}���{��㲩�̄�X���~���o�S�x����1H�7�+���+ݎ�ί��
p:��遍S�>�^�˅�}:aX;�Ά�*�=�8Pϼ�l���L�;�'�UZJ;|��qꑘ�3���b}���\_����?c`r�A��3)�K�(����$ޙH�yH�jB�hg�˭3Yiގ����o	�[s}>Q�}3�!�Q~γt����᝝o��ɨ�/.�8�F�2�3���K��L��v���ñxgi;���xj+ۘ]��a�d����U��72s�z�\j�´�{����YR.ŏ	טڽwe�/q�G��ʴw���?R�9eT��U�T\�&���j-�m��\�G��ث��G*��#��\-���;w��tP
G�d��G�B^�{ϿcT���B��9����N�,�~��,�Xt���c�d��g@R���o4ӺT`���cȄ�x�_C8ʹ��#�`�Y^�ϭ�����]��Y{rN�60�F��[;�I���Q>饭F 2m�����4�i!JSy9��u'�P���pBU��`N߷{��%ɕ�C����I��ע�\6�B���)��B���+Xs�����q�K�mUz�E�~�q��	a�t�.'%�����<�Č�H�rZ�=m?{Ey���ٗ�^���Xy.�&'��Y��O3��Ƶ�b�&��{�[pπ_&��m� ��/V���{'�;÷o.����<�Q�/�$���YȎ�0��ٳ��K�U���
�o�To����;�
|}@S^��7�E�3R��2�+�:�8P�3�Pu�u
���t#��hW3�r�p�c�o|}0��裦�;]އ�2@�ߺ�*��O�w�U��fx��Ӄ����:į�G	��''���@;��B��圝Nhd��͘�p'|n\�9n���+4�.�E�m3�D��N���Vo
/��M2}����T���^W��W熷IdY�P=yע��+�w`�ޜ���O�]f�H�6�(j�+9W��|��Z�^��e�dk�s��C+i͑��j�q���8���zU/>�e¸�L㛌*#q�,e�&+�r.�-�f�CGg���E����/�#D8XR��b�)^�X�.\����oT��2�o��0mf��8w/4�j����Q�Xd���u�dyP�O���:�W�C�]Ώ"8{���-)f�ӕ:���䌛=�{Gx��|�_F[u�=W'M�f�;���.Ӝ��S��;h���BAO�����T{��_��S��}�BW���浱ٸ������{��P��/�s�o��ˆ���{@R7
�H)��=�*"��CĮ.�r����-03��:�[���Nqb���O����{���QF51.����+��T\� _�jL�9��0�s�lg.�4����/�����¾S���N@�wP�<bR6�\��z=+���x�j;��vO�@Wג�U���҅˝��<�<?Z��t��v�fc� 㨮�3�7�ט���1l�����]�x��W��ʄ�^�B��{mɿ������W)YޯM\�rM���:����@qV�$��r8�^��G��Q�w��_��W�kڇq�\}�Ny^:��N���s��n�ܖ�(|��TZ�rE�U���n��Ȭ�&)Oa����P���o�\�H,�/�*����/\��a���K��E@uϬe�>n�N��a��4�w����=mu�C�sGN���ӌ�̒Ǣ3�;��N���ʦ�?@YpCVMu�/���C�������>A�5�?Q}�k3VW���������t�b����a.������M���7�MϚ z탷k�7_�\�1�x�e�.�D��w]�>ʽCh��t;V���l	(q��MѾ��X�{*�������L��ˮ
�����7N��De-u:�wO�b��� �%��+��Ϊ(��u['��P�6�lTkb��T;G�k����e�(p�ǜ�.F{*:��Xp&rrP�:�1iUc#˩��F?VI�D9��@��&�k}�g�.��� ��%�.@��H��e�\G��N��*9P\�̎����V��w$���]oE���{��K+8�N�_�{�o�O����L��#L���Y0֋�d�֯:�J뎿@�V���pѾ�͕G"���<�}�x���R%�|o��x�3�8�j[_MvO]VW�O����<�̅���B���<���L�J�\e�C�o-�v��N��bW��r#>�{�>q5��'���2ѿ�2�/FՄ��u�p����������p+��tiN��Qӏ�����p�� U�
�s�ߦP\}�k�B��Wq�����i�Lo�L�p��qɵṾ~ڼ�:���6VRt�Q�Ⲡz.y9U��g��]��l�-[���s���;s���}��a���hze:+�$���y�uC/�Ub�!���|ova)���
�����Y벮��,�Ps!X��H�R8�W77%i�X��\��9����<4��o�������=�	��3E�����/�#�]{̼��L>��m��.����y�55�F����	�U���2��?½ն���g��+=�ܗ#�as'�����f������r�x~o�x�e�
��T���%�q��o�,��6͌������A��;��=�_�����g�ҩ��D':�y����T����+�0t<گ_���7��1�7o�5E�{e�@�=],�;���t�|�pO� R�juQ}:F>�،
��ǽ�6���Fk�a0����8[����o:6S 7Ц�y�GNPD�t��a\o���.e��З�\����9�L=�e989�T&k���Ϊ,�'@%peǺ�J�]�q���z-��ׅO��SO��i�@+Fg�gW��?�� ڄ�o�!��EF5�S�2����+a�>��d��O,�޹����|�m��d�q��Xq�;�F�9^�G}5�n�u�e�]z����>ʹ�?9��Oњ����1]��Lr<s�J��zk
<�Ӳ*mα�t����H� {�ԅ�L5�Y�&T��������<ay	Xv\��^���k������\G����3~r+ڐ�_���_.��g���Yhh�ϴW�z��F���nRy�q"!zV~�+�.V*��å[`���4&�#�9�*s��/&�.Ƹn�"�~u�h�ߒ��v>��}��4�	�*�3@�C���w��l5ө�����g0O9���+���g
��a�Վ�)�L���ڽ�=��hʗ>�S�������L����A^귇��V�-�ᕀ��t99n�˯woT�4-��[�i �*��x��p-�#��!'>�^�W����{�qS�M����W�YÈ��g��}+����(����Vn!ʠ���eʫ���,Mǧ��c�"�yu�R�Σ��]��+�����Ӑ��o�У�Ic�*|)q��H/�wC��f�\|��)�;[̝ŗ�k=�
���+���E�'\T�$f���E嚅��Gd*�.����ְM���y�A�>�w�z}���:wJ�ѵ��Yր��"b��>�>"�fͻ����o�9�v���]́����1Kg<r	L�z����d�*Xs�k �\�(��UV����㷌	{�����=��D:���5V�į��0��ٲ�A:�Ev��ݷ���Y@k(�ɜk�d�}7(eǲ�+��3_d�&MF� g�|+�����v<r��^�q羪91z�Q�|�?D#�~��(�
��?�&d��R��w����@�uG��ex;� �2�oxec�1�'�����K)+�q�&���J��_3H��h�uӖK�Z�s-�wEB�8�2��&�J�z�}Ó7sz��#����}W��&����A�qV��_`j�,��\�6'\�Y�c-��\+W<�*�۽z�p�@�J���:�^Tʛ��M�����5�}'�r���<݃�h]ז̿G?λ��H����a��e��t� Ws�`{�T��s`��N��xkt����7��e�3���Uy�>q+n����oʺ��1��L��E{��3�^�֯�T�T�՘��9�ë�	�%���Vw��=��+[KY��c���=��ٖ2��ʹJ�6�^ſ{a_w(�����G�����E�X0�?"p'���X��9HuY��\��{~;��a!�QA~����py����s���O�Y���H�*� ���x��=r���3�6g����g�K�u��6���y)�u�|��7��u¿}�A�LS���Eu�
��NQ��0��`�xVV�u��͝��:�B�up���|w�=�2�;~�=��*�`!)�fJ� lukU��z���e���*ܮ.�P���J���!A���#�!z��*��n��^��W}�������#T��d{>�42�����\s�ʄ�E��+��h�B�Z=�s$S){�{b�3*$�������.�+3�P缗Q����4��or�WZ	�-�/z򅴛�oq"ԭ�n^ӒBL߳Co�m��L�$Z��luJ���Wˤ@ʻ�(E_.��ru^v�H�d�3�4���n�NkK���G<���+��;�xY��5r*/��H���P���G} �:�x�0� ��Q��C����&jV^��TQ=���5�~����*�su��VQ�a������l�y�(Ɩ�}y[y�%.h��1�])��t�'��Ϩ	��ӒH/����{+0�� ڳF*+6�9��V�w�%�y(m^���%��7�?F'!��2.�m��vMu�r��P�x6yM8�~G���i�k���앇u΃5�RW]��gUF)d��uC�.{Y��sw�x�m^J�&�Y~�z�SOkƓ�a߿�R vS�1L�"֫b���ǻ3]^Cj.�}ç^�ݼGs2��$���U�mV�Z4���K��������U����wg8E��>��z�_h��q��ZG�k���Oњ�O�9���?V+}��e�K5�_�q�^)�n�y��[�d��|җ�i�e@��u>R��Y�4���<�����NKd��=����=e�{ϸ��+���n�����t���zW�fB��b�}�\˧/IW�Q�1ޅ�T�©�>U�����2�OĪ�f=趋��Jӭ7��_�ݝ�M�̍�q[��\��Q�2{hT��=����R��{��-���g��8���@%�{췻�#��Q��ٌn��v2��FN�2�S��"��*�B�ssUڔ���*�q��U-�l ���6t��*σ���#q�9�6�$u9����4{"S
�z�!GK��
נ��s��x���Z:���?] 9��z�=�*��>%ǵ��\j��qD���{hh�fiv�����)�n;�r�����s�-��"ʪ��}I�Y0��za.u�I�yI�"��<�oo��~+5��y[�=��V=u!#�#��Gg�*�]�(k/㘙������N�+�R&|n�ʟ.�	��b7�_��p�y�V������b��2��6��}��C^����5���+���*Y���@V�=Qiՙ tŘ:�)D�d�Ũ��5��/z���l������K�\o��N}�p�O= TZ�7��j�e=�2Mwgk�grq�U�v{�&}n�MF���!���J��g�М�������p0��2�K��}��jzqK��~j�g�r�!��0i7������°���L�u�!y�E��G�(l癊M���͘�eL�Î���`/��x6�v8%o�qg��=�[��eիq]l�ɓXP�O��/�
6v�I슚��jm�Fؔ4~��s�O�4�g<|x3�=j,]�q���(7+�YՓ*_Vwm��H��ջi:�tQ�ےq�9��Z�"m=�n!����*�=�닩lg��(���#�Ge���;S�m�ݽ�ui׳�ypmi��Ğ��{�i����p8�(���>:�'|v%���u��{��мpO��B*{<��@Ɏ��{��B�_�?:w�`{���;��f����1F�� Y�-�|@���˩BnX�w�e���H�~r��b�1_�R\m r�bR��c^K�]��}��
�	W�?~Q��B���?���wƽ�L_ޙ�n<�WR��w��ҙ�n�����4*���u�-F<�w�л�{�x%�eK�>��\x
���q�<*Ա���A\F�~6ܦWF�{��2���w������^�;�ݓ(�c�)YT�[>����P=���>�Do�\'��ҫ��{�A�y���N�Ұ�^.zձ��x潢�r����r�����,NWv�:���s=x�ޗ��:�m�]�-h�z^��۸w���g�o�@-�E;�仴�%��cʎ���u��#A���ײP��ж#����"�ѓ>q
��EBt���F�D/VJ��"�PW�n;6�
��őR���Pı׻Lю�;���}������;8�� ����@�6��0�6����@�6�� lcm��co����������6�� 61��� ������6߀�m�co� ����p�6�� lcm��co��������`�m�����d�Md'�
d�~�Ad����v������U���[�Ak*�a�P�҆��5�6�� wQM�-h
���U!mTM��[c��G%( 
� ĕ4�͍����Gp;�{� ��e�VbE�vCs�F�n�6���N]�A2F^y�E����w�� ��齬��ѡ��[J�,m|��ӺΈ���1w,r��s�gt6��K��ʋ3��9��)����}�_k4(�J5v�m�{�[n��C����h���N�'6�- ς^ڞ�:[n��֑%�WO������r�3*�n��[v暶eJ�w���U{VQ�9n��ҕ�n�]s[�IN��Wl��Rf�9מ����pww*2Ü�k�b�vb�B�a�9��g�/��p�l��Ak,��Vm�����1��|u�;m�\��vj���k4�����qݴ��\�u����>;�Pwn�
�wZm6�vr%��B:�(@      S �J���0   CF��S�0���  4     U?ɐIU�LL	� �0 5<!4����`=P�  �L$�I)%M��      �	��jz C##M�t��J�xZޜ�9Ʊ��`���}<���QC���iV誂/�
�����P.!
�7�
?�?��4���d�1���@�*.PP#Q6�􈢁�P�E.1K�D�m -DP3�ݮ��n�=^�y���QA@ڀ����h�$��-�Y�>�;�x.�?�T�p#��lB���ĈQ���B	(S0�Ӆ��) ȁ�ҁm�a�$HF�Z*x�#�\�U@i(�H��E�������_ĦP�Ah�]&"I Q�B-�P��q�,�	jx�ML*BѐNRP��.\M��I4#<0�T�Jl�� 2�E�$'��9���j��<����Pf[�z���B�\J�nAv�=.�cE�R���۫��R� s!0;Q����iߥ!�ڥ>�5�LwB*�{,\�D�[��*SS�U$�M��ojT���Y&1V�B�-�([�#W���Y�p�*u�tXGe�R�-�7x�(�X�ê�K���Bb����c�W��v��B&6�D7w:QÔ���ޓ�=�����U�o�]�*��s��]��k���$LL>�U\nYc��]�l�]0�k�5��V@�vJ�X�$Vtڹ{Y��sA̭�ԛj�sAF-˴(��*��f�-�7`{n�"j�$ڢ�٣��lY��ZĬ��3f��Ol�$�����V��E���5�a��%dJ8���Qb�rL�cc[�m�o�r����$"�b��b
�wdE��Y/v� T@1O"�h�aV �]kW�&��^�{f)���[z�F��Ұ��M!@�oe������^;6�R���Ғ���:.�׻ m��̈���9y%���7�����ի�3Fͤ�}����g\�Ǹ�2Y�pd����-+�,���R�USj�n�
�H�.��n�G�&0��!+i,�]d�<V��5
���t&V4�(�T�K%T/;*��m�sp�I�c/2�To\zM�R��{.7Yj�ƛ���h;� ����f,Bˤ�-��j��b�o7Q�/q*4��"H� F��t��@��%��.�aw�-�Z �wu�3�Ef�oD�{��c�R�3{G�C��ث(ݧE<�h�h[akw���]�6����ie5�4���SB�a���,T�0��n2�����2[t��(��#x*�b��J�6Uy$r�L�
���jh�>�`��5jUv���Dk*jz��9Q�$UO7��f��M��o*i�ڴj�yQ���j�[2�Lxnj�n�*Q{l^4���
ʂ^��R�T��\b�C+�������E1f�7��.�Em�3[y[�	l*`�T۸&R˧Z�shD�뱹,QH*�b��.j�0����͓]@�2�N�ڭB�FH�U]��B���^ҕ�EJ�v-�H\̡����ʼ�ǣ/$c��?��L�}]�4������+�0�2�"(⥻X�]��/)jZ��؄R��/D�[�V��X݂��t2�-���񊛣E�1�9ز�G�X�
J]��pHF*�H�A��a���N�u0�(�nT��� n��-���(�����Le��/(+�HYX�"��oj�Ņ���P��;N�R#j�P�2)�p���{�D[�@)P*hf�,�j����*n��.  �,�^����s2��A�f;����51`���t��t�J=FV�ʽ!���V���VH���?�X��;l���`�=����RՊ�&�����gwj�Rj/Q��E�boأv�Z�pZ�n�;m)&�e��y�(1��q�(Cy��E�0ҧU�C��$��T�b�[��S��28B1X�c2�'ǚHu��^�^�al%�3g^6ӵ�9/u�F0�1GE�Vt-=هS-���stXs
Q*W�	Y�������ȴ1��P�#�r1T5��T�P�u�l�ku,��Cq�6��6ɩ����7��4��f�+C(�rInѓH��TV��¬ib`�ˤ�i̬x�4�3��v�i6`����0�W�n49�J��)�r�]Zؕ��z�!!��i�i�)������Z�݆��{�fi̠�t�s�9U7vMb��kƚ��p�:�ġ�]�71�%'c2��voװ[��^�����������M2\�VQ-S�!3(KD�&�K�(��(�Z�M*[4���J̋l�w3/]�����d�[��ɒ���b5�x�v�[�S�
R��܈�%�-�߾�aGl\���:lMn#��Ƃ���'P�-U�����YPˊ�`EizN=U��d9�.��#	rhi�n�@ʖf8��!�aե�e5�M�Fkي'uO�`�/wD��Ӕ�h��AQ�8�X �eb:�HӺ�5aDmя�YvU�fd3��m�^"�)��2��v!O)�jVB�zkvk��u��m]���fKWu�/Wɰ!��Yخ�*Sv��b�6Fؘ�4�6*mT��P�MؽcS��w-����f��%#�h��س�N=Vpe���*g6���Ks˓����%WY����k�2 ��%�$�+������S1 �D��E�S(##L>)
e� ��8�q �%  �@L�bH3���
FYH��N�i�8%D�m$��912T���(I!����2Y,$� ��B
l'ab�"h�Y(Ld6ЕQ��4�j� �5�0�8 �(S�6�"$�F!(E�&D��.6�s�(��?�(��u����uY���8Vm4����ue��+h�����ʯ3�]ͧ��3�K�W+�O
�%�cu���K(�q!�E�o_�s�5��k�`��F��O�ξb{��*f��ۙ��A��+�W�Ծ7g�[oE3۲8�����K�Z�k�����l��fbQ�T��Y��*ʼ��Zq�e��o�^-ֺ.��ݼzV:2wpKpe7��xV�QJCգ^��j�-iNڏu�_Wf��9u��)�β���i'�G	1d';;��w�.�
��4�eΫ,�.��e��ϭ_u<}s�,��̘�5���.�k4��bn^Ru���=ru3�)s�yɛQ;يl�DީwF�A̼��c=�b7�1�wQ��	,��X\���b<��+o�<�Y�̠V����9���Y�U��G����&ې�!�`̩�f�7}ːI�4R���7[,-Wa��tnhʩ���j�%�y�}��N���ן��<6m�e��:Z,V�[�Y��k��F���$0��.U�Œ�tΈ��e�)h��Aò�Q
U�Jav�T������u�����9�U����V��Y�%䷇������*;��]��ݎ�Srô�=���_Y3�w/4��\�K����{÷,MJ�!�|/{�2�Y�^�m����>��U²N��PX)V�xV֫����rX�u�]�vl���m:Q�
��jWK��!#t�`��$F6'4�W��-�u;�G'O���d[K�����vr��bL���rN��\�G�j
�x�si튖�<N��5�D��,��K�wF+H���K3���9t3N�㵽>��O<�� }��b��(�.��߳5�+��>�a�9�4�T 5:^H6�Vnl{dY{ǝ���R�F��l��u{��ј�����SH�g.a�RօW�����z��v��Y,�M#F�ڊ�=���������K:�5�&K�3kmi�^��E�X��ݡ-Hї���.�'x&f�u��d���Z]y��/lɆ�����V�R��j�7�H9\{�v�N}�ڻ��1jKZ��ūe��L���l���'Uw]֍�Ov4��B�6��d��e���m��A�ܽZ���t5y�:P��q3{^T�QH�V�vU��2]�cuL�7{�[bI�;�%�s�]0ݸ)��ArݼܺJZ�L�!�	��t��;4Z��y\��K�5�E������Gث�W�ݮY����hANJtG�Wh�(򫗚m���7R�z��Q:̰�-Р�:Se�ŷ�WQ#`�t�:���8-�G�tU.FiK���;��cl���9wi��1�֌�SmV��I��v�}{7ʊ�^v���'�ڜ��U��;o%Z��cٲuCL_v��H�^��G�e%}]�D3��6�-���Řmռ D�&��$�i�_is�å>�Df��6r�t4^���2D��pS�A�c�u����ނ��Ĝ]lg�P����ʽ��>��6�/��w��vo*����{�)���t�~���Oq_c�ǝX$���M�޾C�Z_w4f k��jּoI]ٝ�]YyPvs�5��S@ܾXﷱ'	�f��V˚N�6�T�r�D�U��Y���u���'��r�`���k;���vH4��#�t�5�[�n$4g`�k�;5��Lˬ�����ԇN� T{����H��9v��)ꆬ͸�_u�h�2�cM��W�c��5�2��`��	9wFʆ13,
�:S��ƟtrI��$��})��7;���So�6�I���$��})��I;����)U�wғ�;W�'�I[�3�s���)oj���B�.3�uuk=}]���jC�`�+k9-��y�s3�](���3�妎E��(;�U�81i��J�b�C�Hૢ����[F�2��(��ze�ؙ̼N;�� �vf<��=F-ך�s�R���ۛ[=�$���T�����u�":�ǫO]>oS��ܠ��,u�[���c�`]��uf>̱ז"p�Y�+��wr��׻���yls8*o�zf��D� �d���x��'}�m\��Fe�x�����-�ރx����&.�)��!�ݫ=��܀�Ԇ90Tх���)<�E�ʚ4�2�̦�"���^�U�j�l�Z9}�n�u��h)X���f^cZ���i�*KK���`RwL34e��ϵ�r$˒�t]�X��C5Z���"�֚͘�+�1]&�n�ɩ�A�%nJ�ϫ:�NQ{5�*��v�ܸ�
��Gs�n޼vu����v���y�٬��6�6l]�(�/'$��.3tm`�{�f݊���T����O�ru[�y�.������q�=X�aĭ"R�HM��x��=*ɝ ;�%j�H�:�B�]�����M�+/��ߎ=e�br]Y�GuuP�ԽјU��VC\3��NaY41U��隰T�}b}��|"��*ΰ�]�N���m�L=�A���5"ݪ�is5m���ʱ{�+{��4���Ir8c���V&SJ1�ܽ�����4���7X�:���x=�����.��RYMz�t��:�$d��ݨV���;
��A]ؤC�Ǚ:��{Nt���VQLC{���n
kJȔԻt��{2�Bg	���S���\�{�M�I�j��2a�pe�Z���tw4h��ZP+�U#qa�[K�¸��<N�{��//tm�ͺ�!�B���R��F�,����*|Jy���Y�S�-5���W����a.���mL"e�DD6�˝ut���ޠ�]�k3W�\����X�ݴ����8�����{B�w��]���R��C�:ġɃ*ɾ�5��d��`z�u�yh:�0�H�u�}�(h�I���ݨp��찤^���&����u��Z㯝���<�9��Z{�s M�&�.�)�YҶr&�^ ��լ�[�o7�'u:b�t,���N*[�����|0����wV��}���B7��N�G�T��T���5W&,Zp�J�u�7�)ܾX+/dVp K�x))��EΩ�Ƙz�V�GR��Ivԋ���i4sD�.n���5��.��jns�t�֊��m[Iw;�ߺ�.���,erч:���I��
q�`�;N]�^^EpqyJ����,�����cj�&�::�`�Ud��GP�M�[+:V�����E]2z�^��&��wY�J�\��B��0�����|��U�W��T��D5���em٧L���TĀ��-�x���|�hC�6��[C�����D6�P���,vU�n�m�f�ڌVuf,�\-:�5��f����$�w�|N�y37tV�c��1�n��"\�!\ �U�Z�����ްi�������1tfΒr:��$dI�Y�7W�jU]�L���D�k�۠h��u��]�PҚz�5�b�c��ڃ�k�K���<-��$K�O;2���@��a�X�:� ;��6�Yc������,��yk�X�f\��WAI6f���l��BwV62t5���5�P2�骳����Q���i��_�Zu�wr���&4S�������E��ɽ�<�#:����<�.]�#�P�k)�-.����\#�X`�#�6��Co��++�Ȳ4�u.rKLq���2ӥ���9��8G��@���9��'?��v��]���h��� �BC�U>]���O#.otʭ��	�WL��͏�rk��M�iq5h���̧F��X���)���<A�X� �Kd@����fU00��0*�����$X����Rqz���3�RR��.ĺ��)�;V�_mG�fY�2-�m`�&� 7��9F��\U���3����=��*.M�	�����gT����U�3t6"M=R�W="�^�Eޗ�V���N�j��� KRډ��C�~i~ٵ�^��b��	��"�WA��l�L0�^�Wu,�n�3΍�����m���"U�@+��eїC�<�ۺ��u����Xh
�n���`�&8�tI�%w],�@\K�"��������\픦��S9_�V\��mr�]�^��"g_O&��ް7J�2��)[�Ja�H#s�pY�#Yq-�kq�յ$�Z�����`��5�U2K�#�KW�7���9!������_[U�Wv���f�l�<�	���Y@���r ��ސ�n��ݹ���}�	8�.���ܡ���Дn���<�ou�g=Y�v���'E��������Q,Aw^�{A�5vbO"�en�t�v��+�-$4�d�{�d��R�7��q���QV鴬�K�4;.>ˢi�y,��a_Y���!]b©�t࿙��nڱ�oN	f�
���4d��U%4�\紶�+�a�#Rc��0��a�5K�(:���4)x5��A��F��L�>,�B�*5���K�}ؕk����(v�}0l#�c�Ҭ}}:pz-wJU�6��>Mv���2�#��Rn]����k��Z��K��W�t��PQo:q�0�^�m�Bhә6��K����w�z��X�_9蠋�"��,����|s��b�ޓ��m������E6#�[.0�|���J1F&[H32D`�<R Q%���\�ݱ�@Re�&�|	I�$���	�ČL��i��H�	�"(���o����<��:������m���'[�QQ�>�l��]�y���ݬ�s0�$���v���%b�2Vc�#ڊ���Bh�3�`�WcY1kkI�:�B��\P����w"ks���;��;���:�wM��U�W:�;`�L��W��ߛ�2D������4��j+[kQ�t�ԙ��W#����w{t��=Ǩu	r��5v@-�o���c�h��&���˱�}9�4�b2�ٍ�s.L��3e�z���%� _��j��������^���p�	 'h�@�2���0��C1�	�BDx��< ��/5�u�뻻�W+��5��j�r��n�lX�`�ss��חs~��W�nZ�~�W�����[E|wb�/�y���Qh����.Q��-�76��v�5�T�g_���j�h-˄ld�Q�_-�h��F��y�wvدwkI(�u9�/.W��b~�?n悶7�na]��߯~��~���!<�0��a������`�m�_e``��n�ln4���7{���q+�ǻ�����n�)��<ъӥE��ޞ�<��t���U���u�qI��>^���9���raL�b�b��wk�f9�S�jMBk�N��wv��)����[m	7���u���2|�uf�V;<�Խ��ߜV��I��upE�t�F,?~z�5��Խ�?�b�L+3�R�$=���Ӫ7��lVE�r�|q�\�SM�]i��@��%�Å�I�g̱��̏p#�e]l�9��\�%q�{<�S�m�/t��;�.\*J�o����r���9���,Fa��Y����$�}Ů�n�m�+���$ęL�˴��E�L�(��e�D��qS���B�Ա!��v�Q]t�}v*;�w�=�����z���Vh&���z�я4��bBt�2�3��q�&�ox�c��+�-[�:��V�������4Mն^f��G[����U<�S���9M��ɩ'�f���̸۪|�t����U��*�z.ܢ��fc������pc�˼��J�R���܃��W�׼6:w�ͤa�d歬>����߆n^��	�B���i�W�㞺sw��x��_H��7�7�ë|��@��ę'ȭN�N4�͓Q�w9��`��-����N���f���q4��fy����w���U�)�0���46Qv��7>�xBz�̹GqɛwY�g�0��8���x;=����TS��d~�粆�跱<���{ޞ���d����������8���\���hZp�tY��oy�}ޤ(}���U���EgTBډ�H�J���U����M��#nT�*ɸ4�z��B���ŬU�ܚތ/M?]-ڬJ�E3��u"��&6��/	j�˰�*ű�s��PXS�B]I�[���0!f��S���m�k�5`&R�y���|��}�/"pmHsn��Q�;�H�s�y��$����Nۮ͟z�ړǤ�l��e�0dA{L{2`�˭@�����é+ː�y���_'��s���ϖ�=*r�m}�U(n�Mek�<���g����~]���z��p�{�Hz���y�W�!����*;��Ϋ�q��4�^A����(b�y�u��m�����{��,�<3[K�م2Eў�׶��z���7t�A솻Sz�S��,s�+T�Lp�k��y]N�"w�������Oo�.��Z�S>+V64$����ݗ˷c7(4s����)�c�B5y��.��HXLg��6�:e�</YXf�.^���g�a%D\�{k��O��ڬǋO4��xG����޳��/h�3̊9�f�A߷ڷ����4P�&,�B�띬oZ����v���?f��||>\�}��$@*
\q7�\Y^�,�`�;m��`�EǴ��*{Y�#9�1�z��>Ө��\:{��[pK����ۅ�8����!�������Vo��CWD��&N��4|;a�i��Nߖ��Kُ��n5�s=^�"���GA����E�a�Z�P��u��|��F¤���!V���-����*��z�p&{EUGVyWB������'l�d��1�����"���ѭJ��}"˙�����S+>��U��+!�ɻW���޹�"U�Q��s��ov�e�9��,1�P���a
�@xB뽯\�3�J��Ղ�[���smy%�+�7�y3�[s(�Y��޳�c�{mB���TC�	�C�ѩ�M���KA��C������f�8t�uY�J����)�B8�f�vބL	k`�����V��6iUK�cZ'n�qH���"ߚ=6�W����G�b�m`(>�`]rN']������_]2�s+򂜝��-S�νn6`���8�wG��7[²�[��V��-P��0ky9nq��j��{!���U\V��l=j|���dM(��,`�@�ݧ��$΢�k
��X���[6q�XTl�BݥC�d�.����Hf9�멝�:ɁX���E$�������Y!S��?h��AS��c����lRU��Q�P�μ���e�h]p�E�v���k*Yc�on(�f��7��{fX|S�R�����~��Wh����b+���t��Qѱ(C�6��0���]i+@M����B����N�|�o��h��ag9J��@_Q������b�����ϫq�@0�\�%���#ú�H} T�ۏyp���y;��]��n��x�0ՠ�j��<u@i��d�������Fǽ$���@�ﳩ�g˭UQh���e�����	iNcМ��Ø�!���u|�R��WP�u�T�wdJ0��w.lY��%̸�7�*Y�pMS"�"N&
8K!*Z���icP��8y`�IX�3(��Scy%��q��
8�Xպ��-��Y�r��I��L*�wV�֤���N�l�B��lХ�e��[���{�z��>�=]����ݫՒUwu|2��ߪ@�s9Ԇ��Q���~�G/�{�6���E�׻��)�/�U��]�u�|���~z���w�yX�7�ƞ�ͼ�7���^j4n���t���o��C<$�!'�s�s��Z4�C�h���gQ�I�ý���ᝑ�C&>�xI���Y���~��RIO��?Bl<4�`����տU�f�>��#�H1p��[��2j���>�ctbN�\d�F=5]Cw[|��p��ϫ�o��c�3��{�!d��ֿVk^�]��k{�d�f�����Eeq@��/�}q��}sm6�{)(�������UV:-�S������BBj���v{��|5w�mv*?D��͌�xus��-G��F��-�ᶶ���?��Eu�]���I�1eW[��8:f~<�
k�ln�aٻD�U��+��q�o8C�H�\����G��U�ޮ���}�!��^�ٛTގ�ȕ��G�k�z�V`��d���mޑ����+_�~��a�t��7�ҟ>�������QK�\��>�پ*�a;ۦEJ�����1L<�D||�L�'��kxoP8�<��<<��LD]�ku� �L�7+s����o���:	�sX��摌m�6�'�
Xci���W#wW+���>�NK]�[Xw~;�w�F����D�����o�(�"���\���}���o�y�6sE"TD���)(�t�t�i#�V=�[�r����^!��GQB�19�Z#xGx�0�1I��!Z�N5Ņ-7��<A�AS/ELCCknw�;cAx!h1Nb���E�
ox�Z��mb�*EI1dGPʈ\��?cџn�uR����F�A�iS�>#{ՏQV=Q�����r��M�/�o�M��P5�k�I���KH��S�S:�Jځ��%�j�";@19��Ls���ӝ&��$V�u5H��Z����`� �s��tR���- -�iZ�d�*.��E� 3�'S�R8�NiS1K�6����g����-�J����5jQ�(b)�5�x�@�M�k�����A����"�)Qd�& `1�Sh��!������ŮN%���ʘ��)�b�o��g�*�m��"��[�.�*��Z�9��y}�D9����Ch�D��v���cT���tEN`Z(k���� ��R���!�x!����/8����x���"�P���E78�6*
�\B�@�Y���]mJ�CQ6��nu���4�`��&"���)x�P�1- ��d�&-�w���6�}/H��$"��x�����~�>��B^��-(���?� �8���
c4�b5Hj"x&��h� ��ZZ�	�t�dM@/+��t�u��8S�	h%�b*q�� �zT�!��$V�A�w֯����^*jq�1���Z��Cxm0oJo[f�1z1Z��őd37�EM㈻@�!�R�@vޖ�N`.v�	��Cv�|[��嶱�LE�D��E��]Rff)�@35�'1S��s�7ҧ0��Z�N ��F�0J��S8�x&`Lҧ0 �����o��v���Z/��w]�	h�Z�v`�5�aыO3Dt^<��_9=Q��.	̠)�voE��h�=��n3?,~�p?��:��:�ف�w0Dؤ����uclg��b��T�gvM�Š�^lN��8�/{7@�
?Ü��}����=�UC'��/��M�sR��"�.Z���v��'[U�!U=O$���70ݗ{E�B�U�u�(�y�v�z�4O�[�����kB�������@�BH �g��쉧��+�����T����0����.�ѐ��H�['��"a�Ǔ�]�{����|*�$�Zy��S�1��ߺ�I2������᠄Ek �TOû^y��W(N�,D�D1���13�K��xx{�0�C*�;ԋ��.�FnH���=�ͨ���D�u>���y��oL\�5+_)�v禖e�7u=Z��c�t���ǎ�Ů�]��O��wE8]���ul�����Wb}𿌿�i��"���U��3�^�/��Z����-��yr׋�A�3��&9bΰ��Z�B���u+�����2��X�	�5{f�<'��4������^�j�V`I�a\������f�]|5��	a��[����~��j{Tަ��Ӡ~�gT��
�E����&�>��6�{f<���쮃B[��S��+k:��N/�70�+/�J6�ԷLm���_���6�b���À5]O�D���c1yW��pGV�yW4;-v���p�eQ��j3��?�������0�L������9��~�g�t���{鲕�����=]k�ry%�%]�9�^wrt+>�����Z~9�t݂~ڻٜy�]�|4�N����������٠���0���٦}�K�.��OS�i�;lS�A��W]�����3�Hz���=����u,��>dM��~u�b�.q�HRïk������d46��7Ĩ׶�Q���1�4�ͦ�@b[���)ʲ��rz=���b�8l�����Kvn?+�9�#o*Y��o�j�r��U_� ?�)&T�'��Pe9T��lЩ�E<��d��ó�/�/�S�ŋ�M��ueځ02�z��t��Ϣ��s%0~��ӭ4z;MZ�
��L�wV�b����u�]n�0{Vܫg.g_U�4�bZ#�����!�f���.E�k�E���-�$s(�oK܈z�9Ym�f����/?v��&XCl��i4Pd5�b�D��1&�m��R�h�,���\���
�D�V�.���p�LYq.��bp^˫w���e-n����|6u@�c=t��(�x_6ghA�*ē���幽k:�kr�Z읥&0aD�OfM�X��8�37��v�.l����//n�+F�Eꢰ�r��Ru�����hz�,`��b�*�6Ι��9�v3M`#A*�6dd�=��w,Ҏ1�Y$WyEX��,�&whXF ��2�U�g�?\6;Q��"��']˞����:Ij�Z��4�Svc	SW�VO��@��
%&�!$�J%"�-�Pl��I��
4@���C�r��)A����R��Tn��<���"ՓiRPy�t/�^	1��Pe]Ƃ�R,,�<�h��M6�Ӽ�������8��2�'TLWS+2d�v̳l�KB��8.���e�v.�b8b�S�V�#O2J�
�U��I��A]��{5�P�#wLЫk5:u��l�z�Ğ6���uX32ɹ�;�e��&_�M�����2��-�X�1+�Ł����W�c�k�:`���9��rw_����O���-������W����� �w,|�\�5�ys�W����޺���{�\��rצ1�~u��|���n;炙�|����{�;ݞ��7����,]�P������E)�mz�ǖ��)�]��y��H��w�{�����y̺��U�狨�7�ݞ-��a��+��7�_|��#t.�=�
��Ҳ �k��AJ��X���X���0�����6����B'q���O�'c��z�u�{/>�R����U_��;n��GP�=��`���Iw�U�|˗��ּ��f���U�x�ݺѯ��k-|*���p=>�̘:r&��u�J�q�%i�o<N �8���d�ٝ���M���Wl�� Cx�<f���9���T�ҭm��nz# ��ڣ/�3���XZ1I]�9ٍ�fc����,*}�e�u��ɚ>xl���Cxvuݲn��[�7�U?�(��z�v�LO��a����)f���;�mZ:� �ڪs^ƶ����ڱN�D[��=�k�@��
���}0�@�h�=�(��8�H[G�np�`���r��79$:�q�szo���:sگf��['b����Tn�i��>T>Rs;�e��g���ʯ������w�ϭ5�?eݫ�'��>tmJ@���y�}�W=w�z��Ӽ����`9ᇂ�p�=���6b�F�z+D>L�U��nA�s Cc4��4$.�c�߅lx���;��o�N[����p��(�Ӫ-X�� ��a�m;���K�/�^�>���f��Ѧ��.�	�����SU��jqGf���_��.��B�*�U��V�9g����;yn�w�9qZ8����n�I�U�^����זFC��UW��b).��[5��ﾁ�_G>�u=s>}��6?�����,v��߲n�Y�)�߄k^�k���q{�*�Ֆ�_ɵ�����Z&8�/,�E�
�0�]u�c�i�BS��n�`�y;���{[w��u�yK��)���`�K����C�y�����9���Y)���{��vW˔���n���v���.�?K�Rj��m�������u�-�%�B���"j}Ks����/�����U Da��Lf��4Zt��8�r�4���z�}���;�'P�S�ܩ]Uۺ�<��8����a��mè w	$��z�"j�Py�.M�lk�W��S�{����n]1@��bg6�fz[�3�w�^ר�Z̓o���
�ý6s���W�}�	����G|-��oM��8yh������(C-~�/��J���+�,��u���C��3*�����	V}\t�H��N݅�K�{��5h��y�6�3�
"gX�>�o�Mv E"�a���m�dp�ې!�`ư��By:ƽ�t���D�z��Sݔ9=��S�������*[:��f���RƲ}�����P����� ���t��v��剝%��������� ��e��7ڏ}\z�xr�ϗ��}�����P^���9I��H��'�LN�n�B�_Z�!��D��}�y�0�v�(�y�ӆ�p�e�����z��Rp"��"� S���� �!G�P�i����cZ\#z�aDW�Qr/�}�}6p�R�c˵���򺋑 0��f�(�j�R�d^#��y�l3ύ!��Τ�A�,r���G�l�[C�:Y�d�y�o5��s�lmgW[�,x��õ��"���t����U������Z�}����bt�N���NK�~�����D:p���W�Z0P�7F�� 0��×���-r�Y&�~ߒ�9}?|a�A\x�g��ʅ��)p���������]�0�{m`3�qč}b��R��?��w�g�S#�����vmR�Mg}�%��G��g�y"�pm���������3=��˥� �!��ڰٳ�<}��c���缙�	}����W�>���i�����>:@�}1�C�P�+�y�s�u����y�v��آ�_*C�2�p�8�:��h~��s����S3Z?�Z_��:�� ���W(��n����ؕ�X����gN�嗿0�rZ�f�q4C,R��"��W�����r�������~?f(�t��<�rChZ�f͛ōYg-">!�,��v���P��J?bEC�c��@Q����>H"9��,!-'2��4mr�V�KjƑҎ�tC$��+��G�1h2�DQ�M�������x�!���'�v���X}�F��<|t��E�e�./�
ŷ灗��$�y�@SMz�+L4�u�&�fwi��p��n�ܫ��_UW�I��p�G����!�YǛ�����X����Ф���!t�!��D$��σ5�Fš�����x�,[X��K������8NC̋�hȾ:y�c��x^�V����OU��ʮ.}#��3�F.��Ļ�v���i�Oǖa�$��@�f&/�?)O�FE�}���*/�5��?f��:і��𑸰��f���a�h�R^�b$��!�6��	T��(9�����7��@fx!�#i��a�x:�����yu���bS)6k��)��H�ǔE�V2����Vt҆�jץ��G;:=���-n�1��@�s�I6����X��3*v7J���ܹ�$�t���pf�th�<"�Z8v�8�%v���&A��-\�(���-��^����e؟?ܝ0Ǭ�^��G����h��5[wkBf�%��g��v���ӽ�wVk8��Σ��MF���&b�,v�U"���[�H���]O�W�֨��}�I�Ьkr�m^Tf�#d����v�Q�.ӣyU��b�Ǎi�6�2�әM�w�i�m�7�^�L�ޱ�$]��8n��bH�����7��R�	����1��wx�V[���:p�s1�4����B����\ж&�zJm�ۧ��i�[����Kª}�i~[��(x���t�F�;|����]��HTm��RШ��+�7���}���[޻Q����y�����>�r��r��}�U��/��n_*u�[�)�dp�D��4������,\~�ףo���������޻
�'��j�>�����u�ܒ,���,��~�F�:�K���F��U͹��8J���P�C�"W(���,��#��]���x��B4Q�[$#�ԓS��[#����Y�v�50�c��Ҵ��1�ʁML�DQ�䥰��N�}!������B���z��Ū(}�n�<$�#p�� _�4y�Cz��CF�<�FȠGe��OMg_��i7�8V�0�Hz�ms��.R\�B{��W۵�ŧ�Q�(Fh#�nׁߐ�/�z.۾#Tp��D"��$it�C��7=��>�dY�J�Jv��q{o+m6�)t`�';!WS��Ƥ�T�T{4�,ڢ��/���*+Ý}»�ﾪ)U؛��%�Đ�Z�is��u���!mpa��
�(�˴;�a�-J["E?� 8 x��6�a�����N���/� ��0𛠹�VM�9�G��U�j���aÄDq¹ ����ϝρ�������˔s�P"� �t�:_`�I���|����w�H�K�ސ��@�)�j�ܴ������:��ݞ!`������g�5���PC�i��l�h��E�	ڲ:��>��N:(3��/������ɶ�4*".�M��x���L:I5
J�p˰@�P)�d���&�� aR���4E����ٻ\�E�� �p�ۛ��[��HF���nj�ks�|ҋ�
D�<������z���a�B
���G�B�V���O�W�k���ϛ[|���M���b�#]���}��6/����.������E�F���v�ߟ[�,�|��p�'�d|I]/�"�~��[/��xMd��*�ч����
]�7V��4+�mP㖅�f�D5�><&�±���?4A<�X�>7��!d/�������&��0%��PuN1'O=�s��9��\�5�{7a$���UH����C"G>C�	&���+d-Ż�/�6 � ��!���R=!����f��s���pGwM�l><�D����>�b�`�5��x� �ZHD��W�)��#�_������(8wt�ĝ�AS6�ʏ$�� <C��C߭l!�哇�C�xy��*��y��4��5`n���i�����Ml������.�0�+S
#��"���b�e��������O��[ԟ�l������^=�15����|c;�K�<�so{��<����z�*9�.�+GfHn���UP�՜)���R$#F��A	����٬Y�"�4G�@�0�6:
�ÐN���G����}c	ߙQ�Cㇶ�قz�
k���!�&�(V�'�.������y]��K�<�<�$��_^��y脤1����q~D=@B���\;��33��*v�
Wl]��C{�2�z��@$>s�z�f�.n���� Y>�}Gd�������C�i�C���&@oK���Z����s�aM���L����4/�)�z�Ӄ�fp���N�|�by���n1�٨gk`���F�eu�$��ဧ�:�0�Ǉ��W^\�}l���\������ʒ��z�?��b�}2�k��;���YMq�O�c���y\��cˠ�ګWX ��>�|�<A��:&���ya�f0��4�3�	��Z���H�D|`<G��cy;~��,�]\ ��1��!�\c�7�-��1r�}�D"I�&ᓟ,�dX,���70v�v�ɽMȬ����Ó�aҠnoc��Y�?uv�_��b�̙ƛ�l�� �F��B^��E�ђ={H�����,^�EV�h�9ދo}��۔5�?Bo�ʜ;x�[��#ԗ�6Cڞ�/���g��F���kY6f�[P�g�y�s^Lc����<�Afܳ�"��h`ˏ����~�"���@����Ii��=�=��q�	G�#�����ڦ}����d
J�Qc�n������\�2Y�b���L~`]���m ���"z �<���x�x��������"u
�4w�|V�6g�?Qf����3�k�6G������?�6
h@aDz����+�5Y�[s.l�>�1V�n�G������ukyЦ��mUܽ_���g��B�Y���ϒ"ȠY^ǟ�wE����M��=hKE���g��ڽ�*���ǟu�׉���\ia��k���L��!��$x>�cM%w��ud�a�d���/��)�������ӶW�B���x��QB- ė�7;6 �g�����G�FG�GŅX1m"$�V�a5@��G\�������4��'�y��c1��6[{�c��G���d�bxO?c���n�$u�3�kN��.�2�fMD̜��q�1��='
�[�t��q��/���A[���6�X��<�7���jn����� �@��E�J���gz���	��7`���Dֹ�B���9w7~6���Bp�:��kU��?E��Zد�|���'�B�C���HDC>C��~����A��6F�d'�x�>o'ۛB^����"a��%�H6<��;���:�zGN����g�ȳ�l�B��,��hzh��ė;>a!Zx��>8I��h}W~��<����*�������������Ȧ��ǿ3���b���5�|����Ի:��Άp�oqgq�T߲�(���^?�jA:I���C�#}����ڢ�Fg_7i�<8�<� 6�w�[8A5��R���>}�����/���/�- �JC�񢻬a�(�K�~��W+�)pi�Gbr9�\&�60���M��b�d�J�'�_�G>��x�#��؄NB����CĐ�C��aD	B8p��tȫ�����C�©��|���d7Y�0x,���x�
��<�W鳤2���(��-�|�I$"��KrBI����Q�Fd�ʃ$Y^��_h{�
"��(*+�?�s�+z3�����,�Q�8���顳��I�h�̬�ǜ5��W�t����	]�`յ����n��e�}�̲�H�ݭ1��3I4f�iX8pO�_+�r�{shı'r\�:��8����T�T�/��*�l躹�h�OC;O�J�B�ėx�. �pl��;"ř�m�L�>93���	;���>Pm�Pޥ�l��ά5��41�J�i���jINt��3%���0Z�������x��ޫ����$zvn^-��O�	S3��坣��ކ-�
��r��d�U��n�E��0�|��8Ϭ�C�a�0@�^s/��xm���)񺾣<�$�<cq��ʹHw]�^Ʌ�/;��@���v�+���B��/z�q�ku.�ۉ�-l�U�z�;�s�NN�l�u�ؾ窯��!�����ɹ;��������,��&����&)a�f��u�3;��A
����ER�TA���P�B`����S� N��,�Q�<h67�w�yt>��>�]��{�z�y﫷����1�s�]���uߟ^��������/�Q��7��ܽ/}���;�=���~{������Ww)�r&f�%���.� 4Q�T�H��$�`��D�E�)ƃmQ�wQOk��ҏ[ښ]R�u��pj��ܬ�n<�ms�\��<1Qda�|��ɽ��o��p����������֕�>CG)�����6C<%��:Ak��Xd?��f����ƃ����������5�HX<�!����,����m_���S`�r[SRq\�2���_3�{,m� ��:M!D2	�զ{�|�&�e�oo�A��9���DuS���ʾ�sM^�:��{�e0��Q��o���D]!�NܴGF�Dk��& touܨ#�v�'彋n3z�[-[=�{;nd]6%��v���8�Y�|]���X&'ﺩ��g���>�c�3z��2�_!׍QC�sP�X~#���{Z��!㇟b�m�@טή|t��j�J�Z�<�a�- !�@�b�w�ͣ�Y1Y�#�P��~��7�~7��$3�z�v���c<g�����ה��7�t�<@�ư���G��t���J2��>�z��,�>��
_�!���յ��w�a��v	y�O��pd��W�iy���G���f�ɾ(�Α�>�G��<����uCH;�����w_��>j�O�s�]NZ����g?��[��S��W���P�qQ��ύ=H����&f��a�����KJ��'���2m�V*-۰33���%�LgW���iG�jr��Z֑�u�@��A��6�{I��D�Y���HyW꼯��,�&}�U�� �н��GJ#�N�l�B��Lv�'?W� qa���?�ڡ���C&�U4�h� E�����px�0�R���C}�a�t���ޮe�hќ�gO>j}�w����G��Hq�Bv���Ņ���3n��oYQ���t���6gL�C�����}EfL��M�ݝ}E����9���
 �(R�B#1>?��>Ӹp�_�Y��ĕDr?�"�d^��ޤNoE�=�}�ȗ$\T�<�"��v��Y$Cdi1?�4E;y� a�Xn�i�#�P��}�2-$��j���u�I���Є?b����#ba\��a�Z��O��{�o�b=��g��/��D�����e{(�t4�ұx;�O{�6�/.!F��(�|�hO���������ȅ|�冊!r|I&�3N+�(w�FD��md�Y�
m4�q�2�����.����K]�s7��٩����Iս�~�+��@�i��+�3�0ZFuz|h�M~+���=.'�z��4HgT���D!ڢO�v��8�8����m1�0��Q�ha��m֋�]���xձ�iN1��-\�Ol3��.��Ij ��� ߐ{�A���K��~>K�0ay�Qh3� �����߬����j��Q�c��G2Ni�4W;�a��`�n��+���������%`�YX>� �)*����3t��a��%��xQ���!v�7H�?E���^_>��h^ខ?y�M>��v��2��8l&��{�Q>�� �ý;��'��y+u��s�Z�"B��y�c��8�V� �jۤw:b����C"<G��w����+A�&�Rە���	�A)���FE����>��|��NԋqQ� �K�=)R���GN!4nZ�N5����qq(]�s��jl�,�YA��YӤX$p��{G���O�0#�G��"��#��[$��|Ԅ�pѣ����Ƭ���<-Y=-�:�G��<G��/�"B�y!��p��J�{�G��U"f0M�ƚ,�G�b���ki}����&ge�x��Juv*�C���!$=:�ٝ��Υ�K7W�����@������Ϣ|�<j�����Q�H�ya�B�����T�i�X���qX$5,sc�vv�q��5�l����[L>�V�IzF�-Bs.ZOT:�RF�uo�/�g)���r�^==<���}�D�sU�6�j��Z���Z�k���o�o���lI/��7�Y��v���,U�o_��,�o�(���r�����o��M���ž�Y����u��\> ]]�xW?[?(�/�e���lO4���e�f�O3����>�B"���(w(��`�=돀5��E[�f~��V�N����?��w�Y�
����t$�;.��Ѵ�L.g"[22+/'��8!ҽ-�1.��W֨��c%�B��٦�L�}U�H��=����W�lW>���Ԉ-x٨s�&��"�1;7ގ�}(̽6�X�G��+yv����%��rVQ��Z�{��U,�r�ɸ����5�f��}���W6�ռ��|�W��5Ȉ�þ�}��p��Csk����/�:�a�r��L�7 �T�ݹ��A��PF���ki�Y_z6����旨=�s��N���	T�Hu��oG�i�i.D��6�: O��p+�f�]�vy�v�	��#p;(2\B�ܾ��竱�2�,��?{Rg��S�t�Z;�����ӽ
��]��/$��M٦�.p�L\j�����Y9Ȭiɾ��m�FzL1Q��Ng�Zi�*�ѥ��Q�wu�{���Q9�g+5^t�zD:��/d4���y�GeC7mm��qfT~^��{�h�#�W7.���bؓp,�62}ΫA��~���_:�^��y�Β:2�qJ���)�u�.'4��m��?+���GZ�IVZ�R�����ţ���+jY�,�W�k�B�{I϶�,�_R�Q��< ���U�3�j��	Y|����,��=Z�13�D���9'bJfK�e��ַ�j��/�ll.���T0�2��h�4��3³���GAKN�G5��:���Va��CǞ��2����0[*��YZ8n�k����]]U�O��Z�Y��9�JC�ܥ�h�:�f�ѥ{�#�>;�V�aS���:�r;�۝���F��(��J7ϙ�ٛKY��#ntWW��IQT���nY:+;B�k1V���ݓ�nQ.w��3z�t�H�ɜѬ�W���q�_5���u�a����еPf����K'5G�6�V񫱦Bf)K7�B,l��e��nG��5r��n����>�g�/�aQ7��J[k��U$�X`������P��9�y�y�ju����Yyk�[��v�!�����^fΙ$��&<�5^��6K��c%��/����вF����J��+���JXz�AP �	�Zd�Kl0N�j�`�E�D�Q0�`��Wu���{�ofu
h×�h��:}�	�0���!�ܑb!w\S �%��g��(�wL'wI˦"��ȔH$�II���$�ߣ&g��z`se���ve-�u�����!��qt��w۸���':V�͒�4A΅�3����x\���X���f�D�A7�ֹ>NJ��F��'p�����췋i�,��˵Y�r_<��U5;ȷ��T&�{�	���<i�N ���ܩ�*C���6V����"�������e�߿b)�0yy[~����н��n��tp�?���B{����	�oǼ�5�5?�_�v��̺�7�4:��&����#�j�������ռ��[�R[ے{bf�&wJ��ջ��m�t(�����:�!�!��Y�;�{H߹���+ϕ��`. mm�T�K��>ֿկ�HG{��'����[�;��5��٢���Ѭa)��p�n�r�g7�<�9�B��		X|e��W��3ϸӭ����m�+\U�(o�����+H<��Ù[b��J��G�Kt+o%)Gܪj�m	�tDѼ�i��7�m��� `3���p����w%����I�8e�[���U�zӵ�2a����Q��am�Y��VMC��wa��f �t5�nT`�� ��\�?>�:���o(������j�u2c��v���� ���E�m*9�_fO������B���;\�.�E��-nh�����rA5=]A��_�yyn���ͣ�壙�O���}�tUx:�����~؄e T�n��dͫ��S.32)=��w�٢�#��X۴�}�~1�.}�o.G+��]K�k����(�X/����,�㿌�	��opi�U��N�0H��Yҧ2$C��g���_��K�T_Lf�M�@��[�cF<��o�wU�y|.7�{��w��K����mZ�}>���B§*�ou�ų&�٪��V��\��U�tۉ�;[$MNA$0��?{��L�r��߭9/��r<A��ٹ����R+b������*f��[����V��pjp��xz&�f0��l)�J����k��vˁ��
��6���`��5Pwd{�7wH2��S^o2p���=UpY}�#��]�K�mdOt��#��D?)Z��7sW�����?��C�[��k��,�s���8�T`�	�+�"8���l|����f��ځ�5��+�t�s������%���n���@�?�W�٦�{�S����}���:�a�-�~�D<�Q�$�A�?���gk��w�$�za������,X��iٖ'�yeՏ�yS�O�G�ڥT����ʨ��>�	�i��V�i�Ǽ�F��]�Bq8��6
���w2<�u\����ܲ�=WGNK�c�s�my�^��Y�*�ێ�of��z�����%�\�a���oԺ���ď4��W�*��ˊvd�;�
乷�_Vlm�Ȼ�q5�Z�ձf>�*NN���Zr���2��7҇[Q�p^����2s�v��G�<S�;D�\��it<�H������ާ레�=�9�]o'���C�p�c]k*|6��&|��w�;��b`0���}p��M�4p��XћA���粶_D��פ�Y@T9�~��GX{�؏�Ռ�o�l�UDtla��E���O]����͗�K�� ء����6���)��ʪ�x�dȲ�~����竾�C��MͰwK�M7��N��яl��֌���ۑ�DY����|��nA��wi8h�{*l���'��F���xɽ�{Y��.�ӿ8�+أ����-!v���&z(��+��5�m�7Z��=����͑{�w�xt5wz=<�!��]�L-�U����F�-d�ۜ��� //���o����jG�:�h�3��ꢛ.��OC	��к�} �l���-�S���\�Fg2��y�w����5ş�y��I	�߶��*��N�ʟ��\�q���Ʈ����5�/�\m�ݛS����U\b�'$e@S]�E��4m������guI�93y�)T.p,�Ff�c4tmY�b�����c�f��ތ�彋>�������q]�9�6{dqd������ڲyWc��D���)��{޻����0S ���}�� *�K}J:�*�{a"Cy5�~a8��1aUSb��v��Y�	*goMnDn��͔!���~AV5{�N�S�Y��;�oU��]ӹE�l:Q�"$Rp�3�U?)B\��)Ž��쪂�f&�p)�_2�n��{����*�aw�9���o]���~�!ʣ�����{���FLB@�f&�1Fde���F��LHm���R�0�ɗDt���r�
H����+�%f��V�>v���,ֳgjk�f`�އ$ui��)
�
O/sFE���ȭjrV_X���ܾ�a�'c[Q�5g.+�5(���H[l��pt�+���G�*E}:�J��εu��r:��o�������k�;�A�����-�1Z��Υ�ٻ����o5%I^[B!Օb����Q�HǦTλ�+�+��g,���^[�n�kB��[k�.��y��q�FJ [�Za4[�1D"JM�L$����%!u[��Y����V[�^6l��G!+*S9�t�ux)~0���r�1��,��a��R������H(�G�S3�h��*ʂ���@Hb6�$@I(�R�ݩBH]4��$�
�SĪ�Q�p�.UF�c"���.'n��L�r�R�7�� �WT˶�3��[і�l�z�:��Q	��U�z7�^",j�Z+���)g�F�&wp)��o-c?`��{���n���������;�����Oۮy��k���	I�L�����=�N�W�Z��"�9��^Fv�4 ���'�_9Z���~:g㩞�]�s?;v��I�7�D�h���L¸Q)p�Q�NZH7�-�\ �`0"Sģ��J�/m�b�=T���\#����\��:�u���.�Kk^���8'�t��5/*�^���:�� ��W�:Kz�|��>�6�C�7F4�sh��>Cф;�<���3��}��[U����z�����F&ommҠ:�W~�^M�4OD�;�J��i�^�Jߏ}�X߯�g76��R�6fz�E5iGi�spz�Dq�O�s�{o��'g�b�"�QʬU�E�V����L98�HR��������qw:�}ߞ��߶�Jhq:p�ˠCMn�uik�Z�Ry��&�Ims�3���U��ѪxVx�QIќg���q�Vvw����9�vռŢu����i���8�O2�@����3���1����^��}�*R��&>_��1�ν̫Y����� ��|��H�h��=��f�
TN��+q2%2�c�*YT��o�ѳ;�i7oz����R���y�C��)fZ�����o�����b�m�� �h���ƹ��C�����'=:�� <�ܦ<'��B�����y�
\=T�����uQ���)(�v�8�R'0M��v�a��${ب:���b��NGM���o*�Z'O���6�hԁ�uZE�����e�k�h�-��ݯ[
�٣#"�	u)[Z-�ɼpdN̾���z�ӫ/%N�����R���&W�:��{la�K���Z'��`����e8gL������B8���J��8�����T���d���s~�k����]#d;�=5���w��Wv��l[w���V7bڧ�����*��i��.�O*h+ݨ�2���u�nni&��m32�C����3Ϸ�N�F<�{��c"<+nAҊ��jhaY��%WN9��A;�ȺT���6���5��UQ�E.*�	�&��?������R��Aӳ_>t���g��G`�`ʹ�YX�̘��ft�C�a��GZe��6j.�����	��;�R�_��2���w/��w��<���^�i����91�^4��d�����z�.�s�{b�8e�S�|��2��f�[_O�}����7�=f��/{1�b�7P��e����z9A-������Q��]��b�����gN��黴Z>}=�w>�y����f���w3�Ǵ:vt]�g�w��|FZ��я��O�}�ޖ�i�E�:��5d����H�¬o�Y�?�"ϲ��n��ea�αܧ��׮�n"(E��a��v�]���\�W]��Ev-�	�&���ل�; ��A(�\��]W+��^��e�O���L ��[mO���3��K��S=���Z|n�P��M��V��D��$z�|�quo12t����-K%�R�F◪?4�ئ��܊�yN^�F+����s�U�EGt�Qd('���>���r.�����o�ζ��Uv��ޘ��+?U����,���i��fM�U�}���$�e�\C\s���;TɥǮ*"gQӓ���{C6}13 �`z�f$����4'�A+�G���HM��:e��d=ު�l�̵��Qn���_�O3�0C�q:t���%ͤ��ʽ���;�4 �/Q�Aa�q�}�(+[�k#'�I� G�S��B��Ņ�5_]N���o���߳5܈���X��(��лUKՋ�{{r�)jS�u��l�<�Ό����U����f�D��Ux�({����TUtk6E�]Hi��������עdll�[ּlftM�83�ڎ$�.�[�E�������5��+s�`%��Y�������[0e����s8/��.�K7*�������-���1��hiiR�e�O7�:������d�}�z�Lag�:�Z�Q����ҡ̵wI�h�Q.���r�0/���5^��v_dϞ��{E��W�CmmS�x�;z��#_���3��Y�T�n|O	�ǒD����vV��i��Zu�U�6��q��Y�:���/�M�H���9����{�.�7��UU��} ���,�jNI�̙���W֩Ql��㷸�-n�um3���ʼ�`�f���|POY��E�xn܃��*��]Y9��x�T�!bg`ׅq�\���MW�F<����Zbk���Y#�����zo zd��� F���Yػ��Ŗn���:��0�U�u�Q=[����������&vw�{yO��3�?5j�;&�F܈V\R���U̩A��1l�5VL�(4�}���+���+��LB�Q�Wt�t7�d+jX��>�F�ޱf�5^$��G�J͎k]4m�Χ�@�2�cU����"ʌu�$o�e�ܟK9ӕT%*ቫ�&#m����Ӹ\�efo:^�����5u�b��)Iͷ�M9����+k��Ѭ{�1*����M�O�'������V�=��f�z�S�2�t��b?��(]�F��+�x��XB�%�`:��B�ʺ��Eaۿ�(�Rö�L٠n�ҖC��.avkV��Ѹ/%ܢ�Ȩ��e�H��#C)�ʖ�(���i�lبԧ,�������xM;�6Mݳ(4%(;sq8��� �3��e��Nv���q�(�'YYm޶ZL6ie��d�N�-X�j�x�M��/�y[����oC�0�Xl���_�K">���~��d|�R�����oO��+��,v����o�A�{�ޫ��n����������q;��wk�$򹹧��/�-���~v�ݺ(WK~{p�FC^AF�]�//.�r4;��ݼ�B���oCDo�$�Bb���%Gezm�gv�,Xw��sv?���2s��FS�vb��?��0��\���S�:L��I�c��!��:����>��=,y��WW&|���-�(��#|ʜ��j�W:Yݝm�x�GD=j{_�Z<fCE0ګ��"��9���L�	ț4���EtaOh[��۪XV�_a��	�z�!����R�3����IHT��mr�YJ���(՛ުg��yor��P�jC�|�q|�d/�s�W����gpsC�z�W�XH��Jj�o�__���_T�K�d����<�N��,lx���.�d��27:�����q����Lf�@QQ���Lj�V��l֍�yuQ��Rx��E��6c�f�4ic�D=����ӝ̯9�*�=����^�.�@��Ⱦ���*e)+յtvwj�wtb���̦��OZ�D��ǐ-jK���Ne�y[�Ǖ�C ~�19�����5��b���_b��V�Q�٪�P�dkLN}�5���ȃ�t��B�
�>��¦(AHՇ�ם<�te��]^R��Z������v�Z��Y4�i|Mg����Y�6oR��pY��kd
�9��y�s"LI��c�n�-��P�ɎU���%��L���_l���?��n�����U�T�0.��vm�)P��]��5=+I�[�zO���H���௺��죆�����,I�����dH��8�Ջj�,����Q���}�r���0?e�aa�]uie]]
*�T���'/
���j,���=�'K�ע��T��0���t����/�9/�k�x�����p���`�$s��~Brݡ3l��X��ux����_��)9Rh��Po��*�vΓgb1����]�h���Ԝ�;M�#d��<�"x����z,k����*���ԓ��Q�����p�.6:f#'\����E�:�<>o#7.�R7�F��u�q�"e�X_l�64�;r�=w�狵{�}��r��0�q���z�7�W�w��G���� V*�%~G$ľB�g]Kf�� u������i�5C �/l4��E�D�F��jj�oN����V���齮��G-���؆1���	�S�v�ӢO9���=f����7,n�o;t2A��1��j���oyU~P��0�� ���������K�� e�����p�=���C�G*��pdXS���8𙎯rU���V~zGtI:;�&펟wj7�?����C(y	�2��q��c��e�6������3)�Z-�0o*�K��F�f�v2ō
�mh��M)l���>��5����-�;�}�]�.�mA��gv��p#v��܉�!��<EUٻ�OK�踴�o�r鯻^Å8qom�<�tT�m�{'[rp_4��.Z�_s�9,Z�t�׽7B�IV��Wd��i���Դ�6����]yſc�b�
�gԻ(׻)"T���pP��pD�\�����w���\����q��r.���_�[�E�b���5�-��d���	�����n̎9��p�s�Ҷ���5r��4��f����o{!��&?w@��0�������]�S���J��j���J�#�bc����y��m,�n�X��h�'��`��,��37��v2�4�/�񳉻�����*���j�WK�h��4=����vk�Xu0q�D�l������S2��ٙC+~����T����ߖ|������z*�ͣ�7����7T�I}5v͗�sy'�[���F�Y���"Z��}���c��i��,�q�=�]��,���5=V�䉑S��k� �Kf&���UA�s���f6֊l�ȡCb�e���ΡZ��BFA]ʔv[p�m�F����`�X��o<�3�O���7�V�O��9ՙHc���1&^�W��vv��ݮ��f�����]}��fJ*�c蒬����M��j�Ѭ�Z�"��k��m�Q'x�/�9z��(��&fy�kv�6��ǓVq�OuK�3�}f�\��l�v��;�H�:P�Qr��S��z��K�iy/w�'o׊6u�%�u��WVt?Li��w���p�v��=Qk��&���#�5�[�g�3m��;�:#%^�2���KL޿P9ڔU�e'�Ή�ڍ��<��t�8�>7�R,�QI����(	?_�~�OE� %��:_.J"���泳�u+6�����d�[ӴN�r���|��I-v��k;�d}�v:py��X���g�I�*W������,s�7Ì�hv�*��=(�N�n��f��N��f�w�Vj��#�~6dCF�+�ff������WV�@��p�)��h��e��"d��k$LN�¸""
����-u��婋����.�j0��E/���y�h���e,,�A�J�c���4�̐TȌrp����'$|E �d�Z�L\� �1��!���ge�&3*Օrcȩ���*7X1�%˰،^]AY0�Ln�t���,�wC P\$�J�Ȑx��R�
�X��[ж�J��-�yY*c�
�N�to2�L����yn����!y���'(�Y���U4��e���Y���Om���+���Ю�YGy�"��`E�g.�����%P���a�U�I�Ө�;n���wE~�Ɵw���Fs޹��Ourď��+ߋ�S�ݖ�+���F�\�ss����X%���H�k����Q��E�*�;n�o=�-�8�b�X�s\�-�����$�`�X�q�eH���q\Z؄%��t�t2�a�ŝ�(Aa���{�<���
`���ɝΏ���k�'�'�����`ݺ,+�>cy�>�O��a���EaۣՈ�3��	=RO�t��[|��wB�Z���I�R�V?w*X��D���}��O!'��U�V9�]$�7G��~�u|�k�ۿ����^F�ڗ�g�v��6��	�uK�#6��7ԏNYs�i|��L��1f��U�]X�5=K�&���N�䍰�,#ug.ݑ���pi¶^j}j��'�c�r���QޡF��U)�P:8���S�*v�9���E���
��>^��H���4��A�ܸ����*mV\�xsv��mwH%Ʃ���P��N-�d'���=~F��0}t�'��=��(��>��5��d��y�7�W+}T;�~��-�<�e?&+"�X����r�SDlco/-1pu��E��v�ރ[���s~�����)���N�4�Z�����K��e�1�1�3/xc9�3����ֽ������[U��Q����ݧ�$�#�O��|z|�抗Sx��ۮ�ʓ5��^�`K��*��V�O*�&VG��b��g���qu�nc	̗-�F��C�}�ן^�WU���;�fQS�������|��eӨ�!P���T;ϋ�b����������r�x�r�Y���2<φ�����B��9d�z}KVJ���Qf�.�:Bf�d���MK���q���<$�v�+�����{�2����kҹ��W#����Z����ܽ��-x�=���f�[��v�<][��2�ڗT��m6K�AM#dRV*6t���/�y��{�WQN��O:�:4e�:V��P��7�E�v��
�����j��=��+1fwQ�����F��^�yg6�mdC���U����:@p}l�j��Ov�_ȳ��ܹҘ�V�T�x_�����r]�� ���0���<�G1�]v*�r�c�+D���lD�{��%�
���Qg"����Dg�w��d^�,{B���M�|��خ �J��J�s#ŧv��<���;�����gj:a���JGT�*�v��΃cI·	Y����%`M�'U��Q��x�r�8(�)ܥP�f��n���ڏ�:�O���z;��ٰ�0�Gk���N��Y.�*��&�|�ޅy��۱���=w�Ί.���^j�ϕ���f��`����f��{�	�՞v9�R�l�2�`S��3�[έm�W�Ԯ15u%��^���ԃ:�~�h"��'���a�+mG�a��ӎX㵠%�zƵ�Ѧ�,[r��'H�d	M���r{�q���R��͹!�sr�Lq""L�7�ӏ�3H��6����m���C)�z���ᨅ%�ޟ7w���[[z���֚7}]�ߖ/��WZ״��n7�2���EoQ���zv�,O�Atf�`�`T�F;	�,�j�&"H�j��>�[8q�p!�NWq���,�w]ƞw� QG�b��ۇ�9��s����>A�hB�}�*��'}�E� �ڪ����3�.�*�;�Z�{�C-nV���J��:/g-]�����w��B��}���i��V�
:Gcj�2��fЄYz��;����
���}W���*{��ת�!�i��8(�Z[����I\�/�����eI�u�r����]��,noq���T��3���'7����g����)�tI�#*��?s��Q�C�<K�ezkt��P`�2��s�l"nO�7zb��r:~HL�!>�]����c�Q��S0���^M�w��W=+����y�ѝjc��!�&�\��~�rx��v"��]�j�DZ�Okh{}���l�F������)��e��� ON[��.��z�|7,��7Qs�j�Y)[º�]!sYW7&�@�"s���2	��QU��0�Y�,�g�jj*@6`*2���������2�L����g=k�-=+�OE��oD��7�h��2j��n��-��i�E]��J��e[*���[V��.��f�
���h{��AU�u��*Wpm^��n���T^��[N|E���S�|ј��WS`��/���	���^Q����x3Q$G�������p�<ܰ��Ҹ7vS�^o+�8���3�j�7(LB��"r�| �h�M�幊�9+���Rt��4��dĐ�%�r��)�q�;/�3�_X�����I,'@D�(+�u�7+��D�9R�hL����V${���*�Oٴx��:}9L��t��A�*����M�I�U�3��f��ڋ�`����w_'spKw�2�	ʵ�/��\Xy�j�ُ#���J���ӃDf=�/��]![���F�\f[u�Әz�}[X��
x���n��x_b����T�RL��NiGصi��_�Mw]��@��NJ���A<���w�-����kS����l�ɰtwõ_-��/�}��$�|7��$��$���Y���.^h����t��������dϕu�f+e_Ŧ(����`b��h���(e��^y<��p������X�wF��yo6��뻽ί��/���쓛y�^o����s�њ���{���.so+˽�.w~=o�]������o�y����+�:�o������m�{�@H�h�1���)-Z��ָ��ͩNӬ��Uw�ǫsQ���i�M�_�̾�b�w��)(�εQ:i�����S�h�Zqk�O+F7��[!z���!��y��ӑ�EX��CS��y9GQ�qH�"���T� �Z�
ʭ4��ܸ����!�3�sf��&���nb��ʟ��p��"[�Q���R��'�<��{�'^�ɌQ�_��Z��g�{�Ba9�Ѝf:�|^�ea����f��7�ੇԢ��J��T��7��]o%��u�d��{���'�:�]�����1���%��x��#�������{ Z�v�Da��������߈��{��@ƹ`ۆ?Z�!u�������U�����^�V9h�J�nw�s��W��d$C��Hj��o�i�ylL}f�w3b��@`Pof˜����;��\�/�L�v]�8�`F�>�7p�*�eU��i�2{S�+�B��H������m�ew��v�l�_[�9��vu��G�d0-����9e�K삦��#j-ކyT�\*zR�A���dU��49k-c������N��
�7g]+�uV]�n����ڑ���뭏9���z+,����to�+ޙau�Մ��+��Q��mt��
:vl��&w}VX�iQ�x٥V�Nq�c��i���{���BK�ܮorႚ��Ƭ8�3W��꓾�Bt���.��:諎��v���}igU��}͚ذU��y{�->ݣ��1��M�-�&;܌ۙf������������ȯ�p�~s�}�m9��@�f����E�c�S|Y��"��íf�{B	��O>�˛�>�n�V�k{�Ҕ�رုm�W=ق������Yݎi�N��w�'�}/���*��)�n��lh�2�w�S3���i�x��c�f;I�'D:��P�J�x���������`�K��.��\3��x�r��R����;��GxP�҃7Ksj5���i�1�O�Zm�-��i}��	<�5¶NN������Y���qK�ྡ��3�F���tg�+��U\ר--�Y�yp��d)\�-�V��Px���S��JK	א�e�1��rz��}b&sf���fnR�ݭ��];�r��{=��D�g��/l�ݑ���'.�{w��g(��ik�]��8Z��z�a�z���R FM1�������5��)F��I{Z|��wol9�?�2�%f��A$�_k����h�r���P�֢Ҏ���*��\�^꽧j���!aѝ����M��/�t��� [E��̼����fq
J ������d�wP��7ܨ��G��j���]���Z��a���;O�EZ��/�n��8M+G�������m��l�o��	�E5��	���m�ʜ����c�����&aKVƳ���|8�8�n����{��p��s~�v����Jxi��+���W��a�⎬��BO�Gn"�]~!]:wtc��y_�bFF;a�5jr⥢j$wX��e{�6k�w��Y?/�E��/,r~"U�w�\ ���ǰA�Ӱ#l0k�uB����3;;a��އ{�P���HJ,��'a��^`���*r61c��8s����Pƶw�c���	��}�"wM��^S���5Vk�����ԡ슞@_h��C�ˬ�/Y�G.�#J��{=~���H���Y�r��!�FJ���B���e�Fb�D��>߷�<�T�$�U���<7�(�2^����oM����!�@��7ϩn��4��]?:��~X��`�n�r��.i��8��]tZ+�|\0�������ɞ�Z����<�R�$��W���Q�^2�l��J<r�;�N�1��\���Ӕ�!2�jn�B�.����>Y�J�}o�(h��K�Wz_T��7�����z�#�|mn�JQ�ᇪa�lx�����:�.�V[��w��%a�	��_��?��9��ӑ\� 
ڶ���������=��E��Z�PP9����!�����S[W�\�Tp�����>�q��0���t (#�m�MZ��K���RV��LE(��ΊёUfhUh�����C�L@+�)� t#ll���(J��;�"
��
�A����'��ʻ��t?ۥ��_^߿~��'��$I$�!@02@�d�BdfI0��D�A�3"2�%0$%$�� H#�2H"DM)B ��$3M2L�@�(���$���������!&F�B0��(Ha!�$�"MHI�`�!�	Ld�&dQ""��e3����	?���_�����q Z�]t��b�Y,[��.߬���D�%�<8z�d�HFBD�L։4Җ6�B�*M0��H�J"&�1�e!���m6J32L�͓Ri�Q�	Db�I�%%���2l&�2��*i�L1��Ȕ��,�Q�RJA
H���Ƙ���6,H�"��H$lH4D�H�(�1����2I	!&���CF:(��~������� �p�]�UA@�� Ȫ�'�B��Kc���������'��>������D���s�Y=?��0��<�e���
��ҿ+��$��-���
�� }�F	��v��]��-�@J�W�Uz� c������N�H�:��{2�E�ȇ�?�2XEo��K�j�l�����
��""�>�J�\"*����/$��
,Q��j!V,{������W�!�������t��H5���Dڽ�䨂����gC�x�һ�B}�x���;��'C�\r�@���`���g�y���5�����Ty��	�D;3�_�/jv~V2\��a��p%A���^�O�Ϗ�}R�0� ��>GR����_#�;O1��� M�>^�!�>��m��bC�_yM�E,��?H��r�|�2R����`Q���͌%
�0�r~�"��d2�a0x͉�K�lY4��ޢb� ���2���� �ӂܜ,3j�h��D�g%�h5C����Y6�~� �(���=�'����	s�z��B C���Să�����Ó����;���ܶ���������@�;�P��O'ϙޟ �v�o����/��YB(('���i�;�	>+Tҧ���d��D��)"��� ���,V�m��m�j�ص����m�m���lUV�P� EBEE$"�#e���ݱ���D`��9?@��|�b��+c�����Q!d���ܰB���Q����g�n``Ϙ;�>��O���X4�� �tQ��̢
(k��>��)D� (.� �,�ֽW2���(�a�u����:Q�Nk�c ]��z�^�,UA@�C>e����
�O_��>gs��=��(�<!�H�����Hd1�d)��5ou��k`�B����(Ϟ��:�]��BB����