BZh91AY&SY_`��ա_�`pg���gߠ����    b8��  >�_lU��)�kZ�֨U �J�[i�ٶ5m���f�����*����YR�m����-j�[5FZ�Ze�Ś�ZJW�v�U�������L�*�����l՛Z�E��[0UkZ�k*�R�aE��T�Y�I4ʆچ�V��m�Ue�h�1�v�jk6٭�m�յ��j��T��kFͭ�5,��L��5m��iJjIim��l�ͱ[[&l[Q���KfM(��Y-��*��eRfm�5�մ�-�`��V�y���j�t:	��e��f���ٺ�])�٨�ݶ�����@u�I���kbTR�msl�j��������[2o��{��
��m�ף]3wt������ҷb����*k�kL�V�ڔW�T��9��Q�lw��mw���ogT�.og�[5�ۻ�8�S#^ޭ��m��z^�ū&�J�kVɵ��$��� ����SJ��]��{ﶃ_lݒ�W�ݥV��p���t�^�D��4�Yܼ�{c��t7��ｏ�n�]u��{�o���禙珞�_m�uJ��7ןU�ݚkGǽ�V*[j��3e2diC� �]���P�R��sճЮ�ex�g=�Ҩ���a���ۮ��V�mӥK��ם-���Ҷ���t���Ҟ�^��NULy����{����Zk�v�v�[ZSel�j��m�i��� ��+譱��;һl�׃��j������zhPR����R�;�[�R�����];���[���喳m�z:{�u�k��w�]�����]��z��t���$@4�M��5���m� 7�o�����y�u�����:{���)��\S��n�v��m�:iUZt/Q��j���s�'�ܽ���R����/u�T��o��޴�4y�a��V����H�b�Y*�Vke�ٱ�V!�  ���(�[����:���<k�zҔ)s�=�JwoA^�{���t�;����v�i��4�I짖�\<�=�ԩ����@( c��Ԫ)jm����2�� ׂ�U�v� t���Gwa�@t>��[w�@ �U͸���ۀ�WA�=�:u�y� �Wz
 <w�[(��m(�
d� ��
���h ܪ��\�\ i���� 	������A]ZL(n��� ܺ� �wt��Ƙ�4T�eMe���| �����]u,� jt���U��p=��;�W���w���C������g����J�j��ѽv���        � ʒ�Q�      )�4b��� �     ���d)���� �h 0�� ���J�S�2b2i��0�M42B&� *�{I F	��&���a	H��#D4��I�<I�����0�d���>*����!�G����~Pkƻ����̯-5�,y�^�=����Ey�{�B����@D>�TW�x~�@TW�S�?�� ��?}������G�����O�G�� ���UU��E�%E��EDW�ׅ�!
���EG�"�����!@����$A B
���P?HJ"�	QA(���U�J��_A*�$}"���Q����G�!S�B�������B�	D_A
��$E}���E�'�J�z	E���@�(��A�H���A��� <�
'��P=*/��E� }*���A���  ����� � ���T= /��E��=� ���Q���AS�J��C�J�P�'��=�� OA*z	�J��C��A*��J�����|���!OA _A(���A��_I�G�<��=s�������8���H�3��1��vE�^<����O����ݖ�p<Bm��+mjދm�nGY�����,��X�3�-����\�;�����Q-a�Ȱ�����!!����!OI��`�8h��MѸʡ[Bz���X�Y�$�r��������Ê����OB��%ի{cb?�n�UT��@�4O�.єܲ�Qi�v��&�&ç4
7g���KB�'~G�wt�Hf�6���p��Y+g�tF �2J�"`mf+� �ܗk!�4"����KVR�ff�\8�������e��{[����%~�cR˷ �����ON�v����օH�-��(7	3-PV-)��j�$oC�	%��ˆ%6��#*�u6���Y���(ޑ��s7v�Tj�4)K �b��T���gTb���3���nU�pU����Y���͌��l5���-x2��(�6$h��F#w�2<�.d�/UCWqn�Q�	,#J��vh=܏�GZW(�14DDb�$��ql"��&�l*�#��L�mܶյ32�#l�f�f�sk/@q���`H�����b�'�I<���&���;l�6!�x��Ǯ��%��iLY��Xo��d�xJ��!�qG���i����z�0^��6�Ô���UA�UY5I��E�I��@.�+.unn3/w�ŵ��j���\�>�Yw��I�]}�,D�Z�X��V��$��%���VUv���uk�-�	+�T�6?E��?����t�f<l^�똋�Qn^A6^~.���b�ޓ��2IJ��׬++���T�|�ZZU�Fn1�O��ëewM衸.\�B��Uyǐ!�(c��Ԍ�����ޗ.ݢ� ���C�����z⧐��&�Y�	�ȋ��2F%H�e[5�� -R��m,a�K;t�זQ�6��/�k2b����s-9�`փB�ɂ��B����r��ś6�vr3 �5[{M�lR��X�t���j��Zt�4Z��ͱD�X��"��6M[�V���Ou�;e��2�Jf�*�4L۶�q��X�T&Z��m�HfJq֡����'kp�3E�r���4^i;�~Lm�3[Wʖ���ӊm�o��e]jט�:ݛqG���I=�FX�0F1���y�V2���i��a�xoAh؟qU`p��@b[�e�9�Xh"�aIW�pQ���w�wQ:��RՌѐ��l;���ܒJ��� ���^B�d!y�(������iU.V-�I���BS4�b��%���E�;�Έ"l"�-Oim�e~���!�2sc�3*�v)�\��Z����d@�DI��U�����V�M�˧.l.�
T�Gf-(��jt�ytѹX��-c�(M�tӫ�j,YR�mF71��4E�b���+Y������"�_�fA�*�At�7SD��>;�oNb\(ڪ�U��wki� �̎�q*�	��E�0c(\m��3kJ�R%�?8�VA�!7�y��i�<r��(�����-�/LRR�����ˤ��q�!A�ͪ��stݔ4����Bh� ȉ�R{Z;�wi@����\��wq�{)��:r�k�JYwD ��{6��u�S$��h�Fo��NQ��T˦�顱~��틦M`n��(P�0l���@���(�ǖw,QX�2�Qe�6��f���d?�@��*�Ǥ�OT����ى~n]\Р��ީ����V�7�zkZMḰ%���65�)Y����u���64,���R���
��Է��(bVFJ�Qn�Ԩ{
Ȧԃc�x�ho�"\;@<+5hCl�o�v�XGi����%]�ەJ���n4K
4~[W&�u���('+Q1���Pe�7nK�)h�B4��m��kj\��¯0��5
Th�8�	c �3 ZT��/Q���7����ە���ᵉ�m]Z��H��(u�=���:�v��/p!V۠7w �U���$��ayRB�(k���V�?����V����e��i������r]�8�6����U(e��m(B	"�H�r�n`H��b�BQĻ�M��K�u��1��O]Y����#�T��5ӭ��8V�e�@�UT�"iQl��jEZ�Q�hfmd�ˤ�^]� 3C%ݜn�i�[�܇^ǌ���KB�sZzi��g�K?G�%�	7�{e��v��t����HY����5m����D���\�dmKi�����L�ׂJQ��s�km��h���/�q��+t���t�V���1���1%��"����xjՆ�4s^���sF�X��֥Y��*��S���XT���M�6�*�@��dV�N�a��E�K%�
�����9����Y��Z�j.� ��rK��_��QmZѫJeK�`v�ʆ*accW�;��`�ƃo�bK�u��g5ٹ٪�ؼm懈�����K2$��Qҙњ��	B啚�X2��yv-LгѫVe�J�-����n����Y�Y���1�:Ԛ,a�`z��Ǣ� ^�����u�*ݖ�R����/��6գ,�Cjܛ��Tt���qlݻ��Ltxq�v�heT�(�T���1,��u��ǁ�-u0+ʻ�)j���|�h�1���sL��6ZׄV[J��RLC�6bTb����0�������sv5���*���'���fK��܌/k������Yc�4���ۮ,�ū%Ў�^fc�s%�D�ٳ�G���E_���dPNŸ˼?��I���i�4��IN=���k�UR�Z�nj5w�C��â+���(�-ôՕ���m���l2��D�jL�dÄ"�x;b��]�:VL��(��5�Y�؇m֡]֚|^���P���N�B�V���7X�)�FK2���u㭸�����{���7��yw2)Z��t��u�<���p4���M��v��֯��⽳dZ�� 4[�	��e����1͇p�h4�l��q���2�Ƶ�j�H^A�W6n����l�t�9�*]� �/�#v���+��#�����/]����w�J5�~6���a���]�Bm��Ƅ_��[��=�QS�z��9<U��iOqЊ�r�M�Ǩ�~Ym���Xq�p�E��.é���q��ƆM"y���[Wիi�g1�yg/�]�d)Xf�MՒ�̣���_�,C������"U�j�X��6�xd��<t��O��Oso՘�k����T��]�Z�=�����x���Y'E-�ب64V4n� Y���dq�rZ�x���m\4��N�0�PN!�0�cY�3]!�f���K���6��MQz�0�dw�Ee�[ݗN�=7�l@���k,Ӭ �U�֌�܋ �"��W�
�y�a���� ݣ�R�����%(v�q�7eR1�v�T�+wC��n����p˘��/e�Nb�p��lf�V5���Kmn����h�=>�i�/C���g�5��۹,��QRD^f��L]�P2��r�ś$mh2�.*�vl��v���Z ۓ1�]ʁś�隒
d�h�rV3���nSW�3p�n[Ï(��Z���N��N��u+�9�M4l�t��h6֚<�[Y���
ܧ���W�~9�����ԣphkV��;�i(���]5kV��bׇf��[:��&�����eVAn����Jhj��{�j�Ɏ�!隔N5���M��\͂Ĉ�VA����)�Ll!Уf��WoYtJ�������)P)��}�f�����E+tN�b����n�[�~�$��H�Z�!ع%��c��	�:;�r����%n��v�vſƨ��ț���z�H2�\6q��^�¡���!�z�`rGX��d���mp� vWY�i��:�N���	Or6�̣Q�	r���Z��<@���r��0� ���շ*�6�E���{�p�u��ʊ�R�3�L�jk�^��H9KS����)�2Mr�Aoub�V��;��Ż%�^nikN,�mP�w0�'*��C*:d�[Y��VXu�re��	�AOuKx�\��D
r�t�m\��c:�YU�R+�[�-�t��a�a��\�O 2L�Q��u��΋ݙ����5 ]5H�wx�@�B��/^f�n�^�r�em�6�c͉�B�n�Yiǻ�Z��љxFX4I���\[y�c6����NM�V���S��F�Z����z�j,e�Ln^�e��Ws���XI���wH#�.ƛ�d��� ����42��l��#3s@�J����m:)��1"�zퟐ��=k� �<�� 4�<)4��C��t�ɱ�n)�v�3n��pK[%�բ&�W���6�ި�kKL�p�e�>k��VK8M׶���rՃ��t�Zk%maL�]����R���^V,���Y�v��l���r�L�.��Ɩ0b�,nUi.�	�mV
����f��	p13sAY�.�&�v[��V���ј1뙃wTX��r�.���I!z3u�y��R��ٻ�*�5���T1=5{� � ��{A\T�wT�f�̕ŏ,S�"�,i��B�,�b01,Ô��l5qR;2�r��pډ��㊚��6�L)I�!х?ƫr���D���&�IfX*,DN"���݆%�%Y{YI�ޝ�pvh��,�Q�(Oס�y����J�Qj�C{E	�1n\�eۜ�VV�)c"��C��#OB|y�X���9Ss,�&)��`�_�zm�����+\ܱR��+5�i��:�r�ctZ�L^�'q���	`��kU��f�()L��*���t����� �.�<���x�;-�sj�OpC#�3&e3��HF�mb����0ø�`����J�±�'��P�ʹwD�eK�f��Ԑf=�B�S�J��ۡXAJe
��C[����B�A��/F�9����&��=��B�#B��uե*0j`o.9z�f���n�H��Jy%�*�^	N�8n\8���V�԰��-���~���,
��/Q���,�2K{�	��op�������O,�yC%u��p��x�k:�3Y�btN�i[n�aP'�+)^^�ʱR��MdZ�a�27�m�p^�/X�n�ûR�j�t5�&4���FԯŦ���1���Y����{V3N����kU�/�D�,p�t�#�*lR��P1�+�nXhR�����{mŕ����纳1�U�����s�H�[wdD��4��i��X� n�e��%�W[7��o&40�Q�VZ�Y�݄���r��hI.:Q��J!��t��^���_c�ƭ��Ej������0��'P*�L&�!R,,�0�ֻowHn"�鼀l�N���hv%ԥ9�YW2�^��n=1���`�w�z\�eh�%76�i��rF�4�9H�� ��!��H76C�vVڔ)=�C :������Xp��w���,�{�Gf7���3�L3A韲
�n�!j�.���D���U�*�Fc5Y���Q�AqZ1AI��B���wy�,U�x��C���ȼ/X��s��ף�Lz�b��c7nڄmd�lj��)�8�NiW�R`x+��WC(�YJ�EH�wN�+X֨���MLh��� `p43u�_�$n�� �FUL�5�8H�e\�a،��Fi;���Q�re�$~�!���^+ Z�ܬ����%١.�63�F˙�R2�]�*�jǃDZ.�������l�Hk�g)_2��]_i8��z�u�u����Y���4��ܭp��[Y�	)(�E�bJ�eG��Z)���;��dWUI����5�!3@ܘ�+ѯb���y��p�-m�ú�g�Y*H'^e��m"��e��M�c#R�l���vE�a�I=��ǋo\9��&It��9&̥v��H�䩅O�hmiYO�$���԰i|C��j�3�{eiA�2���r�{%���Z���F�X��ht�f`%]����]\�튒[	�&-�R��2L����!dʹ �y�su�r�[{q�r���F��4�	T�4٫��5��gu��nTp�����ݱ�N����Q�/]k��/�`�(m�7�q�F���!Q��EH.�m#Bl�$M�0��m͉^XJ��ոK	Z�J�ޜd�ئ��j�|�U����wK\��y����
��i��"ĩ!�k���a�F��x�6�jd�f�SE���v���+	Ք��i�*�7��qd#�a��Щ�ݺ�ɮܣ�"C!�����N���
�惇wBGi�"U�f���@�Mc�^�Z*���F�޶���@4�ƥ��h��2�l�8S��N��:�̏�����]�·O5e\� 3^��8�0�v���+��Mu��oec�wL�V�u��*�]\��g��fZxS�����e�W���������j�{m�3E�f)��E������x�۸R���\qM93lBӅR���C�K2Հm$F��e�K�sf�x�>嗫p�w��V��F".L�NZ�̢u7jj�d*��F�eK�a"rdKM�F��R��ʲ�ͫ.ZN#S]nBu-HMY�mAH !��w��92�:�Sʎ��MT5���]#����4!��'���B��r5�Ɉ��[P�պ��?��v]��q�ERⒻ�ćPIcTU���kumUL�uY�U�R��y���[N�)�$���/t@�-����,�#��w�&H�9���w�ۭ;��G���y����+h<{CN����W!h�/4J�x;@,s`��LV��,`�`O�V-���`f���x�㧌�+4���q�g_CFf /�H>��|0�}���X�`�`L��C�&��$*ɢKH���M��æ
30��j 1�E��V�PQ�V��]!�����4��vg��n@}�?���������F#A��6����vc�S���^ѓ$���W&�WB����$0p��������xχY��9�m���z>oM�n��5 e'Xח�9�,��y�&���z���ѡ�����έ T�LV�%��U�Q��Xx�wB�9O ��`w�vM��z�))��!�3���ܳ��p,�f�1�0����OS��s����R��լ��c;��q��F�H(1�G��M��oteɹyʻ8Esv����V}'bv�5�kf�w�B�a�Q�y:��v
���U��%yj"�Ü�չo�`�}�%s3h�c�N�a�@l��B�۾77���U+Z�h��	�vJ���YYJ��tb��{�S�)�ʇn��ubN�Zf��=}X��XZ�N򲢘^���Er�Y[d9���E�K;\r�I>9��%l����4��BN�D�V�Yݜ�ٵ�4�����=����Y絟��m��X�)!�1��c��#w923[��TX`�	Y�۽�ucB����L������W[Aj����ᴐ�x�ٷg��Rf�K�����f]#�����K�b�\U�7:AYx5Ħq�3-�b��	�!�s��aݬ?`N�14#u��Ē��=:1Y��c�Iu��b�i�l�7X^����������D���
�e����sAsn�֥��VD �عʐ�wN�ٚ+ �*�'�P0�.�]
wԅ�,�5(7����:4��fX��x�gDq�D�&�|D�Z����:�w(ذ��#��N9yC�ܝ)ǣ�Lb+u<ԑWw�hm�T�]F8��z\=��d��Vu�4f�jԿ)]Ri3�Ha��H~��)ed�g`�zSɼS��}�ev��}�����!��0c�8*�f�7n�r��b���ૹ#}P�S�(MN��+O;h�FW^>�`/)��	Ƕ/cwO)䘸��6J�B�ge�d��Wj&SrN�Xn鹮������
*0G(�v����5��A�"Q`W3R	�W8��]q�V�o���"�"h)�U\HȀ���]F>�Zح�z�wj3�o�=v�Z�̰�*Z����G���R��-��z��N���A�/��83�8��z�x�:�Ԧ+�3�lѤŷ]��e	��4ޱ׺�&�ԏ3�Y��Ɖڶ�wi�{o���B���Z�Y�4;���j�;;��
Wƅ8Y�3m'�k�6Xt'u�}בցP\{(��gt8S�7{aE��u)��|0�Dz��v
/�2��v �*?Y�[�%�<�tm�n�S�1��%foF�tY�S;ͭ}�20ރl����؇յ�J��1c�r�5k�[B��.�/n,�Pw@�:cEޕ�%�;�i�s���YX��pn]�O~����^�d�3;�h���L��-����T��ӏg;qc��e�k��	m-�-w���]�n���n*V+1�m�{�������UR�)��!9��gs�b�3H��k�]�9qgD�Q��Ӯ'�$��Ǘn����Q�lim)w��d������r���p�*9Ԃ=Ӧ>�}+q	y�G��W3FN�`�#ւ�p^��9�ʛ*#[��[�ӆ�$U�m$e����.l�M�u��a���ȳe�}���\/���\���F�ۡVlP��"��nf쮡6A:m��<�[��]]�ǃ|!�����1H��cAudP�ً2�:�K�"���kA&��{�
����uw���&Q�!=HM��d~��� ��H���\2�j�"v7��=���Q.�뒊��Oa�T2c�]��Gk�-�8��;YP�|2@�խ�D���G^��E���ܬ�JsN�1��f�)���-r[c]B.O�^ٙ OT��C��b2��Ԭ�!��q`�P�0oV`��lhϯf��O�T�[5�޷�tb��9f�܏�\x�]O���Y�˦빍F[���V�)�[���'���:���ɺw*�nbYB��򔈷s]�tmLx󙜮��'m:ȧPN"���N(+��j�Ll�X��f��ތ�4f�&5�5��:9R�!��7y$s7�7~8����7��9XC���y=�i]LCD�mm*������N�6�wS�X����N!�f�.����^r����8�"F;��i*�,���e!\�Т��8�tH��b�՘*�(�>z{)��k�`����*o���:����()8;:seepۻ��ep��Ć�uz�{dڍUS��,.�#����,%,�n!o�<3V��L,��+�mQ�)�m�����R��9�b]Ak^�9��#�g�Ut�c����3Η���w1�Pi>V�V/�g���-�0���F��z�&��I1PA16��a����^�D�E�_4�k���� ��G�]Z����rB�e�or�g���ެгQҮ�\i�.��@ˇ�\���1��,���s[O۫���u��V�Nk��n�ث���e�h 9+����[V�$T����c윬�~�2V�`���S�s�W2¸�[.AqP'�{ݐ��:5�Ŝ�μp�$�]�g��}�S�ty��@�J|&5��6�crnU=�|1Z�ʓ��CU\ꚁR�N�-7��_Ac�ܻ%1t��8K�[p;W���!�I>'�)��q�^6"��Pr�&��i��{�n�v�� ˍaP>�ݺLmw]�*�V�;5���N���z���gCPu�7ԐV��U;�%�I������bbZ0�r�0�ܑ:M�ݟ�W@)U��*�f�tb+��"�q����v#1V��1�c�\�*z�x���9J�a1u��L�Տ�'X���Tם�{AZ#�3�u�f]=�l�N��v
��{.��Q�w�pKM�}����&汇v>�b�"�;�>Y��(0I��+�4)���{�vݴ�� �DY�*@�x��v�L�
�G��^����
۩�_]q�˰�������ꇑ
aȹJ'wK,����f����1�rT	�.��단�3�CXG�2�@���w�$P&.`<�\�8{�}�qJǦ�<��l�h�u6ej���o����[m�V�Tw���p͙�'Ȕ�/���Z�a.�w�\ӣ��+*R��Wr)�K��l7��')k²XW�ꗫ�_.o)�j�ВŝC0�l}����� �$�V�T6f�U���tu�s�� X�z]���&�jr�o:��ɝ����K���r���E)�{�]���(\��uòG�cgVTrËe��<h�k�Ʀ�;X���U�ol�����n���:};����ks���N;���^��.8�q�34�-6;h݊b�7_S�,,z*�wS�6u[m�W���lE�6���u茫iB�5�k�ݙ�eE^�Jq��iV�[��n!|�"j�f&lX��׻,/ڑ9Φ#��K�Y�X#�.)·7��s,����#٭[c&��=���V���k�8��<���m\s��<�mF�a�YX�N�s�)�b�����| �z:��d͐��6�qr9�wY ��l�b"f�/�"^oڸ��o��/�{u����o��1E���.M�3O6{Y�\���N�Y�^�r�@3]o���K��]U��9C"L��+�94�b�!��d�26��/oM�҄����]॥-�����*!q��h)g1�-������Rd̒��su��4�P��+&r�/��;�z�p�j�� ��y�!�(鸷k^�ub����j2:�]o�q��9˗3�<�$�RR�NWp���R�>�^�v����)�Z
��j����GՙI�Mq^Gқj�;�u�����a�D�(%���<�b�C�{��_Q��N���qǹt�}�Y&6��N��"b�]K��!�==a��(���( ��1���15|P'�b@m�wGk{"j�b*ƚ��y���,�`B�ެ=�3���Q�]f{t��І������K/�AhQ��A�W	J��+�+4�YG!e��{zn<��O��6\��Y˺t�"vȳҖu0��=�R�v�R��$��n�(�h��y�P5	[G��7{��+�����2�zh[��%�u�AT}9e�MH��#��N��C�B�k{�N��΁)�s%:���O�@�6R�z�m�z+q�ms�)Wee;�̵�_U�8����a9����`t�����Z� ��޾�X�εn�f9��xg0{���Q�P�W�d1�+��u�<*�^�l�{x ���?�f# �Z��qi�'qJ?Ҷ�Au��M��.�W/lu>wQ�00�<׋�l��0�^� x*]˧}14�9td�����;��t���-�9�.��=us�������Şw!�i�{,<J���NM"޺����M����%Z�uyZ��ڴ����q�ğ,��# �z�rU��F�5�����XW��Ν�6z5MX�wEu�ə�6��]��p��Χ��LJ���<w�<�se��h����U����AU�0�k1�Y�g�q�V$ՖԼ�s����:T{�B��}�h�aU0	\S�:���ˮ
�����oUk��<U&tE
��oA��^�jl�tW�^e�['J��O
����:�sE�w����c��>��r�umFl�2Ze��F�ڲ���(�թ��E奱�#���2�Ay���;n:�Z��:�T֜mlU�M��b��R��@����m�j���IM�9i�Q8�gY�C˩w����t@�/�	���нӟxwǩs�g/�A^�=˨X�s�9���5��4���SN<y���s��J���B��ĺk�j� ��IE��m6oS廫0V!�5e>o$5)�j� l�~B{��a/M�ӛ��s�^�4XP:�p�[W�d�����j7xXg��F�7�Ӹ��**F�k["~nP����8�46*/^M��qe�٘.�O���i����󺜨� �����Py���V91Y;�W�6�wJu,����cm���7��k6�Gon�vu[6�AlN����[ʯot ���?��tbG^�i�l��y��w]�A��W)�� �&:�T����{Yn{`��D��Z4r"`�����������|7�69^M`X�ۜ�ٝ�:���9�YΣƯ����KW^�W/���؟3Й��خ�-�W{c����t�g_"��N �ὑ��ی���9�gd�[�#��ï���.խ��ɝ�n�ޣu&y�M�J��Y
�EkIm�hK����ٔvf:O�8&'ZCY�=J�:��[g��ݩ��E���a:�t�l��0��Y�"�Ӄ'W[Z���ƞr=ɑ��fq��p[{$꽂��֍�o+�CrS ��nQ&�V[�
�&'����e�v���3e�;�]��s�\�Cq`sPS_J�+�,m��n7���ZPC]'����^#��D��r�%^T<�3�RTސ�2��7S�6|���u�Kۣ;�F'iQ�f��Zj�z�r�\wX+Mk�ES�e�v��Gw#׊��=�
OR腼���j	[`��RȦ��{2��E�0�����]u�Ғf�n
���֢�1�Kbn�.�V������ue�-���9�ȵ�S����bpؓ���N�;�gQ6)�B)K��,��Ւv(Λ2�mVC���E	N��W1�O�ɈɎ���\jo��ec� �&�	ך��ܜFuBK���L�v�i��e!�����6���Y
x&�Y2e�)���%e�7y����l��k��/���'	��7�f[��EE40�3�u�s-��њ��f�=�%���mE��y�kre��PU���ӧf̠])�ZTf�`�R�Ț�X��*X*��� D /��q3�;\���q��{Lڏ�-��z��뷂���$s��0�S_� K������`c�w��]�0��.��9��4oghv�ȟ2l��a���q�
"��҆W_:���J.�2��('-ՆY�u
��q�0�e�<ӆf���]Y.��X��U���5��8q��z6٠��Ⳮ�P��+:�)4��0Vl
�!�14�)���i�$:��N�tʎrx�]#��!ȷ^&ڈ���)���е�i���6$��]��h�s#�ה��m6��UtϞA�����7i�`�.,�:	-uǱob�J(]�q#�0D "���E%u�AlwC1��\�oDu�q	���3o��	��֠�*R�	f�`���ֻn[-B�&S���eҬ6o��"8*��>�7�������6��a�P-���h���J;�wkSvV�]�˙�]s4�YN9�t Fų�9ta[2�Yݝ;����c��3��SV2ݷ�n�.�/�[������h�ӂ���{ph��l��s:���s2�+wa�t!B�x)ag�ڑqĆ
�ʼ�:�\=z�8p�S4�6���8���+]v1s-��'s?k��2��[��js���l��=n%����5D�p���x�S��ͧ�X�	\�U	ώ:#k�80�n�c3'Jf�؟�F+�7�K������RG	���m��Vr��5:�ڹ��4��f�*䁽U{ܗVոfAXj�V� �F�b�+F�T�}Gqd�>%x�z[mQ�kOo�:�$&9�0M�!ѹ����t�(շ��#5�Y�t��gi�*G��r�dٷ$��l�2V��
C�$�rJ���:�[ܸ̣K\|�z3���mD��:�n����s%�9V`.dhD�*��;�"�[�S���EnR�L6)�PoQoGxw����;��ϯ�&�[�ݻ͹$sj�C!��{��I$xm$�y#�]�
�m��D$F�s����o`<��ĭ�z�ׯ�Êvv^1X�A���'��D�A����QD �( BD���E
PI ��W+�Dx1��ˍrw#�8cR�U���vv���nR~m��&�\�n��Q_�������~[���ʧ��|��b����A��������3�����_٩P��.��`��շY}CXrڵX�٢VG��z5�[�Bͼ�U�w�XB��Wb6����:��B=���$�oΞ*��Im����[Ī��k9�}G!v,P�O�e���d;rTL�o6��]��u|�
���8�ڊ��q�BpA��z��4�k�� �3�L��b�7tm�Ӕ� X�m:�sOH�@l��l/3p�۩�S�9R'#�ַ�7����ȝ�9�����������6�7a��p�Ecy]v\�r�Usu��<��r�ص��ɽ�vʹ�J��;���R�o't�s�:գSK%~��D�.�q���"�{����6KpL��;�Guf��h\.�Hݬ?eMm9���`sM::Ō�����Z9�l�hsEDd99SW�����V,�%Z=Q�k����bPB�J��9(^�*����A[x1�M�T�A���3&S�x$y��tKWeK!=3:���:m��C`�H���r*]���M��kS�QJ<�1#�/c�۫�X�t�ڛ����*@����T�+��Tɜh+)�U���U�)H@0id̗�K��6�Q��)μ���Z��S��w��f���ofY����k�s�Mm�Y&]�r�#:�R��[��6�m�zew#���I]q���d��v��MMT��r�=�WhV�e�t����8M.�3;����X�����X�2>Fܮ�²<�B����8�e���o��u�S����3-�G>���z������sf��֐B~q��ű���l���s$ݱD*ǎ��[�i>���� $��aި+ub5Ƶ_`��^���_l9�38�FAY�)n�x�Ea��Ń]��q���n��Զ=;�'�A�HRէ=t� ]��!���6	������a�텋��#���ڶ�i=�i�Κ�!F��.3����h[��w��0��&\�r�<<<��Σ�	R�y��Q3�L@��v��۳��ÛA�m���Е����ʃڨ��i0�+|s7No�;&@r]hF�G���ڇ\gk74���*f�]Qӏ)m�\	w,��d��m�ficvV�H�������"���+Ш!�����eXo�j�ɥhW�����g�N��bn�V��j�a�r�;��⥗��3k�ȹs������3��k(0t(�<�쳰_͝�/^FuP��k��ţ��o�rT�d:f�`w*���{sw�[X��ު��qV>���.��v�7��b;l*�iv�v���[ےn�/���U,�#0ܐWQ�FPwc��hd�6=�7�Խ��0f4SaoSpQȴ@�48������3���HT�S۩6�%Dm,P��mAj�s6zWf��z�p���1$6�<F�f�u�=��
(le���흨�W���wNx{C��@��!VN�н���ٱ{���6�/��}il[wƏwe� ɴ�wZ�=ٕ�]2zs��sdj��Y۹�cW
�KP��:�A�i��en(�
�ۑ6�X��zg�G�υ�s���|ktN�rm���[fF�Mv�	yRhҺJa�X2m�p�Ś��u!Ô�X8��"����;�sy���;:"���C*9c�\�ֻ+�YY;6w���T�u��gE=g����*��X�v8M�kz�)sgV�� �-Qu"��K�wͅr������U��2u��9�{�.瘹��*.���3T�����R:�\���+��*\�J6�{��|-��=��$-���e#��L�׷�4�*9pܖ�<�b7@V<똙�/��j`��x��| k�Q<�oI9���|P2��I�����֤�j�F���|7H�|��c�p5d,��l��3�����Ԅ�Y��[8��z��-�݊uuL>k']��({T��6��.iɕ��Ɨ�e,p�Cy��e	%�!$�l(Iփ|n<춡=z���w��j�E���d&��x�͌�4�+wV�L�%{�uuMr�SO^~Ք��c6-��gz�h
G%p�^��+ U��1�6�a��u#H��h�6���C#�=�#�Q�w����am]yY�=��AJX��	��:��K�+iUuT��iݐ��˚�m$o*�WJ�VcsW�����]�|)|�bi0n�M���	R�8� ��Y��S:��Z)�$8�[���+��.�ٗד�Ek��/F�X��Ӿ�4�ւ���������<腈��7(��%m�)M�B\�쬦��2�t����;Z���Jd@�&�\�Er�qvT�,k�WpDs���gs4�Oʷ��-(裷3�fT��N��)��ܝ�ne2OH(ۜ�*�s=0V�\u�գ��;�Γ)��l���xVѱ{r���H�փ����)Y���SK��kn�Aʂ:[���9v�L�.���9����uH�i��7�mYKVM�ocC]'��AB�%�л����;�J ��K�;N�\�Ω{��D"me�����E��w�R蔛K#u�:>�Ziu�%gG@Ȯ^��������%��8�¸Z�Ǘ3w9�+�Վ���\#��LNʖ�zKb�k�<fq.�̋O	o�%�K6�Q\򹙌��ɪn��hW�0\��;b� :�����]��w'\�<4K�L�]�4q	�o)��$Tͭ���LzxZ��8ftb�R�5���Up;���N˕����n'�f�*�`DH�\Ww4f\��aC0�+eҼ爕X$�ia\&1fPv%Z㛆��,����KY��܎:��XmqJ�#�˼��d̐4�n�0��u����\�:��Rɝk����;ST��뾗��'�]���̩��U�ͣ1�v��0���)W\	J�`�3�S�Ci�v?��Ju��������)++��ˇrW �-�I��{��vlPGWZ�c;jւʻ� V�#Zf��u
�+A�[6�jYQûi��Ac\��X��ݱ��gKzJ9ei'���F�t���ދ��Kos��/��"<��2�ᔷ��#�%DRG"��z��nY4��6����k��¶𱵭�ژ1u������Kw�#xiÈ�p¥�n`"��5cJF���֌��ӦuYwGRƢ"+�,�qs��|I�&�J��p�h�%�fVЩM���Yw�N����8Z����4^vu��O9�]�[)>++{�0듲��"�WV>�p3�r&A�����uQޠ`r�b��<�`�����Ws�K_�@qZ}D'���4� �2�Ԏ9J�@���֘�n-�C#4�,�̠t�����W��p5�#��孇8Y?�3�u�7�O]�jZzy�D�eV�ىA����I�gZ��cقn�e�Y[�R��:�2�vl�o�:����.a���x,9Ap����2��v\��,u򁛜�9�va�ۥ�ws�ë.�8^3y����t�:DԳP���JЭ�雦NݛON\V%�:��8��| �B������/�L��
O6i�UR�!幇��8x�h�i��.�M���w+�a\�8�]Ck.�RH�'V���BwY�ݯ����0LB�%����:�v�[B��X�5�M3:벌6�*�8���w�/����S_ �<G v�]��|����Q�3NB�x���(��N!��n.��K�ng_�/*��AM�0d2	�/�^Nv�#�w�^�X�7a�/�D��s)4Zd��s�w�^h��K�{uҠ;)M��R�>,$c�J����D�P��p�:�����]˲�ԸfQ�)6�5YJW�Zn�� �dk�mE���V�(�ɶ���ve�[�S �L���:�T58Wt�v���;�k�FL��b-s���wvM�GV��Z���e�)o_T����f��F���M�tfeR.я�o@���7AhQ�4E3
r
��i����(rvR�O0�Z��#M����aGGU޼{�p���UG��npX�=�z��������sJVv���+�=,1;�θzmʂ!���h��ڸ���/dF MT��9F�M4�.66e�8Z��P/�oq���gC����,A�T˴u1�/�p������5L|��ϵ�N&5��$Lҽ�N˔��[2]h�vg.�57�2���(:����\š.�|���{��p�䨬2`��������fat�[V"�n�nN�1�r����/��y�x�f����P��g8�I�qͺw��h��yL�F�ig,��w�]B#��eN�N�M����k0�N����p�sS�ݽ�aT|h�/f�9�2ɤ^���?'�`ީ��&Y;phdՕ��]G�W�E|��Ū�Y��śj�R���|u���G��fQ9�w��hM�&_��{�F�%��Z���:�b�����T�33�YO8Q�N�ѽI:�:Ꜳ�G�pwys��d�������A�r��ZCB"�6���%����d�{�\7�7t����G�Ʌ�kUgV�ە���K(D�r#�++�Xn`�c�*rѱ?:%J�{E��og'��Y4-di=ʕk-*{�lcմ��(^釋̦�P^��*�(���%��ur:��p���"�'�����խ��:e�';��h�|�O�l82�D��P�]�pĭ������8[�l�@��ZA	w[�I��B��59���<�F1�&#�)�jPzT�3��`�ăUk]i2u�u8����/uK�*�殨� <�ك��ݻ����%`�������Wbgv��$C,�#��;�G��b������[��r��^4�������3w�EEǝe-g^��x��'U��}8�JX���,�+w�wÎV�HN�O�>���]�̺��d�0o>�U�[��¡3E����@�¡Zz`z�s/2d= ���*���:����2��=Y��Ԫ��Pp<䖞��+�G34�F���h��%7V��A���`�w���D��G5ǀW9���A�T!j��l�i^��M�mvv�ǒ�<�Q��68'G	�k&K-!�M5�����\�;sn�ɚ��N�:��T���E���ae���!ٽ���m0�]j�Gd(�lU���r\V��,�N����-�7Ie�I��
�Pq��7�u�$)t�w:���$^�<q[G]ӠN�'g@H\S��9Jz+�����tݰ-v�����(���F�]c�oR����`��h@���0�8�/��/ �p���z��r��4���Զ�u�K*�;fҥY4�3o:��V����U��Sw5=���w=�/�ҥ��.���'"cY������$���-�R�����Dܑm��>�Qz^֍��%&Cˡ�iؐ�A�iS��̗0`|;�NwqDyf!5��e�u\A'1�/C�sN���:^�gT}"Ј��&f`�.���JH��ݏS֞	�K����`Q�U%�T���Sm�9�3�jr�g+$c,y���w}��p�����6��ޱ�4ث�����ak ��Foh�Z�y5���o��t�}&�GW#��_r�+;}V$�\�o �l��MKv9䒰+A���p�_����f���
���۽aQ�r��g��Xq4�-&��iY�5Q����!�J��c�Eb�Զd��5�bv�x�N��ۖb\7�����;	5[.*�p�1[�,OMf�k���U�-�!;%�y(<����PSF�E��+��&�N��r��]���-��g`o���k���m��yR��\q\��Rv�Š��Z(����Io9kT�C�:s��m���vL��ڶ	ddˮ(�x�\�E ����"�nB�5{g�m>�����	�M�4ޭ������ҧD���v�g���.�D�*�N7��܃��A3�Ũܱ�m�-ɤ1Y�2�u�6� 7��]�mjW"��t��ý�9!G�9�k{�et�*b�6�ۨ%]S��]"=�%ҷ'�U��L�f~r�M���m
S4��Y�aV�X㺋�m򂺉�����}f����X;��T��e�U�'�!M�,�44f���v��x!f*�ka/�Y+1�=�����R���*���wʒ�S;獪2R9�@��Lf�:D�|�]�k�v��g�b��j�-ѳ�A�QTV��n���&C��k
�\Ѽu��q9ri����μ�ot������Ifoa;�1�:G�EhcRH3�^��c=�7$�KP"h}�N�Yr�;�J���д�%R9Fߵk��d���;(p}�bN��Wk�;:��ײ��iK���	���qxucw���M5�@?.�>m]��p�}Ke�5�'���1����e��L��}��fż�u��訖q����c�![J�\9cH%�w�ob�U$��ow;�QR�8r���+H�7X�G s��-�"��wiV"�NkG�3�sŖM.�/U*��*5���yMq�7eΤ)]���T�6�q��ɛ�|/�b�gZ�x�ܧj�F(�#lX�Yr��ڰ�L���p,\q"����ms�I[�s�߯�Z�C�k��f<}�:9��W+$\��,�Л�ł�4\�A��.VԷ4L��s������7�ո既�כD� ��2��X�,N�z��\wn�ĩ��6�& �.S������^�8Ue��WZZ�/vX�ܛF��P���>�zP��5x�v��4];�s�㖷GA��3VX���\��%˵�>�7��ܕ7!�n��sn��K���T�ݐb*�����F`�%��f���~�j���ھ[�h5�����Q3u��p�}�a�.r��!��ƕ������2%�e�u}a��`����fJFL���#4��6��C�v��틸���Be��k��"�~k9�bܱ1Mkҳ8^�A��vYUq�wQR�]J����f�!�{���ן� Q_�K��g����D>��X}a��>����=��}c��txo+���t���׈げV�	��z�;�[)����Ɵ��@����FN�%�6���wp��r�vZ�3z���#kv��q��t˅٭Z�`���W��bb�ʺ�gfh�ݤ�m��e.��ͨ�8cFVu��Ѕ[z�Q����!�����̸��Z�[���e�\[����q�(��0�:(�=ܕ"��x���Q!M�����)�w+�Igw(w�}��VB�Ό�(����6�<i�=�-B�L�n]N������ʆ�j���e�z�]X�Ce��*A�[�q%Ӑ�fcB�����:�y�`���A뫮W�r�ͽ�
I�$/�
͓oUEʏ��g�|�]�椧���D���G�}������#1��k�;��Yڪ6&e�xyK���R�[�,e[��Nj�1fI��s��6.��Ц9��p����xZuaGq��aX��cxk�B8��*ې�X���Қ}��J���Aߐ#\,��2Yp�ol��v�LF\1.�e>�C])�@�CZ ͬg�G5W��j3^�M�j�B@���!���*`�q�w���*�]f�r�\C��m,�(S9�s��έC\4�����Zt5co��noe*U-��p�0�{WR}��KZ��-LאX��1��^cMr��&t���]��c��CCh0��4ҡC������
�J��rF�NI��)�R��<J����Q�B�hCH� ����i:�I�JCG\��=O"�֊]F�-�Ĝ�ҕKJi�hy'JҔx���I܁��f�����J�	�c�Ws	@P��U��SI��<�=��x�JP�t=�u(�����PhN����94��
\��Z�ҴA�@�����BR=J@��C�pc��eT����LȨh������&>������'�hEwy��]������oe�]�]L��Fgʪ�6�s��T�j�W+8�|/$�Ϟ_CT3�`=\�'yOULzvq~%"�Nٯ!#'��[����~OݜW���pRǨi~�N�_��;��d�ꢸUg��T�ymS�c3ݼ�o]B2RW}�C^�S���j�jǻ���U�vA-w��X�� oA�L��x���*O�u�	��Sy�4����&����.��f���U8�.�h���*9
�|�y�[������{^�kd��U4�U��=h�:�?r�����i����(�8���>��1]'����r|I�����-�սW81u�|:{�:���}3R�bd���/g��w4���+��_i"�x�E�h�ߝf;��SF���w}�F�����9no��mE1醞22���N�_��Fį5��z���b�������?{�[�����c��#�˧�k3�bj�1�f��\�ֿ��+���̧WX���r�.�D���# ��kA��Z�-kj��Z���e��|b�cn�jr�]�܌�}�AF�49�$/���,�K�i��ɽ�m�0nݪ�w�Q�:�u�zi�ݒX$['V?���9���3��;W�S貂n]/AOf���5�Ϳ$���]��xGx����w�_��宆���FsC>�_@ǯ�����[��v��I~��<:��`�I7�z�����<9�X��Z>�߯����P#�o�q�<�v;���48�t�&F�B-��L�����m`^�~�����ɚ��=;i
Y��y<�/T=�E�ߪ����DZH�O�W�w��C���3��獜�Y��1���q�MOm�b_�>^�q�N�.����B����[M5���1uu|���=@a�۳�7H�m�l��}v�[�T�}�q[R%���%���p�n\{�O��{�z,/��=�c��c��o	���k�F{�w��9_������=�+��>^��S�ޯP�p3�]h鱆�M�gu=�l��1�ߋ�\^�6��[�>z��alov�5j����ԆM���:SM�Gg9�7����5�d����<��V���q��\ڄ��*�F����.�X|[��̕��d�kY�x�M�G�Z��g!tR=��}��I����m����n�u�ٝL�]���W�k���{t���Ƌ�̱���,��h1r�t��nl���)�+���E�/V�gԵ��\������~{B.^J�o�S&���^=v/��2����	ŏ�O�:Lqo���8�=��J�na�o����d���a{z��BMa㛜5m��8*���������i����~?{��Nk�m��;�Wn��^��cV�����~������J>��缗{�_z7�!�m)�t�[��p(��\�dɯ<y켞�Q��N��U���P;��C�Ly�q�o#}~uC"�S������;����@�t�s��C7���j� �3>$����4�cf4Y1_��؞3~M�u������>�2���������M�>��dT�u"�fR�ўa<`�T��ˬ�_hѧѓ����S�8���]��cAثM=}�b��;��9%�6��_z�'ON�\�J�҉0C����5:˂��YR'�:W�=e�d�S_* V{�S���*�����v�k���ζ��?�};71�ەi�DgiW�3�3�N�)V��g�[W�~cF�Q�[�;�_����@�3y���4x�3��k��1��u��l�t�A�o#No'���\��d�D�a^���z��t~!O�\�^����'3�ҽ�3ʻ��0sE����0����85gl�� K�ug�W�/(����*�{Ol���OG7�x���Ya1��u)�R~By��ND�j�]��z��^g�5��l��y��ݭ���-,ٺ`���g� O-{X�s�|O�:��Ւ�)t��iOH�c��f�;Qȯ`��0d��ͽ-S��?<i｜G���Q���3Y�c�����v�w��.0}I�a����{��_��� �% o��h5��L�fq����𳓦��>���5��ǎ��ڞ�~^��~�9�R� Z�}�a�;�6�xQ�2zm����.���}U�{�ů�#�����(�#ݷ�Mn�R�i�
�T��z�43l�c)I����&�ܱ֗e��o+�0TF �	�n��E�e^��'t�;�tvFt�0'�	��}�2���MU�	����)򬱫�sI��Vh يV�>�����t�Z��ؙ�&
?_[Փ�:��}���׽�B���Bϙ�#}Sr��o�C��ű���<J�^>Q̻,,���`�P��{"3e�hރ.n=,Ӄ"���!�muLY��uٴ�שI��5~ƈһ��v�T����EMvz�O����R~�~��xPc�A�������7�_xgX����&�1�5�M�ˎ�#;zGv�E���2F�;��6=�^���P�kѴs��Du��2	����X�t�S���z����wj*n��Ӳ7 �"��%�V@�Y�޵�m��3zkj_��q��3�����;��Y�ޒO0�<ƻwz��Et���%c/R7���eO_��>'�o�23�~e`����V^u4Q��)����#Md��񚋫i3�̀�Mr�/���;/�w���EI�����~����>o�{Q���&�:�����^۴����9�f!��@�<�`7w��7O������cx�"�~%Os4W�f�K|�-�� �V(&M�ѭL���0V�Z��@���QSד��e���k#*��shm�y_.A�Y��k���8M�#kEK ��0�:��v�EKTS'8o��1@ގ�,�7��Gn�o�`y����z�_P�CP_���p�{����G��{��Y������旬�^:4d~�L�V:�~���}&'���	=:�y����v7���ג�i~n���^��ߩi쫏�ŋ�����C������'�� =�p]��:�8��m�h���`x�F�����o	�n�9~�[��zcԥi��z���}GM�W�f�����r�z
{`m����`$])�:t���S����d9N���H}W�t�bc��_���g�g��_�e�<O��ѧ����'�8M�k��'��V^;�\��:G0�W\̖j�#�b����u��r5�f�cca�_D��#i��.�f����N�U�3:3���կi�ſ½���s�Gޮo((Oj��W�X?_�8��b|?�a�N��@�<�*��׽)[{E��=DV����3p>�9E������^��]у��d)�[��k2����d���ؠ�YH�É<��[tP�82+��0US͑�7��p��[1�\��8S����˘�v�.�M�FPO/6�8a�,�E��8�N�Z��F�a�0�S'h������m����}�s�j�v�<~��^3�笣�Gwv��iIg���U����i���+�ePÎ��c�����P��ƻ�)��ݼ�r��z&&'�z�A�zI�0w������ooԍ�f�![��������=�V���yꎀ��yǤx',4w�a����U�bj(o4�i��v�_��~-�G��&�?�������n���l憼���-�{.���Ӓ�Q/G��a��X�,�J{~E����+�����{�x�%gI6zT��|���곧Լ���t*�ʸ��٬�9�����x_�D�=~�)#m9�{����t���Y��]�_y���^��� -�˸�T�������Q�2o������l�f����/�o�_�9H۞':�z�xz�;����[ޖ��%���5J}b�^��z�#�}�Db�Z��q��/������rx��W�t���F�a
��6&g��^��f�D���9EL��Fͦ�ZͩĞq-��V��$&2���)���C��[�y|���@B��^�)�(�.����p��|!	έ^�@[�`��{ݴ��y�2W6\Ƿ�6��e/�Y0�W���י�������3�:���hB�D����B����������r�����e'Ҟ��fJڱ�X8����d/��lONW֍�UF@EuLϽ׺��LWw���z^��Ik�;�����U;@yj�T�mfm;F�9ч�Pf��ɟD�ϲ���Ԗ�%^�n���h��=��}��xi��M���c�E?���P�����<T~}�7G�K˕�\�_Nބsю����;Q6X솻�lc�OZG0��êEM]e�th�h��u8ks"�=��>{��S��W�����L�������y����o:��B�������'z�U�.�k��;�ha�q��k��u�M�H��9-o����#%
��7�A�{�z����f�����k}i�\J�>^�{��J�j��Tey������S�/8$:���輝i& _�SԾ���>ț���VJ\�BCKwԬ�戯�u'<B����X���;#h���88<H�%�Ь�q����
�ї���s;_d[M(�=6�_��>g.���:���K뼽LJ��q�Q�%Ҹ���;ۛ�Dg��"x^Z(�c��c�@�n�5���M.�����|�^ݲ:��{�wn�F�5)P����������$U���̹�ެ��=Ϝݓ�žL{|޹z�٩���V���Ə5Ǩq�z?v�^��W�`G�4��$��z�w���6@Y�-X{x�/K�|24�����������>���5m9�e��&���{_F�	���<x��t��R�L��{.�k������+���sPjݲ�H.y�oX�d�����g6P�����΃:z� 
aw����qY*G�h>���#�$d�H�Ѓ��}�k��A�)J�	iB=�AL{�<�;�ѣ��H��۴�Ѱ��7�]ھܬ5�S�I�sW�32V�;B���l�M��i$�L6�F�I}�5���/C���i�=�Q�a]�~2��l�����Y[�+0S1�?����ѧ�8O,B-��y�&5��Z"���v7l���p��/�Ch�nͅ�v(�k8\߮�9a
�:��$A��Q���7��v�j�l�x�	E\���7�E�me�҇G�잵]���^C��}��|�4�S���/|��0���ݺ���q���8O^�JN�K����z�����=�~�>�z���6�7;mƮ+�f�́��k�A;|���P�a����Փ|�ϧ�?������ڎ�s��݆���?	�R���2���26	�s&�;��CV���?o�^mON^��x��&����o]�:��y�����^�'>�ǽ!<��n'B4���_�4Mv��'���b�"�ȇ,ݛ��z��	�8��1�T�K���i%�۾=:��'V��us��c�9���+I�ߗ���u�r�Yd�`/�f_�4�F�����m���c�X��/��t���=��.F���ɏ�$����v�B�P�O�3����}�{��P @@o���y�~~ļ�\�M�4�}�䗄Cַ�u���w��a�n�۰h�~}/kϧ��/ ��d"*�t���-�5Aˢ\�����|��+��vk�9�}P�v7����Z���w�qJ\�ڊc����/�K˻n�%f���ʛ�E�̶�mfdD��a:�ۍ"j�����.�)����3��&�K�w(4�l�j�q=8�Nn�!��Mi��:�r��v�.�,�(�g^�uhdr�y����O�ۜ�;��ɸs��D��5]P�ğ(����dd\tt�I\�{´CFD̩�+���q�h��>`ef�8��K����;� ��
b�S�(�FT�p$t	zO	�����v�6���k���^(��.�s�@�Ɇ�-�"CY3�&�ǰԎ�) Wg^��sF� J�%����ю�m<��V8iӏ]Ƨh�}�J=��.����?db��7��!��"r�;!�n�D���RX��*��j��hk�2�YPb pg�99r#�;سf��y��K>��X+qV��a��5U�����0[Û*�m�9:��;@#�r4x�X�c��"�ҥt��"��c'7?a+=��tR��%k�u�cUs������At��9��j6,������7Z��E4��4Qpp!�}��e�����#�q�d:t��=ٓl�]9�N�jvmM�=B�q��5���˖�+�l��gȚ䓥բ��	���v8.66��9�������y���>N��%m8Z���3� ���"Æ�qXw�	��|�R[s�4V�y@g��P�5�lc#�
��v#�q�dJ���yA�^��귽z�C�o��1E�:l��B���u����z��lK�Jr�d�t,T	u�u�!Ԣ�RӦ&p[��ѧ
̃MȀ���b��8ȰL�B#i����cws"E�)Y�jN��������')�W`[R0���UɊr�#"7�_`���pjnPT��!�mm�
��r;f҆��J�I�n���k��g�V-$�7��8K������xS�asm[[V]ɖ��������Z#m�#O���3����S���@��$�GU���s��;�W:������qZ�ŽFrHv&<��F�[�|	��ᗇ% !�{V	���������S��j�u����w�7)
�p�w��f��,V�DN��w�7��9zuܫ�=��)��E�]AW�<8pda�y' �e��F�D�-�|-�O[���'+9��Ő�m��ۻ�Ni5�t^,� oQ�ٜ��!ԑ�]�¬�����U�Va7ϑ�}�1�z�Y��޾f���lwag&-D�[��֧Ҷ�^3OK�nF��g�D֮/9����R��s����7x����%�'�S��SPx#��q��6K}>,�w��J��ԫ�3]�S�V>b�e.�+��Z�^%�%I��#�g����s�G��ȗ8��%�vR�R*1�K�y 4��O����4�diCZ�l'�#�l�(S@���H�4R�:P�#AH�:���RSN�-�N�+AT�hJ�
4Prt\�i
�h��+I�t4�l1rp�ɡ<Iʹ-#���E�ґ��s�)@�J4�AA����Jp�P�Γ����nc�<O$�H�ѧ� �T	B�*i���2h�N�y{�u��vA�rLu��i-��*N��c�
qi�� �����:�v�U�-�h��.��P����9�����v���ˎt�1��!�é����eįz'�=���.u��� ]�~��C�����t�e߀(��P�����'b��<3d�͙ʎg����V^��)��ߋC|'rSP���fl��+�#��v6�l�ZE��������k��A4���S+-���-y�)B�Y�=5.���k�ӻ�P�7�Ӵ�*Pm�R�1��Y�qRW��o���l9ژ(���d�6qS�������+�]��ϼ��P�sn���7��u�|C��π}�خ�Dݧm�ft�t�b��~E�}��n��W]��%���ٝ���է'4��xYN�L ŨZ�M�L��e�T�<5�eс����m��n픹�S_8��3γ�cr�_
�m�<��n��\�q��D�s�Z滲����j�CeG-}����A���)[.�X��C8�y� ���J��TZ~:�Vr���������uv��ޛ�sQ��j�����`�O�С���s5�K;V�UL��TR������ϛ-�qu�T��b������0AR��7Pn�|�=�'�'��-3�|�3��}L��.�����LEt�dT��<�V�h��Ⱥ��x�y�Rѽ����S�;�.N��f�>.��]�1�joѱ���~�Ґǹ��Y�d�{�R��R�H��{��ש�3x]QZ���Ҟe�{�
{-R퐝c_s�V,WCv�lT�l�(:�[�)�hN�tt<`�����gMWv�5\��QP`�fK�tvK�Z� �t�q�HG�ׁ�۪�� fV�5����h�����!�=�}���^%t5�0�'�H��o<4k��KYD눲a�v_{���P��*�]�T�m�S����>���ͣ5��Gm~�Dc0��rB�6�%�b��\��8b��K�hK��!5�"���hFE��щ��ꂪ�z*0C�,���G|<����kӦ��/�w�xH�2��xcG�bPX�����e�����p\0� �\���l<���U\y�Nl;�c��yE��d���ބJuZ]V\y���.�7}cN}L8��ٞ����sP}Tu0~<;�����@��M?�&����_�s��jV�E�0P9�qs�X��u���W	M��W�e3�����3�����S�SЗ�qm�F�"۶��M�w�V�����
*g����]2{�D���q�%	\������}�3 �4���6��_�[t�P9T+y�u�,n�Z��tk�y;�H���aMCuK���\:`*-Q¤����k�]��YȨY6M+��WzV�q��m�h1��P긟hͫ�����/�<����&Pp�U+u�:|vU��亝F�P�{�;�����]��c-Ld}K�]�nS��|��e����o�Kz���P|���P���}_}tj��S��}?�tZ��O�MW>�C-==�t٢��|��j)>���uŹ�35����ŭ�\{7F'�g'��Uf�;�Vޏj��j�I�[e����VOQ����%:�S٥1%�Lt=Gg�B��D�S;�M��.�ͻR�H]������b�p�]Y ��&C4�)E�[�n��ب�[����D-c�;m���QL��*�k�ꡯζ<��-Ro|~�B/ܨb��H:5����`�����p�:H�aC�Jb�T�G=�<�^JV8�B��$�l��0���_u����=Y�$K<��y/;��(�.:ͪ�����[^C_��T��,Q�	J�ԙΰɽ�e�����KB�E�YБ�y�ܿvwҥ��K���P���8�������ҝx����ۦf��m=)����B�݃4��}��
���d����0�)1qV��P��yd��(z��f_��ou�����e�}���u��.�
o�'�����/.��F,x�y��rʴձ����}����qX���<k΄g���Q��tdD����̟XPjd\}6/��h8�N�$ݢy�8K�d��ap�����][�9����4��3=}�EU��j���Z�`��&���k��-2����a�% ��U�;v[٢}�az�c�{bТ���2egS�:A�(���Lw0u�Y-pRR;����yݏ��߀0��t��m҆�\�>���Ix��3��;�wI�\���a�%N�7Ln(�x԰vn�m�:�8�P��I��r���9�k܄����M�i���Z:|�%cfǝ;�pa�	��+�]�W��/ܩ�Sا��Z9�sa��^��k��9^]YQ�v�`c�"��{�3~����bP�,JXj��YP9����uj�v�܃�O1�rK(V>m'���NجǕ94��<2��ʈy�Ia�+6`_zYDt*��=�˕�ƀ�P��Zs��.�:����{��[^Cٵ.�~�O:IA�CC�B���;f@!�oP3���1j�h��.CkL+�}��,34"�wL��&e��b�lK2����!��y�Möd�L����g?�"	��WAܞ�A��9A�G%��bS�UJn�U�е'����aqfBݙ����:��7�%�U���ߧ��6Biq��=vq�.,RSۨ����-�s����k)�0�&C���вMu%��L�F�R�D'M^a���%�b�oga1B(�\���	tpR;_�uq�{]g����x�K�9F��S�����r��:zv��St;�l�u�/F��m���Tsm7�ilu�fS:�`ͭ�5�wݜ�4V�4j�_JQ&��O���~�Pcͻ�T��<��3����.���4�I�9������Hȱ��J�?�����bI��o��C��'�F�ͽ`T�l��V[R�c�6�-z���l�zgz�!�>�G��\<��do�'x����C��*�����U��_G�{e�cC�1���|��ԣ2���3ޓ��ȏW����,ސ�]�n{.Q�Vi�c�3�1�KGub�t#rF�aR��K�)��GdtW���Oz�kǁ:���'X??�w��M�Z�F8Qiޞ����[ʬ��.�ʇ�T0�Le���aw��)�|�3���3��j���}���ᰅ*b�G�̗��"�:�������Dz�����E����{ff�9^f	�ۉ�����������O��qH�Ի�滫���7��m��t�e�򬚿qA�����:���ݰ�͌�������%a�(�����tu�ot��z����@�[3�f�9�ͩ��%)�^�/k�r�o_�B��dϋG0���Q��l��R
{�������9K�� ��v��
C:h�Y6�YT�emk]ꝇ�����+)׌@���?rm4�S�}=���֧t�n��������/�U�ԫ{���<k4^�NWf��aq�.��x����t�S�v_WT`��-K���Jư�w2GX����sOs��jԘd�Kw�A�4Cc1�F�:��ۜ���S!9{��,�6���7ݎirُss�(�� 7��xx��tD����?4z�v�t<}����QI��JB��L�#OsR�`�T]�f®Â��a~��[k��{Zd�w޲5���\(r���J�����j�z�m�����v��W��9���c���s��i�wh���ř>h;;b����*-a�TX
"����Y��l�����t
�`���n�}@4F84%�sԹ���C�gFT��A�Bs~�2�����ί�x�B��lEe5��cn�A�Z;��hP#�T��+]\�M�y�n�nM��~|}�"�oR�r�4��Q��k��D�F��Ơ���l_yѹ�M���f7�J��̡y�{d��ӛ�EP%Ra�1O3��W�,��6jg�U�Vb���^�6�j�߁@�أ��<���Rd���Z(�3a2Qw_�����׈�~S3υF��K��pqI�Ќ�L�٦<ϩݧ��y�`��xP�6=�=�����u;׸�a�ş���^~w�3�.Lg�B��oצ���|� 9ķ�	���0�I�U��+!�������~`��w#�5��a��Zop��YV�8�x��f�ۃ�S�(���;�Mæe�?�����朷t�S���V��2MAC@��Ǔ	4zޭ�Ihwi��x�����S�cm�v7Ĳ��.�j��%�S:q��,�2T"�5�vJ�p�{�������W�sIQ�y���e��_V<kB�F���r�џҧX<=�'�X#�ۆ6K�Rn͋1���۬��sjv^�3ɜX.���,ؕ�)���V7������N�MR@���%ò�SdN�.�s8�m���Z�z��2���rc/EB��D�.��|�3n����k���h�;�W+�2��sq�b�F+��_���)����k��A�<��Qsa,t��^
�<�G�6	���o��-�x���Դ�\�!���m��Sk��Gg�־0�Z�-d��6!��#"��i��l���������ފ�u	_O�%^���q��7��;��ط9���Il�Euc��>��Q�ӈ9��'��*a}�oz�E��* �1?{�T�/�P�<�2�&W�xW?,֎��Ȕy�b	r��)�?`*}����b�c9��ޞ#���#�j.a�V-��黝��XTvZ��U���ۦ�Xf �&)��*Ru��1o��D��0Ur�,��s]z�Q�b�-Zb�aS&6s�B|�N(�v8ɇ�v�XX�&�%�x�[���QP���/ �i�ݢ���������R�f�G&6uIvi�H5���.*Q�%�2�Os�q�|�#~=$�k6g��aLhdKJh|���Ld<j��L�
	�.���ѳ������X�N��]�R�
�����dܛ�u� kX�o;���x��s;
�OVÿ>� x?m���e�9��4Ak�LB~j��s/�μ�0�P�(,ڄ�,�s���	��ϗp��R�_���<�fe;�*-j�i�r��׃1|k�����[�M�a)�țX[���Ь��f�L�G	y\ϩUSsw=�'������^MA�C�A����\���	�W��a��b۬aT��sW]C�,��ڝ{�qX���O�<�F}_��w� �����9�M��B#��'�g����8�J�W;Ɓ��qV�s�O�����g�����]Y��P���E��_����q�j}!6��垹�Lz��-Vę��13x4�:�y1)�(�3���}u�3q(ˢ���o@����Cyc�0��@�N��y�M�te�����;]��@7�VC����ˡcϊ��8�ٌ��91�[��O
=��.�>G����ylb0�%�������v��I��H����ʟ�g/�ߴ�T3��\bXo�Vl�.���ǂ#\���Do�K��u��>�8()�kB�2B���i,^�Fi�X�X����T�Ϻ�J�V��!�z�]�2lx��1H����y�υ�Q�w�)�L�ڢ:���oA��]�ϟ6��N����~�7P�:�%L}o�Ɔ3���o�w��
���L��k+��BM�qh�e����ޤ,�̒�Iu�W�|�V{�|�M�5�;;��8�d,=���_W�_}�{m`~y=[O���%0�2�v��s��m����Q}0*�\W��M˶:`]��<�уv���]h[L�c�e���i���0�*�1:��'ԧ��:-�_��x�-��\��Ԣ{;��Qw.��(Bn�d݅�=�EŹ�E>:�����t�+ZH8wZ]���]�U-��$\3��'��?�-gό�dS:���K���n����K��|FqL�]�^65cw����++���yu��C̮!$�{�L���TZ���m���(�g��MlrP��^Y���!Ai�.Q� N��4�w@�?>��N_�:%�|a��2��ԗc�#"�2�&�s��-�K+��>&�Z��K����@ր���Y���&"ֽ��3OUe�:�k��#	F���-����&���I�d*�<��r������3mq�ܶ��I\���>"�z���ό��}����1���߂���@�CC���^C;�ϭ�g�Yt/~���_#��	�l��f	�5¢�ٰ�����e��1�[+Ĵ�/��z�,�2>V�m���y��l�k�d�'�Y�	�5K�;�����v��T���ƪ���B3���t��9�nb���q�����Z�7��$M�B���9��_B)��s�V�<"�ܱy�^�e�{�WM��%�����M=y���x <<>o{�����x�q6��F�I�D������:2�>��xj�.տK)���h�;}_��>��� ����$c��+�䎃����&�#Y%*`��[_��ܷ���k�O��K��tq�121��^^)Ks�#<ͯEd���\
���3?����)�I�jt��
��{Uv�F��I�rSy}]��B�wT����1jO��YO�O�d�V�y�W���&F��Is3�(J̹������(!iݮ�@拫��1I�|�Si�l	m�
�/w	V6��34�[�얷+{�n�P�h��1N��'��mdph�k���B�N2�ҳ����j�s�9<��`IP��r���Z����r<�m�R�%���h�]z[Z�]E�Ĩ���.Q�=�,�N�p%AbA|�芖ź���t�e�Բ�4�ސ�!�]n��E�H���s���ֹ�:�Ch�:�GI���R��PS��Ñ�^���c��1�'i�h�A�?yP��]�y��793Q�DS�
*E5{�{�4'�WOc�c�ZN����d�\A�@�8 �,6C����;�&��y��{��rB���������$H���tu��K� ����s��6+�Ձ�G�C.���s�k_}چg\���K��r��e��Ā�<	�P�z:oe�-�|ohY{z���6�UU �����3�*���{$�Ep�X��;$�0����^閾�6)��F���W*�[I�"96Ӹ���w�'�KFV�|���jJ�6�5�8�
T;��L�"�1��q�H����3i-���Z���@���s���4U<��!�py�T5��3�xtUBz�q�,U��ޖ5�)�ZD�� `nAyY$��q̦�2*��:�;P����/���̂)�1obc�w��2��}�:�q�h���:�qF8��=6K�nœ̹LRie�}	6֠���p�yvB���l�u��t��f�gI�H�|��١+p��-V�p԰��t�f �Х�ܺ"���5�$�|j�f2�ӥ��[�l�4`X�"-�Ǩ��D�:��O�D�fU�����Tk*͋�U��L6���e��i�t��E|���ǹ�ô�Y)v���!�26���7֙L�GW�5mN4�z
�mS��l��
\qE1c��ٻ���k�η����}�P�w�Y/��jd�gn�p
��<4�֑',�t���@t(<�|c��|i(���v������eW���Q[�t�*�Q;|�i�;���04��v�q��w`�E�-#]�$' ͹M����D�+M��][���N)j��ɻ8-8��b���2*u��Uo�R	u~����{�o���ܡ����f�N��{�ZDk��D)�GWmm��G%tv�pP������2V�Fv˪��<�3z�^]a޶�j��u	vbu����ʍ���W�P�5�M�҇bŘ#2.A�op5��y��Vh=��4�k����A��-�1K�W���~,�ΩHc�[��n��2Z��bf�<��q�"k1Z�{���݌8��[���c'U�?$x3a^�1,I��D&�r�f����S$rټ��@^�y*�j��w�V�m�1�R�h�3!�V5�wf����)_, �/uhW�q^�j�on�%�H#�"��0#�e��Bp��`��,e<7;9XGl��Л�ۇU����B_G��l��Tr��k9��LW�]>�Ky�u�%基��_K��5��[Ŷ^��s M��L�����'ۑ�]uX���	ϭ4::�Q���٠_N�z:���*[���˫��[��)���3��l��f��ٗ���q�=�[�Øp�*eX��_o)+���z'b��ꭗ\�mV[�(A�mzL�6[���Ҷ��c�]7��T={����&��EYy�Z��������ѻK"[��gfqZ�[�JS4�GA����X��&E!}�9�A�����u֐�Zx��m=�Z�-�<����8��W-�7:JdU������hv�^»Mh��1���q�Y����ֹ̎(Q�h�ݫ�QL�D��#���`��	�(�m��.�w��w �45�$bذ]��5JPw[����w�$�C��"&	Е��*�2h�y'pt]`�N �4E{m\6�0w���@$伐:�E-tJlh�$K�i{���R�DA�8��`٪1��	�3��*��(��h���{�TA@Wv"�JV�
�JH��ht銩����T=�1/6�k�Jb������hb�8N�#ͪJ^��CJS�5T�:�T� x�Q�:h�=s+AABP�Z;٠�

Z@���ӊ�֖�hH���C����=�5T�ESQ@���214%P5BU-�EUQp����i���X�5�����y�Uo���f��>b�θa)ne�Ѵ�g;�t�N�=�
���<��4��L-�v7�o������m[?5G�A =����s�zi�K�?�=����
U�%��>��~a���<��п�|�\f���S?�pv��ۦhq���95V�Iݪ�䨋<bӉ�Z�Dp��wa��N7F�7^#A�L�<�]��T���vfT����D,cd���M^�`��u�h�a�ڬsPrslvx1���ypa}ǗvԾgI����
k�j��,��PLL/�E�z���}�d�c�vת�F�[�e����V�꡸�ߓ(����6�SW��3��`�{�YS��	%s�����E�d^3�7��#���^Jj���3k��"٤%u�9Mê�G�TO�{u�e�^j����Z���v��E�Qz��,��TL���A��$e�0k�����m6�s�*:S��I*�֖����׊�E;���T7�����a@-2��a�C׭t�~W3Q�aM`�����&	��d���k1޸av�Z��M�·3�Bko�U®B`ܲ��ܻ�kb����R�m�6�K޽��*�os�N�Y=[�tԝ�ȩ���B��ߠ��L�m�4{mV�n�2[�|�粬L�L�F�z���H+�������I��ｻ-uފ+f ���Ƈ�<���p�G���~�K��:��4	>��cc��o~t?4�WR�yb��R�5�|��L���8�ݫ���j3���ۊr�;6:Rǵx��;�K,����>n�sǞ�n�>�]{��
�A��3 =��W���C�a{���q��/N��K�L�q=	E�B�S$�o9D9�˫6�$����Gn-r��������3!K6�=��)���S.~�>�
��[kD�U&/��P��c����So$��E����:�5K��!��=xU�(���:y�ˏ)��aB�
9��_"���oNq7O��d������/��"��<���OB���Z�ae,��a b��}i�;y,�����8��5"��_~HB_�OO�#~\h!����Ggd�R�moT'�Q��ֽ����pl�}&��K����ſ]��M�����(h�WK|��k~^��g����3�+�hQ&V#;2���9�4ν��ZޘB�{��T��^��`�K�mx���FƯ
�TtN�Ǽ}��8�}� �&e�T�6��M]��Cq��%`�݌R��&���0ƺ6�vmztg|f#ڂɹ��}y�ɲͽ��RY��XnnVu^,�'Z�2^)	��J�����ètc:�hz�&������nG��M���f��	�����������r��(7X5�>�Y}�E|�~ .��,�:/�=��r]Gf9{ś�ڴ��_T�\�&�Z{C]�RZ�mc4
w��Vl����ut�n@f=gsa�J��,��U��)~�ދcQ>�9�{��\)�|[j��s-u]�R�t�������0s�����L���w^����M� ����(Uq�:�=��\�"%�c��@�5r,el�u��2�ս�G���	�l��H��]:���"��o~�<�<7�qF��z�lh�'@W�+5�����q�}�xs��/�<m��z�6^(��̉S�Gh{C���:W��m�*(�F�[�f�hNta��G��5e��J��g��}}�ٜ�[�t�rb�Wջ3	�Z�D�h�=�՟�N_xnx����樮A7���o �)��&���S,u��냽���~�Ŋ��X08͔�<�p_x|Gz�TӃ�;�t].T�ۘ�������*��2?T���u��b��|�3\����>�'�X-{eصJ[��7ax�es����Q^<'�p��:��d�g��^l����k�&�h��w��IeC܊�Z�fH˲����'	�D���t��0mO�a�޶�pd[��o�s�YzJ�j���8�!�Bc�@�����m��E��+y���&��Řm-1:����LO��nZ��ǿg��;�	�И�Z��(������&V�>��lR�Sr\�t+lA�b��<ԻFnt��=�jK�i��$0��q���燳X�y��\��i<�J����`��R�%L�r�m̛2Ьt��^Rge�U�L�ʭa�&�e��/v�]�M�}3Z���L��N֪��<�C�EnvD�O������  �f�`���JB�0��63ٹ��.J��Ih�Y^�y�3:�Ų]���@�n0i��]k�fT��܎�3��ųp�Q;f:Z����V�?����ox��x�l2��^��v�@�ƅ��[�]�����D>0^��JJ�O^�lt�M�&F2/�*gK�0,o�M'Z��it�5�A�F���!����f��l��	��J�-R�
����n'����e;h範���
�:�L;�@�'���hz����4!k�8��������N����Y���<U�UB������}
�sk6u�n'iIJ��Y�4����ӧ�œ���qR�MR��]c����W�=LS�m�z��	���e,
ޥW�.��y�WHN�xZ��Q��FgL 'Aj��"�{����Eth�&�
i���fO9ut�B�k�2j�Y6ߑ[v݁l�V(�xl�CA!���T�P��"w(��1�M*�+��%ٮ�@- ]bj��?��]j�O�1H�Ң��1ƺ�\��Q�N��Ә1[L:��n����mr��m{#�)�<��B.4Ī�|	E���#b�	�SO��'^�2z���G!�]��⢽X���n�T��->b�Geͨ])b;|�_*U.K:b��ՍK>gh_q��1GV��1]�(���ǭ�2�`�v�b:��[�-���"ɻ�cGٝ�W����I��ָ�n;�����l��7��� �4n����긿M|"���s���Q�P�o ���^.i�V�W�VwK�6�V�w���Y��u2s��u��:��P���1����#g\�%�ni��M��ۍ�SS��1�f�<-��; ,�C,2^��:�oosZ��m�k	�R��j�u�l#��\k���e���]r�ǬB�Iy;���'8�\���&0Yb5�ޞF��Ơ���W&���b�Կ�����_���;�QO/������`�I�����->Ϣ��f��5��Sg�x{��z��wu���LT"�^^b�.;PǤ�ƇX�&�8�Ȧڵ�=!�U�-��w��y�*�ˡ��D:D�9#ϧ�@����a�^r�-@���Vu^�ԵN�T�}6�#��|1�-A5p�4!������@���pd^]�JuZ�Z��ӎQ%-I!�	�[Kw��pp�\�`k���/�kB�_�q�3`d|푧��j��N@�ʙ��+,׺P�n}�����ʹk�%�JP���il�
��y��7�ݰ ��T��{��N~xX�K��:w2����j��|'}������'�<�q�����^8��]kw�N*����!���V�3��'g�>��/SZG�s��ƲA�n	,`�/�*nT
��y�:);�SH3uwn�}��n�ݼ!�6X�k�ʜ؝��x|��o{«�� �?"'�	�8�ӎ)������f_�B��t7��l�Ӑ�S�7P��n�7;+]dȡ��2�>? "=p۲*�E���ꎷ���aKT�{aP��K怖P��f{Y���Ncٜݳn���;N�U��H���Cpy�p�Nm��;��r������]��n�w������h^߉���%�h��mL�ް4�N5	t���=��X�.X�b6d�:C_7H���嬺&R~�T�q������/(m��[b�?!Fc9���X��{�h?fx:�<+`�v������(K��8�.�!D2�e��
�t�Y�~��,O�e��v/�ޣ����
��4��[Ixmx�S�by=��
�5)�|
*S#�tO6�
�o�G4;�ss�5//9}�{�@|��xg����5����y�݉�U_��\�<���bQ��C�^Il��Y������/&(�	L��5�LF�5zfs{s��2'=�R�w��
��6)4u㳊����LR��,-g�_͒��7YD~`��y�LƧ7�e1�E����܎-,���C����Lk%�ϳ঒>r��W6T�!��w%p��Yto#�W#9WE���D0@�%C�Q��6k\}6��v�AS�y�vO8��0ff+��N�Ȟ-]5^���car�F�"��RＨL����J�;��"*a�s��϶�����
D�)f�{ô��S)hʭB�r�j9����Tt�y�~U�ȃށ0u�j��ah�'��o;�>����3�ݹ�5ok�A��0��9��q�l��[<b����^D;kã"+�6jYdSΥۜ����/Uk78:�ŜV���3J�XCa�;Rʹ{�ʒM�[g����*W��M�ޡ4d��5�y�V�k�P�N��;��t9`	M�j�O9���Z�!�O[�϶��������*�ϼ�Y�E4����̈́b�u�_yr-֩&)X�Ҝq�Y���&�E��|7��th�8r~+�+4?Z����\�7P]J�Ҧ��ti=n����ap[ʸ}��:xg�������7œ� �{���s?*��oҚ�^�l!^�Ƚ�я;�˺UkY*Y?^)�]cث�	�U)3�p0�%aT8B�9h��!�P�;��ډw�:G��栬s�a#��e��S.s��ۨ,��=\��iO%<�Փ��:5��u���r��0.z�4_��#�"��%9`T�-�"oD�ǧ�h�D��Id׺_
����~|�)�B%�:s����'3����K��IȚ���ފ����³��yQN��R�zO�iPn-\��}��kc����RZ6���C]=�d��%�𢡊9���������=�'^�oS��;&_8����`�-�����.�!
�(��~�<����|s*��̊ȣ?��+�4t��1�`uh�>Vl��}�P�1i"�_4�Zi���r4B���{\���!�;s�� ����o妄�uuc������C��Q�c�7Ӑ�ч�y6m�E��݈���C�sJ�G�X��-�c�6*���wcV��eu�&��~�M��|���Z��%0��
+ܣ��ç-��.E���*�(�����q�qDr�$.��e�t���[/Le�Le�lu>�Q��>W^v��:�	l�c�3��ll�pu��%�ұkH�z�������2����N4�hH{�J���Xڮ�4�N��eՍ]�՛�/J�;3�r�5d�iu�F�aP���!F�v�3��C�13�|Q]�20]�r"n��;��WR;�[�ԯ�����nH��*���L�����͆p�i���v紛#5�����z�guD>���ji7������WZE�e����vg��|*�(�*�ۇ���}���͘��$�v�PCf�*fԖdPz���K�,*`B���/Ø{���f��}�Ui�!ŨQR+��/�O�Z��|�a����#���*`2c�ݢ
��bT�^��Ǧ�t�.U�-��0W[A�@��mpɀ6:L2����U�]��+�pP$�W�<.�k6�<�����μ����*�o4�ظm�{'K��U��"��")j�jV	Zi�W���z����|{���}{��Ռ3^�YR�⼔�mzK&�/ڶ�N�iL 'Hb�׃9�2/����+�)l���1z2E7e�R8���WT?tJ�0�&�Z�d�a,�m������9.O^��WU�ҖD��\�m�/"�7��i��z$j��|]��C���j��t���H�T-��������V�ٽ~x!y*��JR�ݗ*|��5�%aT�mn��1G0��+�X�K\��q��PN����e�w>�Ed��a�@��z;�����h��0����뼦���:��
K����)���=̟�$�î����@%�+��$�eA���-������w�Y���ݒ�h�O�zqKS +K˴�&q��xD����q�9 ��nv�Ϭ5����ی�ח{e��j����4�q���T�O=�E5�&^�r�4�(�e���!�'��@-ęӑ�u����D榤�.����\�/%�z�|�#���ʓ����Z���r��w�9��fU�f�5\WO$��'*�&�5*��yM�Z�.;PC[��7��GpcӉ��F�7
��{������ou���F��Z��Q�MwNd d9�l;���Ե`3P�c��tL �8qi��^=� '�h��9� �m��Wl�e6܆�5М�������>��e�WJ5z�4�G֋��x���smt��M�c3u�u�Q����~�P����(P�J
 �����ǿ����|T���Jy��w,��]|E
�P�.����	����3��l�(�a�Hб����.�4ALa[�`�P�*�qZЎ�B`�z�-��
Yg�]��c��Z.fpC�I���GZf��+U{{��i���+��_�hS�����H�z|2!c[��\�8����I�fT�8��������gx��_�w�����y���ty�EkR��/}L-#[$P��ά���H��K�N8��Ŵ����ȼ�q����tu�Ɩ�zmPf�����V��>3�J֎:K�C�mE���un�W6�B�T��A�<�J(��Yպ��m��}ʸ�z2b����R�Y���a{!�i����1�#���Y�Z��魣�7�I빰5	�-�|5�9St8��~�����u�N�}�����~��?�~�5�*�����ZS|u�>���77�#g��be'8��q���gTK��uE�X#"@�L�����,`��VZ2��±�3:��^2h�:�5�(��BN��SrT{x+7coh�lň~g�� d �( @���n_U� \qgEZU�Z��H��4�Xq�/b
�Vu���g�V�&���|ͪ��E��X�Й�ד ���|D�D�}G;��u���#�|!�����7���8���7>�Y0mr������N�lh����+o4a:o���t��&+��F�ӄ:��C�0S��VHYo�4�f]6U�Yh"1��O�l��nTzk����.�鹥�&t�u	���b\�.l}��K6t���[����B�koZ��H
�X��p<:���M�xJ�u+�':՜K�*�]�:�9V;�r�gvgXa:k{z��`
#y��T�KJT���E�� ]��!J�k��h�2A$�gs&H(���#��|m^=Rv
6�R�;2�}��pl�iQ4w%�.�Mf՞齚2�o��:~�����B���E�uWvYP�R�&:n��*҂��m�C5�q��ޜ�X[����̵y/ip��H*�m����q.�"�*�s��`@�O,�Ҽ��*.b�+��M�o�^���]��za�V**��l����s7n������M^�21gXCN���`7 Z�6;`�!W��t;��4�k�[��s�-�1C �d��ќ4<��OILl`�F5X��	�;���[q�[;�W��E�U�����˳.ӛvv�Ѹ�\ƉQ�urC��[��K2ڕ��KUܻPX�q�7\\]��g�}�d����\�Iޚ�[�ӗ�����5G:T�x�W#� r��	���׳y��mX���I�˻&j��%�oԱ-�tou��rT�+���<�n�l�5w8�����I]�D�/52tW]��庹�acUmN;-�y9��V�����p�m��[��=��&�E�B�Z�c��e�6`�!b�.��)t:ų%_9b���g siԳ�_ME�/:��c�{��M۱�O:�vܚӲR�	%�y�]����4���gm�O_Sy����u�v�ζ�Z�q�3gmk�o4ړ�Mَ�K���vc��2ݽ:���l&&�S�����c9�wEW�l�4���9���x�ѳA[��۵��ۙ�f#;9�(�f�1+q�M
݆f,�l}[I�+/[O 㛻-�링\o�dk����z��p^P�f!+�3N�쑣o�M�-����]��-5{�ۊZ��m4�T�yBT��P�t��kެ�jA��٤�R]E�[�v��AKym�u�|�ۍvRnQ2^1��8Y�0s�V���ʉPL�b�i�N�F"����w;mv��>xI�4q��5,y�i�ב��ѓ��(e#G�Ѷč���vo^8�dԙ��)���W��dt"�R"��n��Ж�Դb��3�����>�O7!э5<;1�s4n��N�n�+9��˧�Lǭ����"�ǣ����߷��ߎ��CA׃/��Q�x6���;�QH�:��Z�ESP�!CE�A@��1)��$KQ�i�^�u{�$T�U]N&'cc�Qr2�IM��UE4�RQBR�5T�DH̴�AQ�R�D0���ATSIM��Q4�U%s��z�TQ�&�������������/cH���j����TS��IT�DST1�������"h�C���(�(�$���9��mU%5QSQ����*���T�%P��1Qͪ"�����"i
"J&3��E5MD^6������H��Va�v\�[����e&TS4��ޢ{�mKAn��:�I��!2�;W&�L_9_�SEd͈���6K%���Q����1����]]��@�	O}w����u�]{���o7W��ȗ={S�ay=�m0���=�EJe��<�^*V8�$a.^�q_�k�eq37J�w�h�<�6�2��H욹�z���Ȫ�qf���9�\���M�IF��ۋD�L�`��S:j���c�f����"fs/���6.�Jm�p�YMvb��J�ZFU��8�\_�p�߆$<�=↊q���Ëk~G�)��N�YA�-Yp��2#�rq��pⱹ�F=Z�g�AUSkW��4,���`���/h��^L��x;*�b���ݽ���ʹ�,`��mL�8��1��q�gǡ&�x�yp�ͥݛ]['<__z17`˱���!
jt�.����{b���z��g��x���01�BUI��èv묥�eCS��i\�{��8�2�g���1���B	�=�GPb�%K�t$�^��m�r,&<�r�w�p�>�^m����?�Eb�uE�$���� � VU����7N��45nAc/3�Rypt:���+wi�SMPR'(oVC� ���th��p�+�++#��8S[۶>��g�{�e��*j�<��e�S�;��Z������������-;L
��Մ�q uv��f�6^�6�/+f1��/��iޮ�\��x�ۙsdᢵ�����mЙ�M��gW��k�}�>��o�Z�"��M�GvO���`0�mU₥cZ���HO4P�k$N={V3�G]@��4�������:�ܓ%[W	��N8^޲��׋.�8��Kq��\�s^��R��zjRg�w�����.��x���&��˪������H��&�h.��ÌBc�*�\�=�m���+P*/&9�v���TeAwu�f?����Ƈ�ܷ5�3�����j߇��|a^*�7v��oe�L��7�T��թ�+Ҥz�%���ڃ��	K��ptݣ &�v���i���'�㣺��}�f��k�/g)LlyGظ��9�uQ+�����@NgWb����vڹoA��]w5�KB����s;�Ff���Nf�;h�L�/���4�<�9���E�C?0؈M�e���K��\E��ޥ-k�j�[XĕCR�
(����>x��=�]#�<�9��cA`.�K��Ȋ���X�E�y��q��jyk�x��;x�Nw��b���5Z��-��h��3�z��9T6i�>]�p�U(s ��,�`ʺV�Dqq��KU�g��7_�J�,�������v�$'���ۊp@�a�U,щk��X�KJ���EVz�Ƹ��_Z��@px]%�YYC���-{9u�<��P��/�.�ٗ��/&V	���-Vk�I�һ��sd�ŢMLӏR��}+�]���}���<�;�n��NA�n+��t(����<�;W?z;�R��ַk��K�S������3t�6�$ו
&SC�`f���!�a�	���_F;c��T.1�sf������1
�P�}u�k���u� �?��N�
"ƶ�qD��??`�M�Z��ڊ�T;a�lg[��d�p�:���Wh|�����&��X��xBb!0p�pe��+���x�x�c�!?a)�>m�f8��
.���^�<�m����i�(A�}�Y�i��<�#tq��p���c�L������[>#g��3b6*��J�%�t��^�=�'�Z�ң5�V��g��}n*=�=ВD���_�����I?s1<�:�Q�LL��jA��E��dƔK��9T�`��k�E�9�ƽ�i�ڜ�P��\1ؔ	Yt]�JpX�9zb�7Q1��l�n9���q�62^�X{�����F5|7�b�o{Mi���������z����MR�?|hVv���� Ng"n�wZ8���p�c&�kI7&^�ǲ�1��)���0����3e�v֙�jǵ=�a��h�u��TY��TG��S��T	zb�r��1��9����{������V���8>��Udy��8��8�䁶���GLYS�V(3F�x�-�V7//t�H|�N�r������I�n�ׂ��Q��w�*�y�:X�Jv;r�˶�v	MP4�jv����p����^û���r��UW���u���%���	Ṥ�yv�v%R��"�3�OBѭ���6&;�ma���	�a�/�eoe�b�x�%K��З��ة�#�H��0e��.SJ{ �%���ZN�j�Kþ�K���왇��ԣZH�P3P}`�����΋�=k�i�\T���x���� ���N3��s��+c��z)O�|7��h'U �&�zT+�\hE]���᧷!^�~�|u�~@��vp.m{ʴ9�0�Uk׹Frԝ�b��V�K�W)9�aΣb���A2�$%NZ{+����NM+��;�1�2�^B��*�o�0u0�a�瘛�������~�ޚ�cu0/.B]��5�.�C�z�X�nZ5�N#�ˮN�SA7i}1W����D;=�~��x�3q��8|_��\�[4�u0ܦ��e�����fy�qdȽ�����t�x�mxk��)_V�hfһ��tC�	B�@��k���j��q�0�kzG;l��+�\�k�zᒑN�j��z��`�B�8aP����y�*�E^7,7���IpՎ�$���ߵ��e�O-K��,��h�q(i����_F�KÎesPm>r@�г-Z�yv�7ڭ�>g#�����C����7�jı)̳���Cw��ţqŔ��I�+�h�K����'uyՇZ$�߲��uk#��-4�SzZ0s���V^N�n����o>|�|cm'�هL�0४Sd󍎫|���C������;m�)5�������rۮ�v)>�-�{eV답�N�o!�u4[z=��q���3�v6��T��#�9��Geڥ܀��b�&��M�[8���am�נ���}��%�y�$/��--U7Np�].S˯K�e�mF���T��u`2�e��G����co𞗑�9�)�s�k3+7~�ϙxp�*�b���90��������K݉LS�T�G�9��$"���b��or�ˎ�����4��3^�����:��R�Υ�P�	��c�<��xd�krk�e��2��k��ѽO�d��1)�0�9��QL�>Zz�oW�#���*=�;8ؾ���m�S���gK�bȝ��aŢ�<�)�Z��a)�⽨d�= ]�/O͍�x�b��*=�z3f�\��_j�~[KZ�Z�oW�R]���PY�8>������A����.�N�O�M��������9��y����+��Q1z��S��|z�RZ�b����y7��eޑ���b,a��&�ܦB�zP�^�׻|��}������X{ˇ]�h���֎s���R4p�ӝ�o�����@y�;�@:w�L�0��*���@#���Gj�Z��n�A����.
.���m�F�+�k{]Y���xU{,�V���ȉ���Ի�a�5����3�g��\[25%���u��}�U��7t��?��)��Z��=��ؠExJ�.*k$��v�//)S�9N��:i��W�k5�ٽ�{�����Y5¾Y�Q��k���~!����[S�R�V�}��C�_����M]�:O�����F,n�IB��ޑ9@.��(�"9�s�83�Q�{冃���G���S14�X�;�����o��*���aBS'^˯������������=������vN���ν�uYa}C3Gx(Vb�漚�J�k⥓�(����8�Ү�Vy]�ĭ�v�u��һQ�O���Gyޚ����e�C@�[@ߺbK
�2�rS,���Sm�ec�Y9L�#2{1j���2I�Ki���Wţ��-z�!��!ߔ�r�%9`T�m��f�<���2���oK�j^�'�,�9�@|��n�,N�Ռ|_g�
�H��ѧ*��v�)�.���v�[�,�p|-y7!;��ş?2k(�2FB��2��K��֙� �g}�r鿽�ux5�jE�yR�T��ֻ<z5N�{�n�K�W�ҭV�� ���:;��Z������W�9EN��
�����cm�5:�g٣%�0F5fuh}�OK@p��A�6n �&n�/0@��;���[/n���vlC{+��{�&�0�T���NۋF��
��i���<����E������H�;4�qd�+͝J߁8���IJ�9�I�ǥC����@/����	g\�Լs��"s�t�����:ߖ5��e^�%���U-G l(�����z��\�m����)�[�9�����m<�!j�E<�,���n�[X�S���-K+��$�kP��.�O`��lD���9
�L�@�kP��v���ZG���2|ct�;��]O��P�u�a)�;�n����6�_~�f�-x����"v������1P|�ʀ�ls#9P�L�d_y�-t���T��
)9�1ˋ�մ0P��/F"�C	�u���ŗ�?�"�~��[�9�Y�]���t��}�A�t���vq�.��������q������L�)�^�j:ۇ�v���m:t�uZ�:���h��UKf�i��a�Y�/d���F�2=��r�k?;�U���90�P�zs���}�yl:���_�P��ARY��q-y�i�Jط�7$��l�k=�\f?���C]�b5�r�H)�����J籆d�j%�jW!���sc�I�K�Mn����P���|��aq����q�@ˉo�� ��ܽ��u[�<M��QΘEn���Sۉ��Ҩ�@�B�{�V�k.�w;U[���m��&��
r�04,�v���p��/��.����ca�*^g:>����i/�v�\+k������y���̮FP��wk�4z�W�o��u蘤��]Ĳ �5���#V逨�»9��w<�vR�v>1lA�����0:�z��X�Q��»����H��C+2�lt��v�Ș���G\ bv��%���/h,�a�D����� �Ä��o���i�1�7�������Ҩgi��nZ˄TS����H<��P�u7@����phb�wF�l:[7q�c�ڞs/��H��摳j)ڈ��U,�E��r1��ֹ	��Hw��Xnfi�>E�F���n|���lB'�*)/��D���C<1�{��ҟ�G2�ϛb���Mm���]�mz�P�w���df�VD9�Qѹ�Hq��'�F�Y��K���S�jp6dUo4(r�C>t��f�3<�y����L5��|u��̌eU-�FE7�jǜB�]�(��l̈́���O�9x%n�Rϔ��^�"�W���#�jEn!4T\VZdE/_�s�к��i�3b{N,�ښ����}z���'�Bܡ��1t�\d��1%��0^��t���$��~7Z��(����F!b%���2T^�[��7J�k�W{�����1{|/j�1^^w=�ȅ�~�|�~�4P�!������/u���IR����m�ϴ���B�5�������9F��xy��$%�ޓ�cz�Y��v���{��j�_߫��	'��䏧�[�K62�0�zw���M#5��]N�~X5�N#���r�a�EK�[���w�WS�#9����H��b_�?��a����r�=���J��xg�:^Z��Ϳ�b�Nuw�6<֢@銇�a@��)�S,����T�x� �^�P�k��ɒe� �4��>�{��+ ?8x�7���ǘ�B"��˨�z��a`-R��,B�����5'�;�=ͽٌ�1�^J(���:{+��S�{-#|��83)��?���S��I��a
�e���f���ׂ��q�˞�ؤ��m���AnS��^C�4E���x<�<���&����5�{"��������f5�lt���*�ny#^E`��!]��'��S���zaJ5�O	�e7K��U�(��tuxd�a��=�Q{fRu��Sl��Q퀫���'[3�vi���坥�*��M�8F}E,x{�P�=X�����.��a$Ԧ�������Zz���p���K�=�l5�����z]�s��9	˚_�|2�t����ůL�³5nƤEc�O޺��"�p�D*���/v�(ΓCB��fe�)CM�.���㗘.���[�ˢ�B�w�����&�΍a%���ɍv{L�ac�ss��^đ����3N��z�+8](�M�WN��eyA�'�֬�]
9B&�������xh����זz&���e���8��3Ei�娦K?==@F��f7��\������)�%)暻����}�jv����Q���.8C%��y{�
�	k缯=CÒo%�od������sQc�[��E2��E�P��u`Ġ��Y�t�������`�d<��
�u�U�����bi�9MQl2嬿S���#�t�ɭ6$f�,���H�0[�DCrH���5�aS3��M���6r��I��'�r���H�³׿M:��!����}��j��=����xWSP�����ĳ��G�b��i�R�.(L[�bؗT���6�h�.�z��I���wuú�ؖ�N���f����GO�FΪ�t�{ʝ[S�j�:���rm�d+�"7��^*�es;%��eW|��| ��Kh/�QÌl�8p��`�;Py���#���Փ���{�����P�Юc�,�X��ZE+�����;�Bz���r��^��uW���+ӟh��5�u����Ls��,�⩩�#4�O�q��
�b�TC�y�`X��|32'�^B'+�=�.1k%����cQ�z�I�WO"TrYޏ:�*���د0L��u�z��OZX�oz����jA�����O1U�'r������.&���ɧ�s�W�7�=�]m
�F���f�u-@�gI�Jj�c ә�����S�,r�0�A�6n��R���6�b�*��@����������w�)ӷ{9E�|�I�L�qXعu�x'G��7@V�t.�l���|-u ՞��Ұ�t;�O+���.����)P������
�D��q9t�3Z\Ls�]����1+�*;�wf�n)�����-�O㣔�ƅ�� �+���V��ko���{'oCH�N��$��h��A�M_j���p��C�e���sa�U��Ui=�qS�Y�S���Zc�C4�.:H�s���v���{�l���}d܅�:ZP�4�B]R	�XX�v�}�7tUue�������0D��+U�ʨ{&-2U�g:=�}��z�2�pެ!	��r:j����%�V�����p7�dN��͑����6���q�8+o�"2V�)�pYƜ��V�<�^ձ\x`ɲ�YUǦR��r�����Y#\y����A�/;-��t!P5m��Y�lϏ#��l2mR��m�Y�g&	P>�yl�7���ӳr��b�*
����i��X �O���!����6�$��ݻP���aY� 7�+(f�ަ��N;8N�t�3��ڝ1"4�0���~�|k+(tϫ��.R�Wi^~�u�C+���TwF^a�Q�#1��*`��n�x[��I+���QY���@`���i#��+4H�p�U�\�Ja�9�dڜ��~����{���Q=���-c��#�D],9��wO�h*'Yl���k��y�3n�
��0m����Y��C�k���18��f^V��:ak���}��M�a��H{dm�G�c��iAo[c1�l�iު�Cq�uw����׶�k�F����/���:�x��W�1*G��w/Z����8>A�r�jZ�˭�E���T
J�~�%��Sg<f�\&ީy�L��T��xÅg-���S*w,'7k{�&��K���i��q꼑�jDF�o@�d��2��[�2�܈Z���RݏYsu�埓�&{@���1#}��[N�i�7�����q�U��Oon%N�Tб�U�B��Y/�

�����@�mV��#�nj<Ǔ1�kI�'E��rӡJ�	����n��t�^i�΀���J�����G�����PX&�%˭Z���p�b�h�Ŀ�L�LgҞ�F����B𶺱(�2p��N��Ι�3r�k�ddjk�&줷̛w�R�n؛tl�o1�O���S}+����8����@�;E#�b�sL�Y��V�sT���wrC��ch�)�1 �{���b�ȳy�P��.�g:>�ۈ�2i'Fp���t�<�0�H�1����z<U{���TS��z��U5ED�h�Dն��+mP�45A��EATLU2ERn�p��Z�f��*�9:$�QAEՉ��9�4�Q5m������AAD_ �T�ALEUTESD�Q4QLV�=Tr���&����mM1X�IM{�E�q���f���)� �mT�( ���J�b!�+�����UUET�U�DTUU�1EIEU��(��j(:�TSEEU$�l�*`��*�b��A��QU5S��bh��餢���)��nF ����*<�"�"���GSÑ��tu���Ǐ:=y����twi�)&y4u6��4���,8m�2��p��wIG_Ӥy�ܘ������9v�73AV�7�~��`7>Ƨ��%��T�����8!��W��.�Xh�2��J��9�Sm˱�_0�湕��Xު�l΋ɀ�#�2po��V���E`�~����b�I;3�,&2nƓt�[+Z�m�t�{��{'�wOK9�&�߾��'�&��	�����B���5\؉����۪G� �d���iPq���̩���S��'ˋ�8�|�O�s��c+��L��wZ���Pޟva3b,����f�/�Y2��T�oYA[�n�72���.��/vT��,����j멖3�h���ԪZ�@�QEG7-��(-8�˶׌m�y�5��q�(enMU�Wr�H���M�G�~5au���xT�fs��t���>f�&�Zu87.�o6�Ѷ9>
2��}������	0�/���Y�y(�͘�kc�^�](���k�\	��ꪝA�S^�ۖ�M\���3lPX;n�{f�$g*��
�eS\��T�Om7E;U���u��h`���_*�t"m�L�c�_�3�~,�����gqF�I/s����v UR�Q�&싴�׎��çs�������pY����YT-�-�p�˴,��P/"X���^�?_]H����)[8nL�e�n�����QǊ�ꔆ��+{8��P�(v��۟�Q����Z\kE.�ܬ��P�j6c3�_Oq�c2���5o޾V!��f�\�Zb���b#�8Z�2ө82��f��J��R�X�3�9��dq�^��5�|/�ӛ�Rս��������0��.���ӧ�x��t^��ɡz�#Rt��
I��,�U[�X���zN)d�E*,���,c���EZj�eA6?+^�<g����`*��B�2AL��7��Tܺm��P�1j�ɵ�j-֞`MWc���'��z$�޼E���!��u����*���u�"���S9.o�D|���	�&���[�t1I�(�����Ƕ6��Ə�_���󤬿|�����#�7Xۡ�Ur�o���,�ԥř2�����^�ʶ�	��zc�t���h���3>��u�)�Y�=yo�����s4U�=�Qk`"��E'���XE�j���lG8W�RO*aI�]yu�:�q+�^/��ML�[}���Y�u����]bx�#�ؑ��A��gl.����έ�ے@�R�!_��G�n�}8�H�~�[;�z�˔Ҟ�2q�;���o���;�l��I���J˵r��&Et�u⥼����#3��/�w�lh��h��9zyyM��q�M�V��r`�h�e��t_�/��q:�/C��C�c����ً�B�Ek�y���A̛m;�!ۤ�He������V3ZR\w˘N�V����=�c�N�_���p�w��������D}^9�yǮ~�2*��0�i�h|Y��Vȹ���}��9s��n�b�y�+����z��X�����x���1X��;	q�mwQbT�=�����v�A\�q8�(��8���UU�S�hO�����Zo)x
�W>��Ok;p��D���	��c����koj|��c��L��J�6<h�:3i^���E�����0�����+�K�0��b��ԇLMeS�1��>��8�:/���Pb�L<�:�(�i�V���D�bt��V�Ƹd�LKQf���� ;=�c(��3�{�Hp��[�C�$�>Vșq7.��F�
�[Ɯ~e}~��j�w������2{�z��n-�w�O1�2箺���}�P,"��:�ؗH��Ӑ�$ͻ�O��i���u%ʲ5��8�
����*�
��3�_Z�N[��1סj�e{�����L:�e�z�젰e�d��j��*����P��VNOlEO1�Κ-���zY�p��J�\]�Gݶ��V~�����5��PyJ"�*����)絀~�۽�[�f��A�*v��7J������T���枡ڵq�����9�Ga�ה�N`��j�2xr��g#��R�Vgs���=;0v&�5d峑X����:�g:�����U���6�X�茘]g�߾��p^��6a�C���(Ak�{}Z~6OW����}���e�B]�9��Y#k�Q�T����E�2�����������Gm�(�9�8!�v�ܥ��e'XE2��O��F۴�7"���U�p�������s���<,"~�<r��Z=�P#�S&�1N_&����+/��}�����M�
��(Q���o����&50��<���N��	1�v]v
��L.��5�""rit�C�mRai,�x�3�h�4���Ha,���⼾>ܪ�MQ�i�5���Z�c���^�Yb�jT���[�	��w>5�\W�������sf�O�ʚ���}���T9fC�o�_UE2��-�����u&r/�?3ԅUM�CLcG=`�IƞR8ˁ݆;��s��<�S Pb/� h���d�X�<���c��g[�3��jKuL��&��1�X�م�,�@Pڀ�����{�:�6g�D~ZD�����KU�6��Q#TX�qR�T7��3//�u�z�~���h�V�:K��^�8\P��)�k����YQ>�ص��=�Xa�=�^c%��킗$���*q�]I<�[����@�r��Y���0w�3?��s�`����дO*}�O+�j�l���iC��D�`����g\�1�R	74��/�Cv��_nr��C�F�LZt���%��L0�`�_�����U�^�YW�������D�Sl"?zQ_*��7Ï�F��0�{l����X�V�4nO�^�1]���Z��r�\�A��'+˫!��F��OL;���������|�7����9xfm=�n��j�J��_�*�汅	M�A[�wu�M�R���P0�.e�1h���r�g�M
[�qm0�H{����w*�[�E��R����[�m��Ve�>��7<>q��̱�{�����FL!�&����K����:O��oǳ{�GOS'���.ri���tD�jW���,vE�2D�	�[�ai���&�E�J܄(d�w��s�)�W��l��pF�X/eO�;ҎW�v/�zYȼEe�1��F��|:���BwU��6ug'�s��u�Ə8Y
�|���^���I��~d�Q��H�S��[��#��[��z�5i�G��15� bYO����vˣn�ޚ���%���Ja	� ȶ�iq�Ss��"���%Z��#�#�*��g�e�}�����J��8�PS�i��~0g��:@{�W���%ao9{5�7!��kDSr��ܫ���,��Y�f�}��=�0@4R�`P�jJ����Y�n��]5����8r͂�;���t�e��7��mn4S�+02���hR��k�
�L�GaY�б{����݄�s3p�5c��^��f�F	�A���x<��<���^�珃�64]m�8&w{���?o������>^��/�wO-�E��Nv��!C��2Z�k �v����*�w�s!c1��"�.��oj�t�*�_qV߽��&�:-����2׏gR�Gh�����1wAL���lt�h�p\)�O�sPC����4�L��c9�#"�O@�Pha>؇9�<'`??�0K�����2ϲ}������B�fK-m�m'eۨXr��ͳ���ߩ׼�ߋ��g��jh��u�o�[��
��ŀ�,]�-��Br=	��9�1�8�ʩl�2�<���C��i	m4!q��nΥ��v/5^ek�g ĵ?,b�v��Д�~��J�:��~��Y<�RY��%sM�m�ɪA�u5=MS�]�C*vKH�rC�$���VJ��L��AO>���oL*ֿa�4�Ѭ�4����[�R��ʦ�v���׈�p��+�`�>�XJ�����G�`�2o���!Φfv86�B4��%�:rM���"�hRU�a)��|�vU��$û�O�M��r�q0F�D�3���g󅞘����SʞPf�;�y6;l�k��(�@d˗��އg��h�o�fWyb<��^{������v.;�m���}B��� ͗����kt�q�)ח�uuޕ˚�a�TטX�1�+��4a���s��5i����~�~ӛ�d����u���$�����%�� ����l5���| �{*��h��ȅNk���'cK�E��.��噆v]�QksE'��UCxX��_�ȶ*d0�Sƻ�M�R�#|�YHx���L��O�l���;r��O�bѩ�ڳ�Hk5$и������w��~�I2��'�ǰD��K�~;R'�ӈn�2e���.SJx#�;a7Y9�n��ա���oڻ�7�P`�Lkm٭��6*?��4�q��&���о�w�c�\��=�;o4�M"�>/�W�����q��6W�8#���G_����C�ͩ������K�E�s��8�F����-q����T��H�wEn#EE�d )�K�Rr�~�#l�֎v�YH}/�$cz}��<�sP^���疕��2��y(?��Q-�%#�ގ�O^�} _z���|�"��G�\�D��nM���y�A��F��&]�i	\�����=���������B��j�oRbj��ϠpO��?8��H{�T���m��w�G���Em?}N9�.�H�7��0��<s��w��b�\��4�o�"�*�G:�:t�gN,x
��sSfZ�|��{/jj�%<�ZG����,�Z���Sb��	������7�FஷhA��X`��9�."�1������{m�F6����ѝ6�+`�g�kG�_Uscw4��oAK7ڮ��F��:����ѯA�Ⱥ�S�k�l�Œ�Wt�|��)�ёV���Ży������y!�q�}��Y�����:���o��|Ħ���Xo5:r#��
a��q��F����T�{�2��QE�+�9��k
j5\3����µ-:�'������/q��-�s�3�?0����x��ld}+����&\�al�~�[B���[�-vK���vԱ��=m�n�kTm�pm�S{j�1��!��ܳG�ڭb��d�x�_	O�[b��e�]l5V��i��v�����2���
3 d?}*���Րx��	��*���N��S.~�ϑ�9�:)�v��ޢw�z!�|�6�`��ؗ4X��/asQs���}gB������Ƚ*"]᩷ ���\��R�����6Jw>Б�����E��5w��Q�)��4�7�WX��s�F�ʟy�o:寪/*H7j����`�CS>� _]��Ha#姮7���������A��b��y]?*�( �#X1˩R�/�e��v%v����0�Si�mDFۖA��LCr���6.�\&��)��#�m�S�md�#�9�BȣM+����y�3�.�.: R�t	m�%�͕��V�m:��b�6��!�&>��
HM+�UnK��u����Ǯ�88wT��N�Z�˹��L�l&���w��*��;��}���w��V�6���co�����1i͊�e��[��걸��ױpQ��4>�`_~���z::�����
<UQ��7C�®���ɍO*�'kX���ƹ�D�ܞ{g���e\1[K}��-)����dӬp��-�Gqx�GIBWs�փ����xݪ&A�D�B��-��$��u�Az�K��Z�M��z�aqBj<1�{�mze&��L�k��znDckb0��`�t���9	%X�ל+�F�}��������!�3�4͑p����Rzlku{�����t�6����]Y|��׃�P�ha�9]<ʆq���^��/�=�;�/����o^㚦��۬.UM�xP�вl�%�+�kH��ܧ�O�7��3mVi�}+�
YW�5�+
�
K�Y5N\׋W�J�k⥓�(�Yjm���v7��x;��ضn_�@Ir�+�����.�<C�B��o%2j-$��k��{ze2�硴��k�9��*ef�w��[����7u�
z��������i�v���L��l����Ml�m�y�X/�T��6T���C��DF�"�5�Ǩ��|3a����XڀN��;J�*�t-v��
B���[_}����[�f����nb��T��z@�c�/WA	ٵ�(#�[r岖����޾1ͭ"�7X%8�+rX�W�7��k�c[�_���0�-WI�Ц�'��ض�K9��,�e{掑�?N�߷��[D�*�Zf*��
e����2K�iWb�[��9����~k�9��z�<x؉g�cc}uS�`�O��U9d%�9���e0���LP�%W'N䝋̗G_5)�i�5�<�g�t�ʷ���N�w�u��9`���.��p�ik�r�8�Q@��屃Р��6]�s�.�ޫ��J��;�~�1��������D�l���6w���r�O��RY����������3O	�^f�������A�����z5}�#�<�����9�b�F󠞚�����׹O�3׭t����ơ��`��g�������ny�|�˥b�l/څy�e����l]����$jb�X"��0��F���,�v"~��Π�8>^,��ĞԶ'W�ߒ3S7?[!.0�3a�~ݏ	�78��h`Z����BSiù�ts��_�l�Vn��;��=��/��3�y�j1��z9�ד0ټe�t%$6׹K0��[�w���H�� 6�</e/Q�%�$�e�L�v�qQ�%6���V��0;Z����͢zK�rޮ�����]��To'�Ɩ�x�*(���)�ݵ)/pIQe�nig��}8��y��	�+9�[F��:�'k�z�m.�s��_\�����]���T�P��f�������{r�B11}!�cC��\�����Tݺ����Jt󐆟=�9VN_8�K��es�q�{�O]���F5� ӳ �3Wo�z�%�^W�'R�[��`K�F��Ř�PK�ht͖����><�6��Z��S�Y��+V�Hrٲ{��tyҤ�o�8c�Ҋ�}iI�:�b���O`���Ύ�rӔv�����R���R��xS����^��ٵ�̼ө��Ӱ&.��U���%N���&-����چ��!욜��M쫣�LK5 ������iu���ŶݑF���A�V�v�3\W��=���|���g���S���F.�ͽ�ȝ��i�۳ r�ۻ�n�1L�L��|Sqa��t��7�%���rgC�@Ꙕ���	�j�B��n�����O_,�gq�6�;���{I4����w
v�oo:�z��FT�)%��BA$��W�[*+��]wH��j7�7�`1�����؊u���-��F*�;��K�E�7�X"b��[s;���I�4��K�r�M��[v �cyNˑs��Mn;x�*�Y9m�Hh������ܵV	G%�W��"
�L0Q��b���[V8Jm�7١�ZȌ���|w�!n�Cݕ�Ҽ�pS:2�ʚG�P��w�u�(�����;uwEZ�c;�i��#}ܹ�ٸ��J���3N�U�idb�[,�l�Jc��_;�m���	ĝfP�W�,���㎱=��nk8_[{XF���A}���ދ�ʛepfS{2
YR��[ۭ���n�������j����}��.�l�mM�H�xV��8�"��p�ą΅���<�j{�����w�U�oH��-�o!��Rt�n��sGu�2����t�^qɽ��/���K{�Ͱ��T��2ol�+lYZc<�/sV�	g��Q�L�t�՝�3H]t�c{r��m�k<�����|�%�dsq��B���YW��_&5�{ �5/. u�Sª9�����Q��U}�]����-������x*K/��}K��W�$!r��9���:r�r�U�L�%�i[Yq�&���	���`��o��:�;����8Ğ�/DF_"1}�<2�-�7��d{XqN+j�\.�ܡ�O��ľj��Y|�cܭ��L���F�u3�+�QH�vϭ��Cx��4�h�����(�}0�Lw
�	�]��XF�l�@�=�35V8��X�Z����S.<w0D�E���M�bM;�9M7�okn�\]֔�_4��?����Ѥ�pY�2�ܣwV�ނpo&�q��76v%#u7dqyPo���@cN"���#�1
ѷXf�*"*#�j���9�QD؊����!�� ��j(��i��lbb�I�9��'cE�D���DY�QAD)� �b��"a��	آ��*i������1GX���nmR�D�US%U40DW0j`��i�&*���4E[1Q�M5EUSR�h�)��[%DQA0`���(��&
(�($�
�)Jt&*����y(��������N(�

������"�j�"]�	����b������&Z&B���?���H�
#@���x��c1�7d�t'e\��V�{8�k�|�>-���70:ܡ,�K[s{��В�x34������.Xuf㏙�X�5�B:�K|4�<G�ڽ�Xè.�W��P��|T�b�49�<oI�2���d<�S#ѧ��T��tf�R�d�G0���ʥ�L{#����ɝ^�?p�N��~�?m��(rs����~tŐIM2n7١,��b5VC�PaK�]�X܌����Jf�W��P�g�*M�}�!����6����+G�:���;��D楦i��o�+i[�f�I},�+$�oI�W�ph�ήac �.�"�
�/��������s���h��P�����7Fc��C��Oh�v�/ �j�nt�;__e���������,�Ɖ:*����g�R�5�Y&���Bty��!�\W􌼯s��u\���B.�'�n�ժ�uL���W
���j찯�C;�dkhl>�:D���~��=�E5xv2�ñ<r<6f���w�W��Wk�7���*1���Z����*�r��ˆ�A��)L�%1����t���4'��>��q��C<͕�pGW,d����<����N�^>������ȲL�OT�C��꽇v/�����1L'�\��tM��ɢ=ob��Jpͭ"�'u�}��7d����J���5�[A|
m��u�]k��������./t#K�;9G�1ғ8���l�VA9��	%��Z�<k+��_�ﾒ/'=��������Z��;S���s�O�cYm��u�*,4'����6��N%/���J��tN���"��"j��_b�� �������?��cn�c�^��.(��[���p���j��Uk�Z�v�,�e�X��/}C!8}{k��z������g��V:����)������v/x��(�X�}2=�W:3��ڣ���q)H{&�����Q/fK|���y]��4���:�����5 ���7�\G��[c��t�����"����t��7�����ܭ7�9��b#Z�C�re���Y��y`~אe}�(�Df���;y#�Ӵ�BnkXF-,w5!9��!�7X�ڜ�՘A�=��Fǒ��9V��y촍�D{���Q�i�M���J��ދس]����%�ik��ϫK�r�r�)>߱m�⯹�`�`��Y�d14N?v[rv�A�[ح�=,�3�̂�6�X��ɨm�OxJOң��[b���Bp�4��sn/M��:�%�>��i|��J_�.C.��l��A�Er�]�BN�
��m�-C�����-�l���'MϚ�R�&���:�B��Մ���t���n��տW8���٥���Y%�!�ͫ�n|)��S�+�/�3����١�uΐs���܏�սT.�f�e=;2�%Q��^���V�XV.7���x�e]0��7��ۑBC���0pv7[Os7ͭ��c�Ȫ��v:���D��W=z"1�C�\�.E�6�?���Х���p�F�6������ �wT�<�b�29�<�IJ�!G4;�"�7�~x�cR������U����U����Ji��N�OK�Z�a~(�b�G0�P�ϭ^�Cø�h�������A�y����Qa�>ج�&59�6��s�
�*�8�7�S�~��N�Cy�0n+22��x٢��g�y��2P��9�;QL�:K{�����/ظ(��%�VY���;�K7Q��.�܈9���׾�O�_�@�־��dƧ�\���3\W-o�JV�ouS���FA�.�W3өU8ձBY���w�4u5��rl�*����eY���u��n�������l��v�7Y��#5I�)U���èw��l޶DZ�FyS��Md��9����c!k��1�²U1�5��R��^��)�>;��#��D��ʢ��^�,�Fg[tZm_z����<gV��sq�����'7ME����c}�T��1�v����$NP�!ãR���h/�W�����_o�I� [�A������L��)�\���$ngp�E��#Ǥ�
��c ����z#e�#�U� �n@�l��X���
����p��|q�7YB�P��Q�-�0�E���wf^90�fC襴�dWX���ϼ=}��,�S�Ω�FT�W��i�[UlNytůP�ز6iYB��j֙T͈���1at��_t��G������y�|�����i��W�S�|>�4�n��k�j�l��8��j��Tޤ˿g�ʈ}�G9P7�h9��騬�=p�)�Xef�`T4�j��Vڭ��q�e�sǕc��	=l@�y�+���n�������2�Z�xUH�~�=�K��F�"��1)� ����U[jΓ����Sэ)f�}�h�C^X^��Y�t�2V4#79�<�Ƒq~sJ�|�b�����F,�2k(�1�'^��`�Wo��E/����߬������ȖR;Cz@�&(E��ߔA.�(��07c5��]i����<�v�O�A�9�BCl1p����[z�e�H�+M��]���d�?7Z��K�(�q�w���R^i��P�-.ɼ(s�m2����(ϼ��S�ƄP�f�Y��|���G��#FY�w�]���B�_�^ߛ�^�ȏW�2@��{�!�}��Y�C|�����1L�M��S{Gzt[��c�f���Q�J���Bp��
�-iu�}۟�K��K��U���X�/=���"�B�*����B��i�v��O�O!�s��<\�w�e(າ��*q
��F;��f�m��(�ͺ\��� �w����1��q��7�+5��jm�V�?�ٲ��,jnn!�lPXL?i��ԫ��,�gX�����\��^߄�sb����˟���K����o�����i$gg��_L�X�B΍~y�<��n�0¢ٚ���7�v�����i%)���̺13���9�r�����t�,��<5�L$��5�,d��=y�wM~L�D�)A�(f�D�)1G`?>�ܭ��W�9���d:cy#��)��8���^�M��\��G�y�t�p:B�#�L%�c��j�wd�Q)�n*m�3b�F�>c�P*�4�e��S�f��e�ZV)PDvV���[��S�g?"��y^[Զ��������r+���2�|l�75��V�z�ZOS�Խ�ǻ���ɈK�C��x���j�No�mV�sҌw�ћʩ�զG�F󣪢�c4wwԞ���g��Dz���fy��D��..�R�O`���^�ʶ�M�K��H�GU�'��;�k�����$\��_j��9�sz����*-~�B*J|�*�.��j����`��2���$m%6�[�?���g�̱0fz�le%����"n�!�����z����2�H�qSуyw[8��u��Y��lU����Җ&r�`��5��k\����T�&��M���{)| (��(�P[�t��J0��mXZ���[�Ӈ
|x������oY5M=�~��M���_ }�*��)3��s9Y��w5�s�w�a��Y��խ�5O�ۗ)��w�t=юI0V�� ��=_�}ʄS�5�
L�t�[Eg��%7�e��;X��)�k�׎ܦ�����s������jl-x�J�sf��>�Rӷ^c,G^���q/��F:�YB�عZaٱ����?v)��}�{c�U([wLK	�9�·���%���)yĽƥo#�`��6"�3���	݈�}�*���Qb5�ދ�����SVM�kB��S����<h@����?��Π��X�=�EM]lRL��W�s�Y�N���������"�)�2�[N	��˪��͌f���C�k�Pc���Y�ܜ�7Q�m�ٺ��N��A׹d�P~�+��Q��1��O� q������MK55-�ZS�ɮ����k8EBf׮"-�R��y�u@ty�D����ɂ�L��31
&�Ϸ)���/fO�H��<v����UK�91���}�c�5��6f�᧲�!��3�&�l��S�e��i3��0�hj�Lݛ킡ܰ�^h7�õ�	�}P[��PlB0�`T�
�WWղ�Z�wE�C� ���Ы�]�1�72M7�M�n���澾�N�e]ñ>�J�e�n1��v�V�����퀩��v�:0cw�������'=���?
�o"���P�ek��2��Z�/�YT�~�=��e�z����ѷ���.�jΘ.�$��p�\�:O)̪��m�<T>�X��M���-s�)>�Ŕ/J�� �i#�;ۋ��3'��	��x?[��L� �'��T�s~�%���/�T�q.����������c"e�#��`������̂?}&|ݹ�c�����&O;���G�����{��=AE2��*}��v6ę���
�GW�ս�����Qs��6�E�wRm�5��l[-/���|�t�L+�Jb�7\�5�ѫ���#���X�OF�5.G�����X���*`o]��>�;u{Ƭt9Ek�Œ*�q@��Q�ȳ�O2���0%*��R�*�tqը��օ�*b-���:*=������C���Bz��1(����%i�/<���x���/
fz��H(�����/,��=�[��YC���9�"�;#�߱�;�e�ǻ�Rzŉ���(o��S������-7����D鬒 �^lO>���b>�ac�CT+9=T��X���{�\�e��<;J-v���O���Qu��=�*tH���Dx"g�M�Xz�;�i��j+��߳4��*�9�`�o�F�Bݹ��ep��T�+�2�%��ӭF2���̲Ϊ\q�F���	ʰ���h���D��^��{ϭo'2�����ګ���	�(>���H��k?y��e�2~Zw�m�֝dYݭO�fK��U�'#�2��K�2��G(�ɪ����l:�F3�nj#�0��Q�âق�y�*v(,���XVSl�ɂ���T��&co�sro�jm�#Ξ ���u�ɚm�ӱ�=P�J���=�����j̀����_YHݭ�ik��c%B���9^]Y�`^� ��X�c͒���e�"}�K4��b�.��t��:{��汅	M �	e
ǚ�K�
���S�k��(�߫��Q�d��L|����{� �ܚ�m�S�=�C�\�Uk�����C�9�Cy��s�*q���s,]�\3%��P��C���%:j+�l����1�s�d�B��q����2�v��s�QM��+RQy*�\3ci�v��	�<n\�.+9'3�ڨ7!��*��x٧���S	�J�l7o�	�ma���Y�+2��8g�g��K��i��iز���m�c�On����"G����Hh��8ŷ�~��S����_�8��A��uy�t�]��5ZM4��ć'�R�[��ʢ4�];�.I$�>9
R��������<��ܐ
C7��ُ[\E�^ �%����x�V��d]Ew�r��s�6�F�86�7��Ο��T|��{L�S�~g�\�"���ۑ,�vR�oP�^DH%V�.���Gk�V˻�	��C��>Y�m>��W$����9��sy�C���S-�7)YllR�o
��v>��KC}���αڋ3�>�^���fx\Gh{`Ev�A����L�_C���g[2��~��<*���o�j��r�Rg�ӻ3��!��k�71�̖�f��ݤ8�V�f������V�r�O�;����:�#Y��oz3�z�]S��w��k����5¾�`�m�6���%,c8�5zw�<H�<�1���V�Y.��h`�3_*n�dA�����_v�io���v���SL���)�K����'Fu���o��~�0%����.��W���g�\
�����?�_b�a���\��r�NƲ�>-�'Z�iT�4�OY���hE�5�M�#�^�0�CL��\9�{��B�!]���G��]ɬa˔O���pxQ-g.wuvk�����3k��sM��i�H[���N�^����4���L��H)�5���{t�Kif�v)��5{��Fۗn�r���zG6�0�#{c|�=�\�;ne��&�-ۤ�\���v�(cnwWY1^ڳH�>ov�V+و RߖS�v�׮s�˖#�X��)��=�N�9I�7�F�m�ju��յڢ9�"cl�4dYBh��e��F�m;��{�?�ǢV�� ɪ�K�Em�rȶ������-�#�X܌ږd�L�f5Z
K�R�4��d��o��s昢�l	m��V'��Q���_W�bk=�����`U[�G���1���߾�t�g�;C����8&%R���q9]m�8+�a���b���������Z��M�v^��<c	�O�2}��f��wG�K;_�),>5����݌H}��7�]w�n����7���t
�nM�0#�WcDc�@K�qr�������E֮�E}۳��	�y��O�ޟtR�{^�"c��{�����$�+H����O�P�'�b��s��;C8�.mo[�	d2��S�T��
2Yk��B)�(tc�v��|D��}�߰����m�/�S�V��ꞓ�J4.��0���	��?ߧ���쾱���"��w�q���|"�|�y]�����ս��(�Z�8�[�I�;x� ���ucx����訰Пn�*��\�P0�m� ܦ�����'GF��c��u��mgBf�r�[�w�2Xf�@ p
 �>h�g��,�y�	���YW�KP̵�XÖlk�j��@�L�î.�C{
��He�ݕ8����0c��κ��SR���'B�C�J���{����V�sx4�J�W��ڏ��N�1$^Lك���?`� �;=<�,x�6�*�獁�ˢ�s/2k���짍�D�����G��A����FJHt78Q�x����jް����Z\�1%��zE��1�A\�h��ݗ��e�7��4�q�Iu��Ƙ�ͳ��
`�s���1_���Y��Ư_s�bgP<�2��5=舢Uq5`��G�d��e�j�����gs�x�rmA{r��UW�1_[�[���!�RA&���'G�-u^���j�dI������+���Z�ao њ�_��:I����v\#���3y�;��;�)��~7f7sB������i�3%vw��`b��,�3iPK��;-+k%�鬮q�i0J{���(�,�+ڈ�k@xgJ��ѵJ=e�����yʧ*k���#��zt��=�m����a�1����%��>���@�-�x����e���u�S/�]jL��L��!��9�J�r�4���N���X{ �nw)IL��9��h�yt*��Ȏ�]8��h��n�h,�;�@��!93QQأ�_ PF��Ʊq�t29�����_���Mb��\ZFp��rLJ�o`���Fh�Ҹ��6K���gp���wS�Y8�I���5ތ+8°WJ*�}���ܱ�Ԫ0X�A!���j�!�
V �(߈��w�K�y�ļ���-�u�B�j�1�D����嫵�l�\�P�M��[�bu�Ä��D��P �g�չ����F�Uw��wm�`\=�b���+��\� o7C�6:D�S����)�_^�&�L4f8��tɼ�]�e(�E]��vX�b�v��v]���K[Z �-o")5��D�C��=j��k�٥�!vf\}�)�ib��xkV��O,�| .����f�B{Z&%�9�v�<ܸ�+�]NK[�{��ɵōN��ְX��;��:��Lr\�W�J�+#���ً_	@���6s@���Ml]��=���A^���fū�ӡ���a���2�s.P/���kzX��R.k��:yq�2�Լ���^��;�,ܬ�}|��I�ųrGf`r4n�Dn��yQ������b����p*Sx̖������d�����{��p]�g�(c@�8�a�� ������<��Bj��-�㣺,��+.�+���O*K&ރfn�v�d[�tp2��C��`�Jmݩʮ�=O�G9[����:�Zʐ:��c�nc�[x^�/MV(���ò�[��z�K��11�T/���7��E��*f`v��k\�᚞�fh���n*��{NL�hlշ-�bޗso_w�Q�J�m:���V�խ��N�+�ǅͪ��r3֯���[*5��M!t8��`@FCɯ�O�a�X!
�J:�j��/�e�/߈$� �]��M'Q������J�
"���:"�"��(���� �	���)����SAEHSMSBPQ�UBU�QAE�փr�D�URST�E%)HRQJPąP�HS�@�5H�PDPPAQI�CLE�R��'Q�k�!�=��1���()4u/ �y8�
(���)���

i�h��
(�
J
�H�>d:
i((Ӣ�B�-�M%ESJQ����IB�G{2P�܍��(�h*��(
��J��)j%��iRD�-4�S5T�P�� �v{���랽�[.���h�Aӓ7�j��ݻC��э5G���׹g��rb���(�Ю�	�jN�`!����\�{���9Ϣ|σB;a8^��DSa5����1Z3i�X���={Ƶߝ�ay�U�a��7l�߳R�~�D~�4�诗�����G�G�;J���Eo�{ō�2��۪�w
�l���L⑂�d{9U_�a�~א�Lo-�;c���@NIO��ƃ�&�ޡ��L�2v/���{K�n�����]��.�t<�	��Ύ��L����Q��oKM�D���<�v�e�gW�(�W/�o �]cN�����Ϧ�F 9V0���mL?mK\l�:k�sC䇥e�(�B�,`�?�M���7��G�����&I�R}�r+=�-hn��&�Z�t�g놧fY�#w�����Ħq6�n�k�4Y�Bcج[Ct��ѣ�ީ��)��v!��3�	w���m�}콊��L��,��Qx���C2�f/�;OFy���kv���^x���e�\�*}����&o&(s�e� ��_�3�{��l����)w����Yy=�n��a1OaEJ�X9�h+l(xvl͋���RJ5Xs�XʞS��H�Gu:�p�]���sC�0�m\�[�f��`zN����YΤر���V��@fm����F�2��{]#Z�m)�<�E�	�7Q�'���~��o�h�� /q� ��,�K1MS9�pb��v�kr.�7l��|��ʹ��n�u���{��Υ�8֬��<��y�dˎ�9j��F"��s
	�Y���g�ނ�XClO]M#��C��?6!1	��f	s/����6/��0����Q��/�NU��X맴�rWf��	����;�/�@P����y��Ш�S�[��'�Ĥ�E^�c/�M7H��QR��Ҫ�ƻ���A��������-k깦Lc��h6��E*��GL;�+�=��/���b��5�B3��	�$N�t��4F�ҟ^sw��Œ���ʹ!XR֫Uk78����z&3H]1�6C�QYԳC�(���ٮ��̻)a
l]��ؾ�5���I�k���̓/��;�e�J�H�)M�i�3L��;a{&��nh٪�YK����b�SY�1@Jw�w���wFQ���z/}�A������:ʄN��9�q���la�+���7�p�>�F���T"i@*���S-�e�$&�<�[+�S����/��' ��m��@��r�G=;��,�
����h�0c�*�ג���=���|���2ؠ&���򊹲(��h�j�<�FK���i	wun�g��4��wf�j]�*��X��s�B�J�L���\���Y���6#��-��	F���Wa4�\�i��m���7,R��Nǜ.�UuY�o�m�_�G���l�����iz�#4�oc{h�wIT�v��(;
��!z�]�&�j�#U�+���T��wrz�{C�ri0���ZUL������Y��)(����C�4���3I�tt&�3S�Um����4ˢ���C��4��s���R��*��t�sbbۡ��U;
�b;(�y�gլb�]��҄&� �v�C��⃚U���R~k��i)X���a�����#Z{7>3E�Q�%�}�p_Z�=���e=���u�LP��*�=�K�Yx��-�51D7-X�����*G�`cD�W�P�� A�!6�����PZ[FJ��Z�W*��[����;�GaӖ�\�m���h-w@�˼��S�Ŗt�Y3w�R=�6�����ղ����T{�j��RMV� H�v5��Ȉ��כb��%��]Z��s������e׵�Df����")=��g�d�}3�nZ�{�:� l���o�l9��p���΅g�!xC՘�
3�����{������\�L�wFS4���ha��:Z�]J.աc��	��|6W�ͫ܁�o�+r�v��=Z�c�� ��L�u]��%�ث]L]V�9��x���ô���oW8�X1��b��r]+hS�.:R����L�N��쇓yT4���V���d���{X� H�J9��*g<��.�����?�m���1�CW�䖆To���v����4�ApZ����/�YL�[���T���Qς���9�1&r�ɗ��	O��U~�2���l�'�����9]�+wm�U��g��,�n���~�v�����{t_&��T7&��(�r�\�����Z��	Cs��y�^�W4�~մ�'��7�%~X�b�{�-c�yGB򊰞ڥ��om@W��M��΅]�U��G_Y-)ṭ#�M�
�ֻ�U�����X+k�	�����I������L�-�vD�錸N�v}�wZ8�)/�8��n��T�n�z�����<�%f���C���>L����u��*�ϯ�S�\\�f��}E��]B�u��eg�k~�����iS��K׺v}�N#@)�=ټl����^�3��%E��Tfm݂�%����z�|Y�xzA�Ab�bUІ4�vS�c�B^;xP�!�_�P�l��w�	7�*߷>�W�:e���I�y<{��/�	�n`rI��i��z�]�/�yW:${6�7��"j���ޙ�/f�s]r�ZY���1���\ �:�/���#/n���P��wf����gWW�K��
���G3f�\�5�Km�
N���#"Dҡ&PnK��dY2eJ�JR3�l�b���ٳ�&����V�][�8d�׎\���⌜t�}hE;���f�}����L�G2L��Os�4증z^q�<��Ξ4.�T�m��hN�SO�E��5�^�l�����f�;��:�����[���R,U	���1m)ߴ����`'�[r�}S3��d��PJ� n����'��è
�J�,��"��Z���C�ڶ��%�ԳCޏ�*�b�Ԟz�~׻��C�����݊���%���b�V�ȶ1̃Dl_=	���oS���=^�wA|�+J"�*�>��\���z�/��w�D��O�?~���Rbj9����{nO)tGN�oZ�X�T�k1�ͅ�S��鯜��R���	���f�����{�/O��|�Z]Q�]O;̷�y�'��9�R�xGv�8����-�ZݠoyMKt���܋q��tu�Ɩ
�v��.8Q�Wc�VѢٜ�g>�ʤU��%ԾW�X����Y�C����YB��U�)���*>�K
u����$S䏹�=��P��Sd����m�E=�Cc?,�i˶msG��_�]=겫. а3:�3���͉�M	.qOy�B|հU^D:�Ս�!��3f]��	{���9�x`9~wM!;���#�GwoM��%�8��{i�[w�ud��l������K�r�֮#ڊ�A��>��֪�l��S��1���v��_�
�TpĮ��'��ǺjJ��E\�G��(?*ߠ�hE��C1x������k�ο��˺=sV��c]6�zs�+�K�0(ߖؽzN��K�Ψ�!(�H<�T�(��Q�~�6!��r{�)�Pra��pi�t�[ҋߜ̤�E2����Y�rf�c��Wԇ���|Y����%�r�u�T�O:�3���2�0���-�ۃb�'s�	�جe��ϭ��'����|`����ʣ�F<~�r���H������\��Q��g�O0���Z�]���g;v֚;6"��uVZ�eBb��2G�1�Q���B�v�jvoN��j9�9��Mp��f=�T*�	��c�b��� .���be�o��3O�F�נK���,���&���k��OՑ,�;�6,#;K#a�-^�:k�y�~U���+�0��
�:�"0�����[�t�\,j�h������J�\��=�W��5�k���MIj1Ba�U�/�-����緭:���g{���H[�v��w��W�YM`��g�/���Lf���W���wU�4�hk�s�x~��t$r|ꇈUd�ݱ�m���>a뼟�>Fe�r��s�؝�{��Ŕ&B|��k�슣5�h��sb`�ܦqG�Q�+*c���� -�8{ȼG+r�8.�΋��J �{�a���Xf���2;q�˸1ԳjS����5l�� uv2�޼�QYݳ�C�����GI��oӳe�Md���v�/2T�s��\�P�mr,%���c�#����7⾚}�����P~�	�ĠT�Yȱ�����T�ݎ[���A���̹��ϱ�BU��ڔK�8~��i��`���p^��5�������y��>�/�)�*�^۷�*h��MLX�'ٖ���.1��+h����W����(Md׋k��L��M��[�ۥ�U2%K�Q,��V7���e��J�bV�=�\�S��E.�Uv>��3<ta{[/݂v��9Ь��bKb⪙9�m��,e�	F>����uN��� �ۓ�}�Ш����韁�#{�.���"�Or���."�����嶎M��E5�.J1�/x��&���̽c$�P%{�O�����:K��^C�<ieIN|�)?5�Qͧ�9|�&��U����2�r�T��###Ψ3�@�հ[3*�k�Օ�Б^%W'���q��;��9i�$�r���d���K#�h�KGC�Mw�6���l�*-mࠖx�17Z�����z�,��s��qf
�����+������s�G��dh�CԮ�g�NӗՈ�Q��ۯ���т�͗:4��33\��o�Wk31���*��o�RWpBE��(�LE������h<��wouD&_(�T���,ae�ò���$���K4���-��B�	-��.�O$8��E\���h�f:	�i^w�t�3X�`��{7@�[wZ��Xim�rQ͇ا��f�N��fu�FK���<}��X]�M�s�=���c6oy�53[+t�)�c*ٶrQ;fH�n��L{-���H}3����-\�����d'�V3rU�E�f�3�{`����P�c׳a�ұ�;�ȿy�Ӽ����i8��i�\��­�ks�xe��_0Ym�	����f��O��;6��!�o�cl`�h�tS�̤�=N�F| ��Z	d������Wə<��%<>�?qw��t]����xw��d!B���3��2Ӵ.RC*�	g��
�t�\b[�A�б�1���5�۶�"�EI�x�4lWu���:��Mz��,�k�If�J�Z�j�v��τ�Uo:I�W۪�*�Oi�o��{y�P��@T���j��u�� ɸ�ɱ+��N��ֻ�!��=��Y���WR۵��g��Sb�+���]��t�t���x;���'ExG;�~ b�M�E�� �	:��6�f�嵰���F#KLs^]�+\����R���8��R�m�:��ҝCyw<.^�xV՗{9�,Hp@��a�U�8�{��M�޳9�2E�"�*j��6�$M�Jue$ԋ��3}�;(S�W�Z��Y�m�N�Yj)(ū땬�v(U���[�b���?�i���;u��j�w��J]��GRvy���T�řRu�%���c���s�vS���n&P�@r�$��̹�ϐ��B���*��}�t����\��{7{S��}��) z(�a�*7�(�[��dC��#L�+�=ϑ2��Į�Ρ��9�a�iu�<mr-��ʞ܋�m�Ym�ׯ]���B�=��+�v#���l�~��}=U�#��ue�yT�1�U8��U}P��k�z;gv�'��"
�=j�t"�2����L����FF�m+��&�3Dja�&c�C��>jր��þ�Q���h�,�byY�G�\�^StW��|չ��*��km�(��@�\+4l�r��Y��.hّ"`c�ۭ����s<������GCa��̓ǣo�"���Ɍ��s�^l�{x;e��uF��#�h7V�-"�\m�r�S��gϲ�`���6t�M7��:m�jW���W�m��N���}���ڻ3��M\�u�iMάc��]�Wj���Y�ݞ����/���wq�Wh��{��7��|����x���Nu(Do��QY=b'��ć�~���#.n�D�įG�Z�%�{�����~�f9q؆���LN����(BT�YjlL�eCP�[,�;y�����6��2����Q:��I�E�]�Ѝ3��I6����[���X�ץ��k�Ur'�=U5�亽����)������̻��Yw��us5L�l�'b���w�6[�Z�*�~������>º�.`���k=�"^g1�Y;gwvtŮ'��(�lR��̄�M���O0�mz�oY[�M�|��;�^	�y.+g *���"��2 r�:��������.=ײ+hd�Ⱥ�^�*�5i&X�(t,�WJ�r5���v����ct��tgI꘽�,�K�B�u�h|�2�)�.���"mW�s�9�7:���+��+w��v�dK;�k��9�����ڹ�
��g!ww��)�qQí��=oNg��X ;R�f�ޑ���'�8�xqI��r|�~@�4��p��	r�r��۱:����c�d����WJӆ�V�F��:��(���j.vgv8�ѳ8�IJ�_T���;`����9�c��`�jװ���{�;��Iwp��e�]-�Đ���gj]F$uuM�:�JUt ����s���d��UIV�g����fVl�m�������o��C,�j� Lzzk ���ø�^��r��l�fԭF�m��[�ݸ���T�>*g��iZkK�oA��^�}{e��Ù^Ҡ0K�W,zk�A���8LN�ox��;�#Q�r��=�u�i�<���Ѫ�t�kqX&$���`oZhNf�:5���1�e��)ǻ�0&���\9=P倻�G�r���x�5R_TD�P�Л�W��sϠ����G��h�N�'k's�Ɉ��D�C	a����_"�tu'Yc9n
�Fh��otUql!��ռ�SJ��k��绱��}0�r�,�.׀���W7{'��w�mH�n�-��� ��1�]�(�8��[�C�e`�Q��B��f���ڸ����p�k�S�އ:PfG}Y�k��i���[���ضV�5��)Z��cXx����!֬Q��w@�o�� 
���[��K�������;h��o+�� _|�.;;*]�\�e㒶蝜�-��+�J�r�eh�}#�|(�;:u!�i�J
���dYY>4^A`WX�%���/+Y�smу	1��
�e��d�݉���l���;�xsPk���lBb��WDq�v��fa��au����h�~⎮��Ǟ�`�ۦ���0*��P�J#!`iS;b��j|��;�.�f51��� �ej�1�tR;�)�ޔ�[��|�Jk�����ʡʔ��0G�-y��qM��jܙ9P�e���-��{i.aM�m��-W=��͕��.B�K{��vh�*Ty]E��H\6tp���:��N�����ѳ�a2�v�'�dʹ3��0�O`�k�����=��W1��Hu�����@s����/adn�W7xvk�*�eN�hm*̆1C�5{�ۺڢ$�Ŀư�JcowW-�C�^�2S|m���J}[�)#��gn�a�5�Y§�x)�Z��8��%��´N����^vec2��"�������z�a��6
Ԝ�]�#ȯ*f~Z�ɽ���U��v�aS��u
�zT�%�i�źT��(�ŵ�dП^C۵�����>�M�棧僓ur]���&�tqo>[����z;A���N��$����+�E=�@��qK�����S��d�uJ�x��@	ϋ��l�!���jgf�	mw6�^���#iӴ�)�g<�XF��WfFԮse<�1��LW*�u�WT*�!�ػo��ꨍk�M.ħ��V^�^��7X.0r8Vr;ݜ�7(%Wfr�L�2�1.=�,��27�*�s%���i6���_�.��-	p1��;���e�Ĉ�3//hhft��:U �"-
B!1�ї�TN��˰�k��Y�%�6�$H��'�t�1r��b���*���r*���T@SBД�!E�Puo|��9�T���UTU@PU;��%(R�PU�u" t�Ziz�0C�4�`&������F�*�������Z
4�hI�(���(��
��iM%=��bV�(���)G;�rZJJ�pS�����4:i;��r �!����))�J��4h{�2u�(N�@P=�r�)T-'q� �pj����(R��:�)Ԯ��]�ATP �M%P 4���"|H�S�g@P�{�GO��c>Z�޿�8���=t����Ro:�]a��vT���f+{Qd�d��F�|9�5�����������<=�	}�����24�n�o6	�ih��Dj52��t���i�j4�$0�h-[���KD��K���^��rF��4}ņ�n-�O�m�ܘ0U�5v��l�&i�i쌢#sG�����q�y�y�?o����~�!���,��l����M��@�Sx�gſr��j-��)R+�l:��$\�5.ʳS��E��YSd����㸦5�\3P�L�Ef�n�Ve���M:�D��h9}!�#���0���t����[������R��߯t�	��0H��*"%i�7��S��ϕ�*��f��;�@WՇ����;&*|�'��X����j�����uW�"մ���ެ5Q�%�]>�k��9�Ga>v0,~G���N�o�~�We�A*��zͭ��eV+w�V�d@v�ܷZ���ꎒ�����Qz4Љj#8?�k���FT�����|n�W�+ǠrmU���+���Ʀ^c�M&�k"#��חZwe�큼<\G2J"�]#Z��'t��!`�hdx��8v��ֵF-�ڹ���V[���`��o���vC��n�جc�'ԛ���%����WWR��^��;X�F��s���-6��[�H��{���F:H��k���J���<���K�sʊ��ʬ���j1kmX�7�M̵����r�WQZ���p�ϣ�پQ���\Q�и׋��Y�}.C:�-tz�KH�,ᙅ��w�6y<	޷�a�ǣ����Ng��ws��[�+�A��l%�Y��rF��;�S��f�+����w[�1�������������n*�o6���2�)�y6��0~��̨� O`s�=�Ϭ^'�&.;h�ŝ����ST���$[��s���a��/F*�]�|�5V�}7%�V�wZ�'���m�3��6���C\�S�������V�8��T����
8/��waG,->(�{�YD��%���߭c-gՅ�����8�nOS�Pf^0��>q��oQ­��<h܌�w��ܕ؁�E�y̲�l�x��L��@����9 ����<,��$�Y��2_��v@t{ˠ�+��I*n��cv���y�cO���wE)nN����uI�&WvAl�!�\)�W���w�uΝ�������N-O���Q����j���r�@�GagT��$�S;�Tk.����h�X�t��\��Ѻ^��+	������GO=i$�D�f����x����ϗ[�#L�<dx5�"o��y�h���ʸ��;G-v���@r�&�0R��pō��E_C~�]��oݱ�dJ���7=�7��FE�&�ҡ�(_ UxZ�������c݂m�K��'/V�&P��tե����~���)��z6NX�K�2Mzʭ���P�o�8�LM�:�w� �Ǽ����\�&���֚~Лɋ:W�Z;�.b��R��z2^*���q��\��lă�YN�r��[7��+s��sCk��ܵ4��3��[&��ݿ�*��4�׃u���í� �/X�P1B|E\l][�ʨ�v;}�=�x�]��}�	�-�����p�T�D��i[�:��ߴ~�;��Ω�`���3W+x���B�;�!]�6Dm�����C*�Ah�"5�BF��k��Em���in�׸�X�3��n*����P�c��:�t�u�GnY-hoK�5��݌\�3���(R�Kr��r��2�%�-��"��m��9xi�n ����˒����)
!�r	d2�3"5�+۩W�>�䨘�[�/so�V����a�+Py$=/WR,�mne�fi���*�Ǯ�ZC��}f�E�1E��aђ�����]ua
�y�-르�DTV�3����ja�����fl���V��{�[�v�mc׌��\�29�܁�v�	�`�����ǣo�*1_s�wb^+�]�c4]Y��٢�R��C��n-���nT�L�<l5���:́��3ح;�v��R@D�U3k2/7�t�"2}�P�U�OK(��wLz�3S�U{���icO5q��16��bG�LO����T�.�j��:��L�p{-ۊ�O6���+���g�F�)�8*�`[�u�P9J:�yꯣy���y=W�g&*n���T=���*,
�pk�����S�O��`�Ȇ��ױ�a���?n��F��ڴ���̙9l�^22�M�`��'�Qu�SE�!�v:s8,��fۄ��/
[�-�W5���W�>��1>���&l�6�{t�����ES��ۼMu�5��f��;�]i)Pq���Ǘ��[A�Ծ���E�U�y�xb{(f�a�*7#�UΡK�\Z6�~���<<�=�K6�K��}Wݎ0�� �f�ǢS�G���ga4D�on��C+��w�V��{X�΃p����-X��_����:�I!�H����˿0��2wlq�x�6!�-�m�n̘��g���d"�꾡.�p�u�h�䉔Q�yK���=śϾ����&�yU�vY��O���\oxO��ɳѣ���W=1��3�]��Z��t�L�CP�Dh����zDBF�'�8�qI�Zo�t�ʊx/�[`�ݶ��׷ξ�h�3�[q��>m-N��Q����"�3��*���<�Z^�qm�F.���雑��:�>��g�ņ%d�Eѭ�qriլ��<.�t�ݐ������ĶH�'���m2n�4����V8ڮk��ԧ{j��.���L�E�1z�[���a|-'x{��)��U-jc�SU�I�F�;0�d:�m�B�"&ʬ�/7T�䁖D"E��qqٽS�ǲ�cz[*窥2]M���Y�ɑTCY���i�C���L����d88kY�e��=�agg	�
���.�vAK�[����ʑɡ�D�/{��}�_���;p�7�������8�|
�)LA/e��&̮�\	K�|����� [PH�gX��8�Kgw�l�v�4��=�A|Geq���o��L�����R�f�,wQ�A����}Q\�}�
����sӑ�b��`�S�w�>�U���RC��\�Ս2�g���!��T�﩯��ۍgki�X��t_��9�X����wA�P;V��Y���eb�|�e��U6��F��ѢG��l<��qz��o�v{62x�A;fqx�IU�����I��m�8	�ֻ!�﩮a#Մ8�<���Pn�<��R�
���3,����٫���7�m�y�j1T��p�6�W�����\��:�9Q��	F��nLW-��"�AJ��0���k7��Dpޛ����h�=�v~�e�VR]yS�������
8vή��<��D2�>��"!oul��-�K�Ω*��&�����Vu�-~��uH}�ͼm5n��\�i�2�:���N��	�b���a�YVu�h���ω����ikM#䞧�z���ZC{��(�KE��~��DLȪ��G�[��k#Yy_:�h��l�H��|�\��1�}{�����?0y� �\)ҵ��-��s��5T��"-�#uF�k�� �˧�7WscZ�2�f�%'�Դ�!���հ�R��?��|��uW��m�6,� �M��z^{�mxۍ@Y���f;{�B��׵D������E��<��'�.�{rE樚��e����� �����ޫ|�GD���u����FY�8U`� _c�`�\�����5�m�����HJ�1�V�b���5���&ͺ���5=����T�ٍ�Z�+�V�B%$2G mu;Z4�{)�H�g�oX��֧�n3�N��rWAd�<��8�����ԮsU�uB�������oUĎ���UU$����1���G.���9ή�HZ����P	fU�D�.�&���m�j��ϱ1�k{���R�<���3�7@��c�i��ƈ��ձ#w/���M-�8�Uq����|�M5��!����O��]��?��\����z9�}^��;�=D����̺�ϐ'k���0��lB��[��~�v��*zN�ٟ$rⴱ~��ꘉ�}�^;w��s��ҡB�Ս|a{r��<Ҥ̓u�NI������]��̭����;��;l�����v>��3����v2u��r2�^�!
�uu,}���\�hv%��ۺ9�AV6&����w>G����'f@����*��ݾ]�]Y1�aPm�>g�0�n���V����Enʹ��%!�z}nz�F�Q�+��\�uhD�Ў"��~n����/�M�tp1������G�Ll{l���b|n�**����BZ�;�܂EU�f�TuT�5��C�Y�DȈ�b;n4�Ee��Eۉ]�a�d�l�f^,ٻ!���h������X;�oi�;-�w���'��fj�k#�l�[�ק����Rn�3�Vϻڡ�8m�6"�Y��^�b���_O[g���8��Kv�x#�M���0�d8��x���^U������p�˻�[F�X�'~������̭��3�~#��԰�e��²g^>���u�9s"&�W�g^����!r-*v���z��Y٥�{��L2t�k�uy�|w���|��r��N�z��$���N8�*g+-�=|��	]Q�=v>Pޡ�Oiq�v��-憫����[����t����ÒO�3R��l��Xo/ �1{�bK����ΧZ��u�t��@vE�.J�%Γ��·��'�r��\9����4�E�õ�9?�^}���D{�e���������)����\�e���De%ϗ9Q��w"�7ks�f�mGnڛ6�o��S�Ya�HGѬ�[^���M��N9��T��el�#�f!j�(�ɦ�;��p��6��6"���l�㜸~��X;'V��=�� ll��v�JD���sY���o̆̾Ķ 9��]t����m�ki>�dY[e5rF|�*�?Ww%�%u�'2Tn���U��ik����~rC�� �үB�.=�k��D��Z9j��f���+=1��&�E�7	A�hm��b��,��~ؘ��Qtǣ<7�KV,5�'K�w�kӷ�*i���)�aۅ��^�u��B �Rz;8ш��^�l���m旊��ŌI�X��B�I��g���[����@�f�M��r��5�)�ɃNE�ʵ^\���"� +ډ�td�+�y���8�X�\�z�4)Ē)5vMkdά���Vج�`�Yj[y>D#�'��n��=��y�IW�bA
�I�J%��_N�l�b𰮙�v�%hSl�1�%%����Oz����LZ��=�"�^Õ�CB�t��ʬOr	K�"�s�9qn�;���rJ���vݞ��\�ݏ�U��,\��}M�2 ��7ua�����kn`�cޭ�4�$h��-�u6�p��-�(�+N�;a��7Y{֐O`��\K�\;=�k�$^��x����3oH~M����]�X3��OqLh2#"���2�n���%��3K���@�}��H��G�T�d5���<٫����͹8�#\��dH�=6�۩o��2�ݠ�2���d<d'OS�5;�9cԉ�yݹ� �6����3�|Ay�v�%�[��s�m�<:Z�^�r��+a���r#_8�'��og�V�kֺ��Zԕ��[��"�=���h�U������}mu�*�tE笇�Xuߎ�)u�#H����S�'n�}W�u�-����YB��K[��k�Eu{0,��Ժ|����Z(0v�]�E��ǃU5rOu���_�\�g�r�f8-y�Q�]���#� �8@����d��~hn^��y�b� ��i��ch
�f��U�g7	�*����N�4\�պ\	�q����J�<����We-�-�r����H�0@S�`�\���< ��-C���)¢�R�9�T��e��W6C�j�:� G:�)W�^��60T���t��w{~	^Z�d�qܹ$����+�z닇�+6ym�F��)8���\�՜2����s`��vDR�"�.�Q젹�j���m�EHyλUֶ�(�@/+2�(%�ft��&^��uc�ۛd�Tl֭Ĉ�U�|��Mҩ��t'*�Au��:��zὝ�e1q:�z��A�7�U��9���3�;јV5`����Hz��K&�������Q��	@_%nWl��ҩ�n�ԫ����ZU��P�WT�/-n����|Q���]����0���ݤ�ZU��1�`���3�����im�Ձ�����G8a@Yϑ��b ��n�q4��f9�Cz����D��N�֧��QZQ;1>�ۆ�ӳi4��̩�'��Fz��J�\\f�,�.\:���9ף��c���jݭr�U�Z��+���B��W׌t�;�ɁֵJ�[�J�sZ�qS@˺BvpHS#��&*�Or�G�
\mO��xلw2v��70���r�}{��+�͟$:K��ω0���i�N�X�
�Ogl!"�ۏ�ֵH���6����;��:��Y��ǻ�WG���R�Y��v�]	���&�9{���FA�d2�5@1  ���h��\.�1xh�&��n�R�;CY�Z��sƌ˗[iV=m�Lxc�𢨭�FQ��v*֜BJ��MfR�}S�Τcῥ/���![R𯸦���R� 3�'7ob�ba4q�^��?�V����N���� Bm�y%X\��l3� �$	R]��v��p�2��[,X��S� ��a<��:�dE�u(�@4�.�7�B�Y��t皌�PEn��m�V~amq�I���)#btM���˼��6�����kdK�xSz'VlVt,�h�q�t�5y���ƣ�3���h�9�d��l�i��v��u�L�n���-�6��Y�Zu����a*�nԹ]���p-�]1f(E9�]�A�8�<F�s�ΐ��wY�����$�y���)��3�� ה�՗��Y�O�rt3�L2oR2�]�G�O�Yc��2亝#���\]wGML(���'~�0��|0�kCf�7�loZ�M�E�C�r��%-S��:��@Ս#J��b5�ۨ�J���%(u����֍�f�{����\�G�&_ֳ {.�|��/��(e)̉w�jI��v� ��L�6�"��=�!�e��v�"�L�J����V0�C�;l_W$�%Y��`l��Am]��p��h����ݫ�۴~��g�h�Gf8p��[|��@�Z�4�E!BQ@> 1!�*w
���z��R"���H�4P=A�
�R�W�{�u4	I�IC�4 w4�9oMR	��H��
H��]BhB��A��)�"-��'��t!Z]#T P!HMi��P��r(tSBk@u�9�\W�=ATR��Q^`t�5�@�$�@�4���R:�!k�4,A@\ǈ9.H�*J��(")�H4�D�A99���/$(��Դhhu�hh"@�B�hB�:�%SCH�T����<���c�Ͽ9���������#t��9�C�v�F:�{��)mm
���)�q�*躏N;���oF�$���]���^��)u�od�o7:�(H��$3'|��b/=�5��<�����J��0�����fl�8oM�eN�>Ìh�|�:HǷą�Er��w��;��c�fv��K��~l{�B��h�=}��!��N���z�v��Ew,e�-
l�ɷ��[ �@J�����e�/7��F15��*�v�o]�Ք,�\�i�I��E�R�;[.cjbګ'�3�R�Zhd����* }ӱ�Oܫ/���P���,]Q�=��6"�.�l�BY���j�;68I��.��ql~��y���L��b��.jrƧz�W�`���gO�c��x�e��2M6��kz�Y��㺳�L3m>��ki���KX��4��S��!�!��,�*l=q��˖Jw�u7mGj���Foú�Y� ����n�ޟW��o��O)k���`�ISKT���M����ܠ�6��x�R���l��UVtɗ�wb�0��^����/�������W;��}KϠ';��z�S)���V�o�ɪ^��尞P��)�'r�%wT�J�����!�+7��t]�i��tj�^θ�ne�<+����1���x��qP-m���E�i׶-+�V�rpV��C�Qyw��r��yH6�K��rJ�M]Y�ur��fHJ��|I_]�anH|�;X�_��̕Y��.�v���[�!m��Mə���hf4&"�t�w�ݳ�*��'2�:X�3-ѡ�Z�H@�K;�7\]�U�''H��ɮ������'&���o*����]�lMw-��{h؇[6'+K�;@�gDf�wXd����o��9Kt�d����|q��u�O�cZ���D���-O����=�+��IF{i���)���U4�z��9�u����}��\m����W�	��"��6���ī�"��fl����h�F�3��x8�� ��t���xk���y�A��'���s+��8YT��}��s�6����>��/��Q�\���u�K�T�Tk��O�&�k;���t�L��n{ژ^~�x�%�wڞm�G��:�.G�e�ܞ�Փ�2X�6���Y�1rR��3ASm��;���ӌ���uu�<��b=x������b�F�U��+�Љ[�s�{��,{-m�o;���Wj�)P1m5�r����`�G�u�n��s�9e�(p�M��k�؁���;��5��w$�k����Yy�7-#{NT%�9�8a�쓘~�"1��O��d��5/����·��pb����2d6�uJL��yq�.��X���4S�r���f�6ԁx^w��3B�ӛ���e�j��v��s+!������֠��&���w7�r��Ժ'��9�[����cn��R�vCz�:ԇ8
��70f'f���\��=t�U��g�Gw���~�E�O/r���Kl5P���Ӂ�B��Wn��[l�I�|�{>��9z��U�)v,�*{j`�X�_�����ȗR/j�k�2Ǹ*㦽�
}�������ۉ�r���[I:x�3
��H5ٻ\��z��z�قvE��M�rF|��ҷx��ՎГ���!��s��yGi}�w��ﶄp]>��e��$L�������J3� �+�;�V�����^3lB�H��ʸJ��,�� 8�^��EC{�G�0[�-p4��l+���˕}���k����u �D�|��kO��hh%���f�ƙ�'*v�dְ���z̷k�Aou����!�����,�L�}�K�цL�n��l���a�*Pӷ�z9��Z�>�dG.5�*E���=.̮�;�gn=T6^��im��n��ح�x�0����}�	�(Г�M���1C)����+[zg#��9d��x�}�ue��ϵn�F��ᴴ[�mG�ڞ�M��v��GG�E�+mey.{�m07�'x�>� >���úm�]V	zj��銡.��Z�LfnSj��iQoیo�"ƙ�p�]bUu>���j��r���`+2.Z�@ձo݇��
�4A�ۗ���9���$��+�\ߨK����gβrx�,3Sؾ�m��)�y����q�;��l��~����T��Q��ŋ����4�M��˗J�e"�m�׸t�x�}� rU�s�P��N�z�o�������~/��6�e)[7�����f�c,������CnA(�%���-�z�sb���H��`���7��]��:����$�v�����5#X�F�Rĉ����lRq��	c (�R��ZM^��H?���*
��}�V�"�팱�������V-V�O�ݭ��HXC{��ޭ�Vћ�nE�8��x̾26�Pp͙��o�y;�: �b^n�A��S}~�178��PₑJ��.���m[��o&沖]��N�f�ܞ�=L"K]G28�H�R��#�e��u��-����=-�{hDY驤�e����`�Y�%���ѐڗrTzZj��� �b���7�S�VA��묑�W��{�)��Ej�79�d��2g�n�}�����Ih6��),��7WHwk2-��h�'6��W�g��\I��S�L<��ʓ�nːJ��~��ݐˠ�Yw[5YO�b#F��N�[�l̍��=eB���[�B�Sf�qh;LF�j�e�v�xwGE����'����uWr��f5�x���3�j�'ʮ�qW�F�e�V�	�/!۳��`I�1Fc���)�e��e�O^����)F_nCh�*�y��e���-�ǹ�
�z�����*����\�gO�#��\F`�������)��/��KXea���r�WȮVT��U����^��hj:��G�2�]-df�Q̸Ira�� �s�ە�����Y�\���1r±�.:���e<��C���Q�U��X����z8V�?��w_u�������o�4����Ѣ�H�l2�73�U��.mG=&�{��+.tu�������E�	Rk��x�|�̃�k�u����t�f	����C��F �ɉ��KRD\���N��.1C����m���φ/���E��o�r�?gN`i�P(YO�+eF^��7u[�&T[�3�r�e��i�J�O&����WB�V���:��R��0[f�a��Ut}ۓ7��S.���5�e�)��>�g�hg�۝�v�J[�����SEΊsJ̪	cE[-��ƚk�4z��®�T��纖iP��=e�����/	c(�Qڹ�mH��d���b��ק��D���r�y��}�+s�����*��ݲ�WN`�u(�n��Hnm\�jy�[���G0]��y���
�d(m��Ĳ'��ܐ�����V^,|�~"�ߛm���@iE�LŴ�t	�y�N��l�)����s*�Vj��8�Uc��ak��F���z@�BEc �������nV�B���:�셍I+�ϐZ�^c���+�;f�*���9O-��RB ��Ô�N��h�.�8������È��}=��o��U��6��iR�~����vҜ��f�R��ƅІ�yg��c�Η�{�x�M|xK/���s]ow�>F:��M��V�ٚblb/���5��͕o��U�7�0�m�;X7`���WO���]uA���@u�oU_ld.s[8w��q՝cnQ^V?����� s�*l�a5���7��z`�Dȳ�'��N����������ʖ]��n6�ֳ�����Y�Q_��N�$��];�[�p1��g�/`N���p���J��d6�H�sjbo���Y������H�V(�i�l���^fF��ꘐz�\f?�Gl5���`&ﲀ�Zk��᪝���[ෳy:^�S�r0�e��r���	����!�@��⮟$�q��m��M�~P������)��q#��^Su�PŎ���jzE�K;����j�Y��+~�%������T�̲;^Ҭ@���^�}�B�֪n�*�!AxM���Cۻݘ����B��J��C��ǘ$ܡ:�^7٘~Z��Z���љ�O�$�/S�y|�ˌٸ�*u��E����/��(��ζ@e�����=~�mZ�����e"�Hk��QY��7+��v���)��6�o��o�WDЎ���j��r���z�aTݗ-�[f�ut;����SVǟ�6�D�><��0�d���Q̸a�]Re��C��2�'m�xw��Uֻ@�}����u��O��以qh�Rn��[m����PڸΈx|7�G�+�cЂ��ͻR���Ljo���}�⼫}Fa�c<F�{�QVۈ��ĪX�K<�֥��fpقoH��w+�N�n�Y���Q1�ֱYŷ|���;�vե�@�-�H����rn%�uA�na�UZ�5N��]�i�Y��qŷ�ܫi�oNN�4}��&q�ݜҩ��t=1�����J��wQ�t�^�s��5?b���{5�Z�n�l��L�8��p��}�l������b=�iWB����G7e�س�d�������Ɣ�I���������5V�c$�s=e_2�����]�P;\463>.�M���Gv/��E��Wr����\�<'�]7a�Λjl0�4��Qni�vJ�`9�9��sj��wdOIau�Un��UR��T�Ot�'f��Ԏ3h6�h�}>~��"�!a����5�^�ȩ~Ʈ�J�p՚u�O]5�1�#xP�M&�i��6�=�j���M����Bj�e�m�<;����/���)�*��v���v[��
w^�;'l������]DBUK&ւ�=������g�/�����9�����&Q=n��4�5R�U֣7{�YPR)A�f&֥w2���c1����[�#r;�u�;��� j�e[�5�U6H���fu�)����a/3cT���������vfP޶ɼc2�e�#����V�%�.퇌j�̍���W��z�m�#ʪ�{�"���z^��������n2�w�ms4^TCw��ogV�ڢw$s��K�f���f@���*a��C�gSǃ�<�}�&n!a�{*���]+_�qfg��>�^��h�u�XJi�ѥ9$Ǧ�KkopP5C�7&�ۇ��k݃��g��y��:X�g�F�v�Cot:+F��;e��"�Z�o�o7��3m�%,�|���q�L[�t䭻���0;G:L�d����]�mڳE�-Θ��f=�����n0b6%���]�fd6���:��N;��%�H����4\C��ӐML:k��C7�S�3�P�𭘍�7rY`�4�7�]VW=*w�ױ��j ��-�1�lZg����7r�ϺtwR������ە�u�-��6�L����=���̻�=���@�J�W\�tln9y���3m��E����4�nyMD��2����2?�wU�U����^�p�2��֩��ݛܜ��Y�h7�$X��)c,����1C�f�0BT��|�?_��Y�@��𘛓Bы̘���䈹B�Jݠ#L<��عgډy0C��i.�{�k��uSܔ��vs�p$ׁ�JDd��X�1�ٹ����LT��wdv���k��ӱ3 =u,���E�ޥx/P)�$鈀L���{h��h�mvޮ��{[�*�����T����g�+�]-�=@P�@p͠އjh�#�a����۲2W�mc��8��oen0��J�f`P�!���-cJC����:gpX��É>���
m��fJ�)�q^��G�����=����zT�-"�0���R��;͗J��y�����rwQ�g'��$�8���Ϋ�*ی���'V5��G�gX.��͓]�p/�c�^$N�9P�=�x#E�B�*1���@7۹�Vɻ���D��d4��D�q�->�z��3&��BI���35$ ���#����.ʋZ��p��:&x���%#�Wz�<�r;��@)r�V>ːSۦ�,�&�����|�^�w�r��r:S���7v:k��cw݄0/�5���T-m,b�۠k��\����2���e�㘰#�s��V[c�sA���U�Tͳ)q��V�$o�r�����1Z��J�K��،�y��Q{���oo`RݣڣԂ��(��	�]�'E�%�+|��-ld��7dL5@�4��2��k�4�|��c��Ҹ�=�`ܕJ�t3X���
�Żbz�F`�O�4�Y�����r���K���%B�;�#`i��0�ࠒZ�_K������TQ�Yw�y��!����+D���]J��۩�V=Z��[�X��(�W�VjT�e���ͥ�N��U�e�F�Wx��h���ͱZj�t�C~�\sWaPL�pT��eeCj�
-ٕ��	��3�5��;����r�1H:�(��q��)p�=��y���?C��Vp$��9Zno���Trp��Sm:�u�Ė�(�/	3%�0�wKU�����C�U\���smd1k��l�Z74��y4>5p�K����tzy���YE���dz�Ya�x���D\xQ�+1����UbN�,�y�M�[H�X82t���ۥL����
a	�e������Ɨl�b#i���AS��Ww.
���gf>hܚ����*r�2��͸m��¹�1���>P����u�W֦���nʉ�{g!�j�����9���ZWj����.�w/�G!R�-���g����b��	�͗[���-��0����ش���m0,��+z���$��m�xwX�PIm�c"˖nM��3Ka��4�w���57��,eZ�{�<�(�mK9d�f��*�sY2<`�W)٦�H�Ig�C#���pqǭd��f��f��6����i��A:7�7ٹ��og۹I�����.���=��������-,�w�pr�a��*��\�sug��r��n9�ۺD��@�"�F �q�ܨ7����Eik��3l�:����ٖ��T*d�nd]y�t��u�ɧfq«`i����8wj�po.�'t,��K��ͻ�GY@-��a����m<A��6����6���AY��@i��$��M��ubF�C2���;��"g����q��e�E��3߯�u_]�|�5�4�`N{et'[�P&���C�B�J��9/�&�6´�u(4굥��JS�{��R�pD��>%�-PrЅ �)JT���4)�NN�� )ZF�����#B� ��ns��H�h)4!�t��TДT��Z�sj�Ѧ�(^�9̕A�BkJĮ�4�M"�@�R'*�G-(��t.��	�TR�!�@���(䩠(Ё����h\��#B����4�"PP��ǌ#��&��H�5����sϮ|^�.��\�WrK[gyᏕ]ŭr5�����oq�Tr��?�������{�a\�W�mdo�;�.�5�V��˓��;e3���?�R=zd��;<�b����*u�װ����W<��1$M;�fo���4�hSę��$��M`7Kv~���l�J��1�:nU绺�����驓�9\'8!��SrE[)[�� UՏң���1��c�YD�F�����L�Rd����ng*�B�@�Es�iV^^й$��I��5��懏��E�rd>ΑzD.2.6�U^�&$�%w�T�DCճ��^�=����~Ε��Wc��~L�� ��dm'������co�.o����t��Gv��-�����!��l�ZĨ��M�)��mŹ�iҢkI��|y_X�y�Lt�����G�c����h��6�*�Zs7qԴ�"�#^��I;�����=�hH#
��{ssM���c|�E��Н�+�D��on���M�@ܔFD�9�,����9�e�˪��7&�
�p�v4͋�۞*�pj�m>���{�1����(�84ޘ�Ń�Awb�~���^��^��3�a���ڥ��}�Ù��)�yġn��o�X��^Ͳ���F����.��ܻB�u�ss��"��gz�&!Y�
��rѳw{:�n�$B:M�w���h{����r�B�����ڙ���z~V�:��oN��'���[Y�f��|��vtGH��'˭�4�a���b�C٧�8�3��z�B5M�'zL��lR�:�����1ׇb�~��U�v���{|V!���E�@�������%@Z��f�BWuNsn۠��IS�"�5�j_�_p'����kd�o$7μ�C�d�, ��G������g�5�^7]���'7�t�}Xʆe��lr������݉��4Vt��;̶9�sL��V����M,�c�Ɏ�Z6]�w��WIDF�8>�9�w�殗�綎��>��j,�
��߷�{7�7WO�dJi����͕�{x��EwN��Sn%xC�o27֏_��9:����t+��X��r�f�&i��yn+�rt�ݗ^���I��gxWT=���T�)�t{(���<��[�����] ���wf;�$DtXi`̚��\/��n�CK��r9M^\3�N�$�d����͚�Z�;RM��g�>ܴ�ִy�ຓۙ��W_]���p=zc#��v���
������	a�Bۤ����vbXf�c�=ϭ6t�u6��^i�>3
}�3���-��{�m;ї�����S��I�܆KH�/U^�>yv�Z  ����ڲ�n�6	�i{�LY��r�sM��ܿ�5�2gSj��b`>ّY�}��e���K��`��������z{���F[�@v���,2.��,��Q|w&����LCԽ[��ōy���d�de�t6��j�EL��ۈ���R�\�<m��;�ݜ�x���h�-l�P=L��'=��/�s`����<�&c�����u�`m��.S\�}�׃���ƬhX���"���>��&��V*���D7]����Sq���f��(��&��i��VO̽���7���x��|L-�:�n���Tr�rl�i�VƼL��K<?4�HS[u#���=�k���mݴ�/-
��e����I霹4��W�oO�es1�a+�t=r��3���;5C��`]��2lg�˩�wlָlP,o�j�sh��U�UnI4�:���
(k�9Bk8�NڹKr�s�m��,�]����;�6Rܣzkk�T�+�hX�j�䶽�ݸ��X�4ݨ�݃�s�V���6A�`�]���gu\O�g�)����8����U�{�İ�͇�'U!5��7�4���K��K:�"�Cut��dv���[/~��SV��5�a��y�R����-�T={�9�+5��}ޣ!qUN&b����k%fWǶ
+|f�{���ب�~�m���YP��匢��Y�\gwc�n.<&�;q����y��Ԣ6�3z�������K?:������Pg���ꞝ�m�fǟ�o5(�u�*<��^\��o^5ǿ%�\��gʭ��U��g'M����t�#0p�_)�!8�K�M�w*�/;��Qb�O��:�l��pɅ����D�y��}��?�W������P�lS]�8�d����<,Bv��u��Ӈ�4ꎓ���+*��];���S��c-��O�G�9��<���2�f�u�=�#�fo�����i��xn��mV�7X���1ln���>R�Y�M[���9�͇���SxW�A���)����*��󄕹jGiո�Ŭ�}6<|���3��n�אef̡�2?�D9�ĸ^�V��F��vy�k��N<���)��2"n�ngH]���9'�)ׇ����pw��x��41.�ԫ�S��g��wSA�T�ҳ �P&��,p.{wcrrj���{�����V�ǆ��&D]�8�2'����"��t�;�w3���OW�����[EfU��1�Y�,�zU][t�B��{��6'� ���Y�J%�+�w���n���y�U�>J�R����g�/T�D �E�[½�WPnH��fh+aWVTq�]O���I���l�����K�dx �<F�u@u�u��\K%�lq1sV��P�q_�DH����Gޓ��o劢��>�.6���O݄�OeR�t�=ѡ�*���؊�Om�E�M�;���;,�
F�����v�ڱ�)kF�g���>��A����hLXT�:Hc�Z6fD����}�̄_�n�<H����uCL��7��޳u���
x��8h����:�"�9/�mhShwq֨���$h:85yNcs�S�"y����^^�08����.��]�f'�g}��[S�ERx����o�u�-���eB���]�B��M٭O,9��9FC���^�yg_��S=%[�����D�c���.��ΊB9�U���D���&����r�2�r��ح��d��/�����F'�zૡ]��y�OŤ��H,�k�����������'MF���Tel6���i�Y�D�*�Uى���׽'�Iʸ�|u�pO�툭�=����	�Gө�K��k-iX�����-DeE�]䝋�G	�L`���+4�+��4�CYc��T��E�!���9��=z���ż_�i�Hn������&��ڝ;��6��ᅉ��7ۛw����.����M���P76N^���JT-\cwTs}�k�
���	�ϖ.�4[��cY0Sd�!�֚w��R+6m[?�Зnj�y>x-�Ǥ��G��y-I3":+���T��'A���o�T���W�����V!���g;d��E��ݔ��ݤK������m�#Zլ���vyV�x7��T{m���D쓍���Xq1ܱJ���J�9S�1m�Mȯ(P��B����ok���p���%�a-�d?�s�W$Ath���i���\��ʦl�^O1S�Wڵz����$tT;�?%�M�@��C4��\�'��GwA��Ʒfy"i#~O+k�M��v
�on�0u׏<k����w4�7G�%
�x���z�|WrV˺q[l�4#����+AGά��~�<�V��{o	�)<yU��on�����-�n�X���:���gV�6����t��"![�Gv��m��y�\�1�Fq�w�����"TVz�>�dXbW�}�%`��;�� N[^=iWk#.�v�K�I	�ō�k�27\�l��B�YąfFq�[\�ԯ�޳x& _f3��yW��som��)c!�������B�1e0;
�$E�nK��w4jq�4-!8�H�(dnt�M&����]��u�%|���e"#k�J�G՚3Z��ɴ8�F�+3M��$� �������M��U"���vz�k>n��v��ˏ��b���(���az�(wl˼�Ց�³�Yu)������&�;��nڠW=�n���Φ4�{4�#[�K��1un�ɾ����ἄ�΁��󚉚)�+�u�G��2��Ú�-�\ַ�����4�y��Jv�EȮ@��]�VN=��b\���;sd�������M[��^�W ��u���q@�(7��y�jj��Qv�i�5���g~�몈J�JEU7RʎM�-T�:��.�����Z�+�)��[+kv�frG�A+Ǽe8��dj��l�5��}����Nh�~>n�Ü�T��&���utO��O���؞cYN���s��y�A�0D��zh�(�ˍ�:�˶W�yַt������A(��y�0��ssn�B�~����9C����4��ʀJ��֍�!n.Ta\���z�I���}�G�\AޯLl{sZ�޲��H`*_�v��{��^�;E�,djlR���\]�,z�j�o���[��TcBM�+�)x��l1u���>���>���l� �{)�M\��i�����\<���l���5Wt�AzX�33+ч��]��w����f*�j��dwN�ތ�]I>q���e�
�uR�չSrU�KAu��������cx�e�����d�BĎC3�w��ĪNXk�ל�4�j�����͇���Q~���s0����ח�3x[��m�8�VM��&#pq����an˹�wkIɸڬ�i���?a�T*�[�n�����r�L�z�l6t�&�`�*�k^^�tv��a�gdB%VQ}�:q�Cq�H�f	R��YUEk������^_�o����}�t�����OUZ1��󺈐�:B��^\4P}��uZ���H�ȫ��!௩_|�S�.�`p�ؔT�:���_H��h� �z���� RF�5�ܯ:nʘ�;#�]�.��y^[�6^�e�S��pmw5�IH�Bԝ���W�ɐ-S����ݰS����N�2O���{�Rn����9˷��5�*��Ve%m�l�X�mO��L��}��8tpih0��kUn��2�G
;���O2�~��j�~Lu�g��&J]��J��꼥��{�3�$ȇ��T{�ͦU.��j�,�.P=aMB�CJ���y�7$���5��~M����#4�fզ�dc��u��]�u+�Vɤ�T\���yD�[g*m�ɏd��+��qg30ɍ�1��~t]�^�~�����r]��"�1��Vd��D_H�˷�+k���x��M��όV؂4��ێ���\�LM�,��%�kI�H�կQq+s�^�nr�^KזtC��
��Eǆ�T�h�6Xf�R�Wdf�އ�����z|N���	��M�c3��e�"�oj�P�CC�)���&<Au}U�1���̢Ve��}8E6��n��{}��g��&8;[�/�t�E�Zz������ֲ��x�t����������hT%���:ψ=H��hj0�dRI�M]i�dn}�� �7p\�� �_���p³�^��p�hQ} @J(WG���onî��/����M7���I��\C9Ά�ӭ��
��������npCa��W{����[��kxP�	��c�ϫϮ���{��[��������/���@���
���UQ�A�_�Lq�N��sv"`��U�s `�  �  �  �  �  �  �  �  �;� :@	G�\ �(�X`�@ �  �  �  �  �  �  �B $@!@9���  A  A A  A
 A  A( A���RdU`�  �  �  �  �  �  �  �  �  �`� �   �  +�A�0����+��A�*�"�
��`��������	��� ���0A�_���:�&|__�@�H%(���&�������W�����3�?�����>?��ƿ
�x�����������O�����?ˠ����~���g����/�� *+��O�����?P �+���0`E$G�~��)�	�0���:��נ�)�@Q_���~j)���~�D�Q�I��h�Op�z}���7���R}vk��Dz�L  � B   Ѐ��0�H @ H ��� ( H@ � ��@  R   R "�1"�c(����I���v���QO��?��
�
P
P
P
P�zQO�~��~/���S�O�����v/������#�(��. ��;��~������8���/!?�����z@Ex�Z��~���_A��Q_P *+���	~��������`ADW�֟09�@}Ĕ���q��}/`q,�yܛ���:��:N	Н ���������@E~����������yO�?0������'�p�*+���������-
�B "J���(� R����* �J
Ҁ� �(�H�Ъ4 -�B�ЃB(�"��-+B�Ҩ� H*�
4�- Ҁ4��
+B� �"�H�(�H�P!@
R*+H
�(� J�(�B��"
P��@
Ҁ�� H��*��BP�*R� ҍ(�(�%J#J�(J4H�H�#C@*�@'�N�S��}�S%/ڇ�����>���FOq�ۉ������O����v�
���"�$��{p�_fĞ��'�I���{����P�_���vq;� �+�����gܙO�?g����o��PVI��p���������@���y�d���0f��*)J��Q)PI$�JTP/�hQUT$�I ��T�/lUR�)�>��D�DT�J����@"T��JG��`��)b�*�m��1��)f����T8��`�6Mm�m�n���vݰ�Z[
��QUp���ѕ)���kl�ʶ[U���lZ����R�6.d�M�#%��ml�6Ue��ReZ�������V[YYd��M�J�[[[e��%UT�ۍ6�Q�V�ֵ�ƶX��C6(�UK��)v`ٶj5�-���̊��) �:����e�E�%K�u�Dѭb��;e��n[��ض��sR)K�N�ɧje��v5vn��40����j�ڌ�Ћ7ֳsQ�����m��Slֳ4�JͲə�	S �H�*�
  E=�2�*HѦ����hb0#B)���A��1�� (��4�#M Sʞ�	�=M=LCƩ��"��	JUi�L���d�a2d��hU3S�=Th�     �����4�=OS4d�� 20�e�g>�o�G=&�-}*
���M�!@M��"�Ew��QZ�@�@J�D�x�I>L|��_�Q�?�t�0A�Q!�L>r��	�(Q!J�)XI�	�E@K������j}z��O�*�a(V�.V"R��L��7����G	{$����1�:�*�g��WS�D�a	���V���w���⻭��.�Z�SC����
���.��XY�I]fk51&iLA�D%��J�m	�-Q�*jF� �%(v��kKOE*�Go	[r���f\7M�U��FfYv2jR՚��T��U��дIj��$T�<[���n��[%X���Mb�2e������!n��ܕh����d�Z��IP��ےj�FJ
n�(^^�%�.e�aZ���g$)�m���kj44�*ս�JQ�e;t�u�l�嶝����������&��32��X�����A��uYr��P�,/�8�l����+vҠ�ge&B��{��.�oax��TЎ���M�%$ͭcq,T6�kVCJ�}��*!,f<:�v�ChcbdZ��on�J�\2�9&�*[ճ��Z�xion���P���pACN�&B Z֕e�@0����r*���UZw҃z�6�ѫ#	'>��� Z��Q��; ͬ���W��v�iaDE�'�YBL�H�T�c$pU�ݖZ�Jx��0�8>��t>7L=�AΧ[n�Y��E,��l���dXN���i����J��y����d�N�ǆiBT�� 76��(A��D�ʁ��	l�̨4�YsA7����G2��V�b�P�shf&����+[˔���	GU�% �4h�kChS��S���F���4�oV�dJ4ܳ��kOr��Q��Xۛ� ٮ��v�H�F�c�A�!�Q�����̘��`��b�<ʀd��Ci��#Sv��DU5&��C̧r���RQ�!z@�j����-��l����ư�cwu��@����sA (�(�ݼH��z�ǫ"�t��Uf\YNj��,���s5�I��Jb��ta.�^Sъ��VѺ�ue�Y	MР1���d�x�a�WsL�n��P�Gk)h�2�!N��Đ\2�ۼyN�G0�Vj��ꪋ���6]Z��
î�iі��e��S�̓4�o��0�DZ�Q6b���ܷKI^ᦂ�ӵ�1$r�st����6�P�dڔK*���
Xs6��d�!O��G'R.Ƣ�P��C��J�Wlϭ(�Ow! ����A��fd'b���J�.:�2]8��MfY���KM��)Apmg�;���z�^]�����P6N�ebrk�����&�Ί�zn�lh��'w���ϕf��h-��&4���!�T�Q��1ͱ{p��xm7���M�6U8o@bT��Y�SX�B��D��1l�6$r�C���-��w0é��Z��Լ�i�8��3EL6� _�[30���+�Lx�ϭ�0����j��2��s(�Z��BJ�u��ņ��w*+��[V�(CNj1���,�4���V�Жd�1^�"��������S̭V>{��tB��r"���=�Sl]�S��Lf��flG�D{�f�ƌ��A�O@9�g��㡴sdd�[r�W��gE
k�,͌�����ea���*��;�o"նMӸn#�d�=F��X�[He,_$F�5��U2ƺ�(��1�f^���v��gЀ�R@|qj��,�9�՘�(�Y�*\��8��6ŀ��kf�'0G>U�ݦ�q�З�ɼӮ�)�ooc��9���`Ѥ`a,Y%�kE��0@p*�[R�F��q˧����Eֽ�T�T�F\u�	�Յr���c )(���Pn���[L����9�c�D�B\3����Ŷ����Qb��
Ɵ�HfJ��6��źp�4�u��z�j��^l
ԔN3���qblޝ��"N-0��,Xu���h��⽠���AjƖ3Və��L�5yP&(@�j���MۡO�wF�l�ۼ�./�4�L�[#�>���cu	V͖A��E2.􁛚�E�ƘYS�h�"��C�Ţa #v����r��Pm�x����e,�bT�h�d�t!�Ycq�&�X�b���Fp2[��[Sv[+iXu�3J���3Xvҫx]��k�$6��9�nd6� �IR�ڷq:6oE�-�/L�^)m7��˱�Ӹ�Rl*�ө�ƕҭ����o{R�uygoR��ݱ��(Se��ݫT�Ȱ}�$�%�ş�RQSZU��DK�hۭH�Z�b�"k)���/ZzD�嗪ѣ3���Ɋ+P���#R�e�2$�C(d���KF�B�ckn�2�iح�%�4մ�(\�ִC����P�LH�B�Aɷ���Æ�A�`zݰ�m�e�,��)-D�q�tHE�f�V�{���_�����K3���!��
4	Aߞg��fc��:��k�+����U�bn�w<	_w)���U��Ɨ)!5�eJ��ᚲ�݊��"�SO��2T����J}�΢�5�#Q1X�Y�#��qP�Q�k�G:����}%�QYt�+��N#z��w��TRܔ�rc@sv=����}V-�dU��n�NJ�Ԩhe�ݝ&69�i�W7��2�콭��F���4�t?��V����:��u����p��/w;��2l�xȆO������RէT7��\.��ӣ�b��<"�E:�klf��RS�I��m�Z�҆���y��:�plK��[㧅��Q�F���_v.w�@F�q5
�GR,���Ys]�X�,�Gb���:�����gT�E��*�\��"]�OÍq"N���[����wu�_:&�D{E�E����э��%�U�LϺ�̶�$��%<�+�Ԃ���Z%k�M�ش���m�����5�]-8&퉎�%z!�7Hnu8;��K�ܜ��(t��r��ѩO�T��@����Z�gN���.m7����$*�%�vrט$�[���!vY#0w�-˹x1Z�s:��E������B�S ݇[%H�f�C�šP�=�4��q�X&�e���59s����@����5�e�t[F��X�Z3��m.�=�aԘ/���ks�XAU�c9Q;F��WP#FL׹�p���kJ��H��rBIE��{��C�ک��S��I�9N	�6CD�d*���UK�·S�Lv��Ζb)�;�q��7���rp�M\���;V��8R��&�.��U�1}9m�lQT.�*V)5��g��ܻ�g�,T�/�<��)x�t9�PC!AemN�_^���L�9�7�hQq����Y��@�<���O$�}٠���1�I�!m���Γ\��2gs�S2�e�$vmunV�����Q���q!��W�m�������gn��p����J@�9�J���ѝܦ�;������qߊ�Lz�}����R� {� �q����7�4P�j��ӗ�E�i.l+K�:��S%cN�O��0Lzë^�[�^EX�v��vVe"6J���zO����|]��i��g=���uD�S%p��v��h����X��w�JY���6u@�$����)�o-�K�:�{���0��R���68e������X��{t���`%���i^��4��*p��f.sF�kR��Wn����Aˁt��y�.�L�uT�4���=@�\Ux)`�T�K[��|%зv�1�rJ��%"Wcͽ�2�s}egD{��G]���oz�[��P�ű��}pwP7�f�^n�rG��517[tn>�������EIb���i�7�c�x��:l؁ޭ�7�ƅ��(�'��U�_}�a�+���@�.�Fr�/����$��P�`ݮ�F�C�M�a��Řd�]��D��Wbѧ9Z+�Fm�]p���G���B��{�ze!9��t-���	�U����yA�_۶�i[�ӯ���ki�W%]�v��ʳǭ awJ�2�ĬQ6���y#1�N��X��Z˝Y�~G�D��� ��md6u��yJ��Ne��L���7��n��濤�u�0�Ʋ���6K�h�����4�V���Ք��{�:�;Z����5���{��x�ol��i]��,�c2Iu,G�6�]�]$��hKrQ������i�c&��U�]��L�W&���D<�U�@\�Tv�� �s�wl:r� a��v�	ޙ�=o%-�s3(B���]�8��(���֎:�u�;a���y�@��~+Sm��ѽٴ�ۃ"�m��_��E��|���@���;�{ҹ�3�+E����0��hi%���J��]�FZ�����F�"��ջNX��yق�����4&U��h�Mf�w+�Ur�v��1�CF�$R�r��lõw�3s���HGu��l�����Ʊ��0bL��H�v���{�Wb�kB�x�vw�0Ȥe��c�X=���)�s
'�c�VU�/u�E�.�x0�|;�ɛcN�[�c�*.iѬ�i���oU�7,v掸r::2�֫HmgMÑ��������2��=]Ykl�E��tB��%�Y��U��!��b�JY
��.K+�U�"���(|��LOuu-w�|�	��-��J�9}��u`���<7(OH޻ݾZޤ���I$�I$�I$�I$�P��*�Pd(GUL�e���������p��7��9�ĸ�훻�t-�1�r�6�[���6ikαWF��tW;3��q�F�'�Ç�7=2�[:{��*I�ve`��ǷţfJ0H��F�.;��Uu�UJT��%S��F�ՏEP- AJ�԰�(&�ފ�ζN��U@P��C��n�]_�p�?��s���N�nqv��ZN>و�UPB,��4S��ګYR�9ӡ\ug��a%<�������!>��ʷn'���5�$��� {ۄ����'s���u:ޗ������M�WY�hc�Ʈ�5�
���U�O�ow~�)F���vݮ9�qU�͆�nV�mvHp�U��J�:(����%.�GC��Y�U����xA�������Tk��q�0��E�+�����"��(��KEYHM�hi��j�� ۸��u�Դ�:�C�a�r�V�A��0b���n�]L�K
�ʨ�<eL�
�^�oc,e-6`%�o��.�Π���+�\o.��:���>�#9@H���a��s���݋�F�bL��r���_��E|�d����_` ����m+;γ���o%�v��x��\w8���K,F�j
�X�I�>+��)�!����6�VG{m�K���WmL������Oi�["�9��4۽v�����VT�·S�X;"�2���iJ�>���9�bK��yғ��i�G&�w2��U�1r��K)k�ם*�&�X�ä᝔��f�w<'��)fjW]ALS��V����0�ӣ,�hj|��<Аw2��<�m�6�e�3CӋ.�Ņ.B�ӓ6��h/�W	���ݢ%�6�w.�Q�Ws٭�4#��{WJn�*�{��˶����R��u5�fh�:|WV���\Y����
4�\��l5/qB6��Ԇ���63��J����s­��oy\�.��7Q�qb�'Q��Pqta8��gEw�W�6m�Ứ=�5��[{��[8�'K�'YR������J=;l�4�+E�5��9��ϸ��ň^�]S5v�@+}Cq;���f���УM�P��t�,�I�R�Ҷ�yZ����WZ���y{Q�RGE��(�1+t�ʓ-�L�`]���+D��vy��}�p�uk�ݴ�f��2���[˻��u��{��~�˯5���C63*M�R�䀫�5�XV�W��f1�n7:�#�]���0{z�c@�=�J��x�yt^�u�*���CX�$i�s�+�U$B�Gr�@܉��5p����ʄAb�Ձ���a�.a,�{�г�)s.��
|*^�e(�֞���$��V��WF'�c�����р6^h�²�slҴrc�����)�{������};�9����YEL[�A��/R�s��,ͮ��l�[4kk����ZQ�(;{���^l��v�7"���d�kGqLvJO���T:̺�X�Ֆ�B�1�u�ln^��M֝3�FMY:*�o1�ݺ<r�\t�y\8�ܢhu(��Vعt2�m��bMɫ�>}(�������[�ȎrAXt�[v������B`�[ѕsyZ`Q�-V���6|���ECzD���2�K]�R���S\ `9a����a�4p��ќ�t�;˕֭(�7#���ݜn��P����J'�.��rVU;��s:V.�R1,蕠&���(�x[mڳ��vu� ��C �|�����l�osC�������|:��z.�6�u���S �k����u�@�.�D+�����P�H::�����9}a
�О8�'V\6jݴهg+%�����+���n;�T�'HM����g,c�u �K'��N��^��.��5�s����ov�t��e��n�$T��a��x��,�c�&�nD�.���B�f��;MS@4��Ьr�֘6��:&��(N	��9#�,AEv���d<@1�6�ʾD�W6�4Z��wY��f1��H`iѤ�
!ʉlǣS�&�,j���Q�ٽ�³�v�c-�O�H��u85:�hTf�n%���!4�2���v�+�A(���5K��.ł��D�ٛ.�=o�W��\��v|��ਪ�:�רK7׭i ��8�J��B�����U�y�Yk��=;c6�.�w]�챜U!@L���g�K(p{��ۤщ�On�����8���Д�f<DPf�Ə�0۹�֖���C�ł�-:��tm�w ��7k��ú��g&��*Z�/]�;1�mu��t��H�"4�����9u�����qu_�Nٜe��]�P6%5���awר�8l$5�[x�j�]^����J�������j�J�*ݨ��<,_4��˽��]v^�t�G��3�V��ur����E�	�5��v���(��U����&ɍ��j�	�١�ofAC~q��^�FT.��$(f��k:�fw��L|@|��� �P�xD�
9�=ّ�;���>3�q6�u�c_.�]d:��bՔ�m]M���z�I�ְ��^��зh�
�حŷAҤ���YZ��-S0#����~7}p˶�R-";�d��*ڱ�k$<�P`'#e�%MF��4�8�v���ae�֊'9>�7��Z�����q��LPݵi�n3J��맩����o��ܼ����S�������7z����x���Վ�[�%4�RA�`M&X#(De"�)
��a@PX��
Ae)9�	B2�
@�K*1K��� �'RAS1,Di�g�)c3��t�<�1y]CgWr��S0��g<����5�+��]��<0gV�r_W.^�'�WPIQ/
�!S�1͊�kw�i�%�J��zߣa�����t_t{%8�X9�f�O��wC���RO[��/zQ��t ݦp���u*Oʱ�9����J�~D�,�ƭP->��f�)Z�(�eu��m�;ݿ]��*G^��4px�����4�oQB�V���۪S9�m{�ː� 
���Ԟ����%�KW � ]��� t�n0 ��j{>�"�kV�y�iN������^�Ķ��`��7�Ν�p_F�����.l�[������ձ���f�tR�*jaU��7�|�a��Y�p�*��ո���0/Z3W�P5'�o��Z�m��"����^w��[
.�k�H�e aSn���֗��E��^��pVD_��z��oud�p1@���(�2ρի1I8R��έP�LVa�fC��^����3��<�j��:�ꋚ���}���GkX��i]⹋�#q[�1E������2/��SrSoi��lV�V�6�en�����ݶ��0�С{*�+[@7�<�[�5�OV�Vn�qZ�kw�A˯�?P#���k,�]z�!7�����ʏ=�a{d��ӣ�D|�����Y���f::�x'
~%��x-Mv�h_]�D��y�o�}�^�8���7�r��#�"��]1<:צS&�LX��Ij½C�B��T��mի���]����9b�q��AyLʉnaA��ڲMԕ0ca	]�%9Y����H���Rh�΁�U��������nȉ1`Qtu��)�;�u5��cy�]���v�i[�ɭ�N_�.����I��<�1R��H�v�ÈK��M�/[��R���tޱ=�F�!7wH.Y�@�/		�Ő�厪�^b�٧���:��d!qZԌ���.�ȹ�Vlb|J�М�6%�f���h{�|��ڎ���cM�2�:����:�
���r��I`p�UK�{�4C���d��j�{��`�D.�,������~F��%�]�����׵�F��8�Nɟrbj��J� �}t��:�n�N<hRzD:�S��,y���5�o]�6��j���}��򤔲wxt�u<}���&�v���)��;�"6��[�wc�8�kYE�g��CiB�n�\�[non��=����5���o��p�-���!�ț��7�i�o{�^��J��]��-�l�X�S��x�m�9�M^P�*L{@>݆��A_��&b��MI����sf�Q��DV�=�) g��X�R�E�ioq�jCͿOmA�n�;}V�&���$�9��������fJF��뼀��:���.TY/I�\���S��G����k\��6b�0�oX��*�5ft瘷�"Y��]�^���	�ѿ�ՠj���s7�8�,{����!�n���5���&^4�SO_f>n3l�\��b��ѽ5�SY����`p�@F���
�e��7�X`{jp�pS�w��4�	����X_wt1���2W-/j����Y4�Cu�1%(z�[R|k��Z�Ӈt&^@��'�ІhM�_!z�>�(uV�o3m��푵��g�Cd�9�P�fA]���y�>���&��oG܇���0��:��lR��0��a�9��֛PS�$��<�H�/L[{������Y�|�Hx���N�{��7���H�m��3H��W@�}b�J�	q��i\
lӷ{��w��ׇJ�w� �b�u��4uN�]�Ȼ!ѐt��d�Y�f&���]�۞�h��u���Wvm�]d�Y�&�-�F2�`��ķ6�z'z���2�)Gs���w¶�u+����b�ǃ�<K} �)�m=Ivz��qwp:��a�^�;��:�;5_:4�����k��.��F��ƭ�����D�f��~D	 D~L|7���ߧ�oH�^
�=�R���ϥӺ�#�|z�I�e�/�^ �\��C�wW+�%7R�k�N@Q���)#�
��� ш]��c�`ܟZ�tiq[�P���y��6��xS�ځ齵��E�����j�u3�F�r7[�h+�	.�7�:�:픚�tN�=wl�������4�̼0�h�%+/'W�Y.�Wt+��k+�-��3�c-��	�|����_S�f��)M����ImB�b�9F�qa��㥊�~^�/ܧ~�C�Z�nAq~	:gv�i���a��ơ�mW շ�h�;,S^��iŵ�5�-S�qT�Č�GSŎ�mئ�J��J����h�9�A�z� D8��T����Y�l`k-v8݋6�^!���W�!KjB$�p����F��_Q��R�Gu��'#�+��E�Jևj�Ec���o�J���͔8�p�4�w��=7�:b�LTĭ�VB�'P�x���Y�3� ä�&]\�M��T��牁��9��]�����u8�t�C��9l����5��`:��H<�SK�� ��!%L���X�JHP�B�"&f�X��a�`P�J(�b)�b0��I���QHJ�ED��LS),F&bf%"�(�!�PX�E�޽o��q�g=^������QcK�k$/�ѹ�;�$���b�=�P�S��+0_��#bU�,��;�[�w�i}��%��i&�&���j�Bӯc�=���:^���V��,��ɗ|���}�����ff#��d�{6']�+H��+B2s�pm��v�]Tᵱ��N��b��O����̞��r���
��ۢ��������$E�`�àa��+y��5\�{��f�>��3����5Q�i+�]�I*��c%���S��x�Ś2�����k<��Ё����\$Z�|��ow�F�=��5�D���������K	8�z�'�B�@ep�ߜ�<) ���+�y��ގT�]�����|���Q�*xUN�1�g"�kJ*��Sy�T�>�� {�>������
c�'�)MĽ���P;����� c��iYt�D^@�uPd^��{>�)\��P��%MZ�~�q��D;�aI������&\q,�ԝ���\,�V�>�|�&7�[������.�x{��'�\Դ��7m�8�R��J��B����j�΅ܩ�ѫ���s��G�Y��}Ϟzo6�� }u�l���?��}UW��w3��py���:;�{���X���;Y���^S���Y��x%��N���W���f�u���m���,l��P���g���n�m0�������_ľWri����S�L��6�e��݁^���wEr���g�z�Ӑn-�����-�b�6/sC��QBWO��+8*
7�"���5BL���Ԭ�����]���ٯ{�VvA�N�"����uv�H�5����%Ժ샼�{V���LnϘ�<�M�����v�VM�,��{�E��7��t���Sgq�"�����7z�F��뤥]�"�yc!��{ũ�d�d�&�����G�����|���x�Cٗ�����^Y�)c�E�����j��eyO0-��3��W������f��\qw�|�[�{��ܚ���Ou�׺���s�/zs���"�Dh��5#�՘�<k��9��Ƞ�P��j�������0u�x���g���ߌ>�SC���&ҏ{8<$�1�<@#�QʳN&�eV$�'{�e]��7�����}�:���V��ś��e�ԖfܞJ`�L_�>^�O��ל�/f�@��2��q�z��U_UW��7�Ӈ�n����hj�d���L.�N���) ��`k��)�A�渉������ ��X�1Af�{���*��\��q�r�O�"AR�7h_���;�=�e?8�R�����7����>C5��q��s�C�Ր�Hv!7���0�w��&�%p[v�?7�����>��{�헐���O���r&��W��:��""k8��>�o{���}Y}ϵ��;���Z�4�[k��z㫎YP���{"Q�c)
��&&j��7���Dy�yҤ�M(��_nZ�D��zu�*|T,ד�89Ė.t���h��g�W�3���ṵ���uњ�W��B�v��_D����t�>�b��1T�Λ�����>$����Q�9K��}�%o��LILٻ ��>��菡���vr���ϯ���]�\!c�1���q�˒+
�-�ydMvT�j[��]؜?�t�Y�����h
WAW�큗徒�:S�Vb��y� We�4���l�>�}�R�˽6����ˮ��Ei��W=쁛`L�v���I3vC�w���fǇS�6�N,����[�y/��UW�DJ<�Cn���o��W�4�y�~)#�~L�O=��9^�#�u+KVy^��O�|��B��6�l�=G��!��xt{wS+�;RТy��)����tR����ƇGX���qZ���ߘ�WDkx��T).�ޝ=�4Y���W�,�?,�������b�fn)����6�ڝ6�86V>�����{�s�L�.��Au9��\���2��J��ЙMC�l�����M�j��y�zڭ7��������>R�y���,�(�fHvţ���7VϺΫ������-0MW��Lbx�Iͫ=��j0�4gL������I�z�EV)
��&u��z볘��Y���t]@S(t �� !�Z/2֢wr��*�-�cԀ-�Sd}IZˠ��y��?��AS�}��l����޲5�Ш�5G�h2)�x��X�*)%}2�[#�lI�eaC4��՗6_,چ����ᆹ9j����P ����Ȇ�QG^VU ��3���K)4P$�ܨ	�q)�8��u�&��)
��7�2wV�Q�vFRH[M
v�8��ˈ�v�g��U�j��ҩ�ӦXɪ�r���&�̨�`]B�n���4X�5U�J\Х�V[8�Ѿ�>]�<�����_�Ԍ�K
#31�ؤX�̙�Q�S$SI�"� H�3(�2
B�30ԋ�1H��gL��������E�)�,*$����V)	V��fdS3"�beE%�V%�SJ�R
D���05%0�
$}@QʱK�����g�A���Gy��cʻ��� �uX�f�5^���'�4�sR,qr^7��o�w#��/'[���O1}������q~s�G&H�*Fo^��u�}ۼc�&J[^����%��xS��{����[�k	m{a�u6h�u�VY�4�;wsj'_�[@�@�#2]F���٣Υ�`���S��C���r��I9�J̩o���n��.���"p��鲳f����T�8��Ϣ#���{��{*�s��4:��٭��q���y�6���P=h�s��M�/�S��(��Xo�Hvvw�/cR�:�?-$�o9����}�UnL�����X���������)�,���� s��zں���7�'�J�˵��'���9���m�cr��X�m�F%7�ą��m���(1���HFk%R����}�E��G��2�;S"B�ގ�8�W]�>K�dgrJ��Ϯ�הf�c�p������>Z�ƯXk�t}��T��Uɪ�r���iԺ6;X8hNs�PJ�7��Q��Gv+��r��FՊ�!��3�@�(�+L]>۞!�oq�Ƒ��G*�2�=�wm'�PK�w�y�t.��p$U��i�e�����������=�7�O�ok ���|ʫ�wma��]�EV�w��8荕��a�u�]��i�/�S����=�g��㛙Q湺�W
NdQ�y�b�����h!S�n�J��,��oe�Y���S=�AP����h�Q�!Ͱ��&��̯9����܌�� �;���`�ݸtV�ŕ�7I�J�[/�\n��u�������D}��i:���U�&z_��w�ZA��C2
�˝{F��^43j����v��fӆ�mH�o�ZX�7�1_�
xu��j'k[�k�A�@�ðu)����B��4*�=ܢ�z.�S�l���[�q�3O����y����M�������أӶ7����~W��I�r�R��<ƫL�6�a���W�T��!����;�����Q�ϝ\�k�m��n�.*��k��N�,�� �s�>��a���{<�Uf[�~S�w;R>�A��jD\�Tuq�9���<��P�ƌ�Ti���XҞ�����*.�%�;][y���;��7=X��D�5��R����U�=�9��_I���=5�������y��+�/����l�yx���o��g\�s��e���j�x'��ci
7X���w�rr����_�0�3���f�� �jg3���n��,�1سZX;5�}ȭ�7s��6q��p*h$�%Mw�u�1�����[ܕ��L�ڃfHc�0�F�G��zܝ�ry%��ؗ��Vr�z{�:Z|/�sy��-1.��E������韬~̖ħ����0�'�X�b�s "_s��<Zc���ݎX�gZ�F�ҷ_���$�gpʡn�����"�4�2��[���p�W�-n؝w$|kr	�=�* ����م,Eí�Z��c"��4���׽x\���Ï*7���A�Ő��Ì9�q��z.Y���Wm�5pƑ��t��}_f�?Q� ��W��F0����'�žZ.��ڕ��F��#`x���%���ts����盆tMJ"~1勽�z.����<��]D�'cW{B(F.��~�=�j=85�lw�v���;h1
���g7zfE~Yh�Cʮ�	�E��� ��ܧ�֡Ǟ6���k���d=+3��s��87GIj�����r����U��~�댑�{�v�n�)�'���#�Vn���68���'U{�N�������G�s�,��jf��5��o7�p c-��T��y��*�����e#��{-�F�i[�ͰK�������滵L˝.�_=��y�y�:�w�Я*<s9�)�T�H,�A���WY�Rl�)92�:�pu��Kp4�ݽX����J.I4v���u^�T%����5�]��kwu(a��d�9����v�W� �Tr�ևu�ռ���z�ME>띔����醘��ڝx��������f������<wGi�7�6)�Vn���� g"� g](�㔾]��*>[Ksf�Zz�D�KVM��,��)�6p��x��4��q�t��՜k{�񻥳�7�a�'�b�-\Â�@%\[r�k���w>��J�����V8*�WNB�<���kBa<6�)�-����0kj�p�ٱ�U�y�|�;'����"�0�X�5��N�1:b��s�x�t�|�جh$����w�o��ϛ��Q��0\ڹ�N"[V��IA��ÉQ+3V�-����][�wz��P.���͜�.�r��o�;���.፱<�U��UB̢��H
y�aT!AaFPD�(*���P�!I���Q�XHAD)��Ua�TDXDB�fHL��BX��.f$a*eVEDF`Q�QY�Zbe�`F"��+�R���-������9j�-�$�5V�K�k�[�w�����h�/(�W����
J�c��Y����e�0�G8���5�Zzo�]���}呭Y���Ef{�ҕ,^�1�+X������j��F�\�z���.��'�����a���`�T�w2-�}BB��מ���g�R6K��m��Q�=�(k)[�l��^u�L�R�gY��K+����=�����ߣ|����xP�B7� �Ң�&�-w1ENl	Şgm�O�_�`f��w���{9�Csa��=�
�G��#��\�o��_��hN�n=v}��{��A���`��"g��f�"�1�F���u'�\K�,V'q�Q�6�5�K�-�4ݭ��w�bo<U!�m�7�ƺ��x��/�J��+��K:de�Gj��:R3�����r��r�4O�<��l�pнS(�����E͓�5A���;ۊ�{���:�N�.~2:D��w�ɷ"�-f�f\���Y���řD)��`�xp�9�zg7�/�e���1�!譾�jf<S3����w>�e?]dU9z,�DЙ�j,�D�p'Y���ݎX�+Ѓ�s~� P�ˉ�j|K�]	[�%�����2U%}�(���k��r����kt����DMZ)){�1$������{\�L4��0���{-?n��b���t�����)���} �L�Z�ȗ����re��ʯaf��J�o���0�m�e���GT6Apau��FYG�㾺=�,�:���%��T�#.��m�Re�z_՞p�3?*�U��,�C��Yu����*C`�[�K$KLn��6�x۸.:aQGzJ�JWv�dQi��Z�k^j����0	�Vjj�i.��*�j�M�7�iV��0���koS�0��|x�[�s=�	�lQ�����CN*O23U_��@��[��])`���ᢻ�P����v��Y �ѯ����,�����ٜ�����>��S{Y!�*zINf��5ַ�n���(��3����-�,�w�3�J9$�8d����CitL�[.�k�U	�JL;fاoM���lm��\fL���eA �dk���u=5�zJV�Y&�V�v�S���i
N���pa����bM`7ע��i��c8�O�{�����n�o���t��Z�C���(/g�tB]|����L`a���<���]���^3�>��O��V����a��U#w�t�z�T�oW���:��3����=pN�!@�����B(ӧ2�2�~>����.;�HqI�t�W�R�sy�س�;�ؾ7�f�ZJ���fde�3������0mvJpk\[�DQZ�m�h#�v����_6��^B[�/�����>�}Wy�A�u���ak�K�ẕ���<%��p�\/��4o��q�炕�\��[~�f���ռ�@�j�"�����a�i�;������3{��^e<��K����GS]���X��F������)ʃ�7��d���Iw��r�Y^���ȴ{�A{�gzd��>1e�p�V|&U��癟w��J}w�+h�Eʋ��E����)JN�.���
k��	y��r~^���Z�`�l��{[+]�J�����"�(ξ�cb�.?$z�gd�6N�r̘Ci˞�mָ�9��W��foV�$���� t�1��{� %oG�����S��`���?�)8�����va��S��	��;3P�I�v'r�,/ma����Q�2��T�=���İӶ�󵏠��O�JDI}z�Nq�ڎ���������uXj�3{�4��L؎��3����!��������Y��R&��O:�h\���Rq��5da��E�A�
ը��[]�G%�p.1����RW]��o\���R�`i��d��I�YPܮu�ja�;Gq {�-�.�ٽ�[n�kjz�2_=��7�]#b[��RK+�D��G{3]��r�ۙ�S�6���+��Kkv�@�K���1�c�}*p�Wp�ժ@r�������2�p_7�*�b.�ks��wx:��Z�[�Py�!/Aμ���(ޖ�\z�v���t��wh0hrwy��5��W��Q�w^�/�(U��"�V)�o�wiO9���V;�:�fJŦ�Z�R�麙x���65G��6�݃�Z4�2*'B	�Ijk�u�%�cMc�V^f�5WK��TWI�v1�\s����F�,g�+��\0G�O<������;R�CFj�ZB�y�i����8������7 wG@�3�ap��	�+zӦ��X���ͨ��!-a}ۃjRJ�=��iwU��+y��إ������rձ���p7\����ml�f��gwT�/��t쯒�"�� ��;��q�1�aʰH�L�%L�(LȊ�"�����2B��#S��Ȩ����*0S�������s2@�RIITXU�E|U��ؙ�[���������6Q俟^���β����u������v��5i��M'6�țc�d��U8�U4'3'�<ae��7�!�>��tw���Y���s���༤ƃ�NQ��h��=<�r����}�X��˧���2aԠ<�I뚽�����-�`#hi���2�9������ :���|;z�<ɞhט\+�v��\�KG�#���ڲ�����ф���+qv�p�4��������k̊+��c�v��0 �߂��\�A��+�la�F�ڙۣ��Q��K���[�sջ�v'qXX��i����y�?y�ن��e���6���Y�tj�K�͉���j���z�c�㨨Юn(ڸ�� �P��c����!@M�֚n�s���+[���P]O��������V����1sԮp������b�]�	��w�����,��+kn��*>F�	����'�h��#;����O�{r�e�9�~햜�<���Q��Tߘ�\�pV�&��L��2з;�O�m�/@y�g��|�֭�&V����L��vືS�)�x����M!�T*��%t$�I��}�s�~��:|xn	^���u�%�mу!j�Z���=;
k�����Q����8gi�I�Y&�%U䥃���#��a�=� ��r��U�uj���]J�&�=h`�f��1 ��$'���O���6�:��Z���v�hc��[�R��W!�eV�E�%,4��$�;��í�zME��TF2��)��v�`[k���t��Ti��u}�>֪��W�ҧ��".E"����A���Kk�p�H�q��r*�6��O���,sZ��/m��X)�I�)�g��/�:��8Ny���3A���Ή�ūD��dּz3��^�I�V�t�v�s_[�8 67�{��0��O2�֠�Y�y�U� 7yG��3���ڇ��f�V�*�G�Z�"�ߦkR9�ך]������]1�l��j�fg�on��XE�!	�K����=����`y�!���[��5Ŷ,4�F�*�ux���ea��S�;����
���/��y�7(^��dG['1L�e,K�c��ޓ���_S��<Mc��^�<E�ۂR�=jPu�r�� \�d�
�km��Z)-��߾�9��h��~B��ٕu�t@��J�tݞ��ezfHir�����ӥ��p��*���9$}�}1Vv�>��s�x��{T�K�U1��C�]|��6�ޅifeED���ng"��E�/�;��{�kN.�	>�\Sڜb|�`(�"�ַ�J�i�۔����r��c��а����
����dr���S�`v����ڰ�K����v\Aw߱�JS�^�v��W|L⼘�$S)�kT���LL�H���u�;)a���օ�!fZ�"�:�b��U��m�+T]�Wf�M޻��P�B�mV�gyU�Y�;��ٽm�
.B�p9��"혂�*�:A�H�u�*hR�ޓM��1I19�1~��ӎ�UL�<ګ�V�mWa���ڇh���V	��n���.W�ȼ�s�㔚B���Abѥ�:����#�=��7N�N�;یl�*oB���yrT#�R� �@v�#�8�Hk��Q�d��1;%P�9mӌ��&P5j� �=�7�|B�}�w&,b�v�Y}�P�����LB���m��&H����x��M�4��$*�G�>]���C�|��bʒ���_��fRA�U�;�oBϦBS��=X�$Ds�է����n�	Ռ��t����x]y �֦h�=xC^<S||fX��%I��.;���i��SF�y-y�o#�,j�7��o�[�R��٩9��������kh]M�U?�T>_���y)��=;��)����2�^�\zgBk�׺zfpJ&	K74��=P��qU�q�b�g^V֓�.�s���	����k;����H��&���pΣu׼��.�p�M�\����Rƺ�kK(I���f��\�(8��܎���P�B�@��Ob;ݦ���sVb�W�x.�o����:ջ��@e��:��pG6	��U�D�jor���b���dvnޤOm��Uk�����i\��pa�e�f�%wU��c*T��.˫��:ȅ��K�+"��|2�ǗYm�y��٧zsޅe����n������fr�� gˍ�j���"�˟<�HR[N�N�*�4�9�i��I�˟(]���T7�H�*��[x�#Q=���[Q�#�}� �Pԅ�a=�t��k�97"��r"��;Ra�'54�J��M�N`�U�����v*�J������]e�ث�
3+���bU�b� URF �XX	b�X0�J����D, �
A�PR?붧���S;�����Q�>�zD���Vҏ��&Ү�S��K����'�˗3������Z��/źS.�_�kK��l��h�=�\���[[i�G�����E����h�0�C��lh�]z�"����Y=\];�wS��xFNq}x0)�վ��EGi1��1\+^N�S}@VD�^��6��(3�󻉛���f+&�o�P�9Z�{^��������x���f�]�_e��j����9PL�0vЃ�Ff��J���Z;�Y飶��O�ĵ�"o�m{����+�߳�_gX.�IJ��ojv��F�{sMXr��Q�iN�Wm����W��9�p������Uw&��*�5����|�g���6p�};#o��R�v�i��E��Ѷg]>�8��j��ݵ����h�ق��F����F4`���ͺ�v��3���Z�92�����M椐Œ�����'�����'��Y~	w�,p|�}��of0�Ky��9$-
���qL$��n��n�^j|�G������W���)@2�Ľ��,��.�G����U��Jc�B�kVnřc5�ʈ9Ѵ�>��d�:�嫦_-����_���A�9}�p�=q(�s�����B!NL�K� O���H�8�r��+5�k4@p]�뚱zz���u�@���$�g���^�7 �wRڽ��\���Ùl\O4չ^��:y���<�P�/ ��xx �nF�3�컘�E��n�V�++z��-�ޣɩ�J=��>p�y��8��|�\t{�z�s]�/�4ݢe�<F�k]'˦M~����Z�)���k	-mbC6͢��37���W4C�j�^
Ӟ�W������|��t��8��P��
��v1�uL��ް��c��=�7W�x�;�>K�ć�Xv��[\vQ�R�S��[�h�cO'y̿���_=n�<����ձ�`e���[F$����=J���^��y�V����w�����j��]w���±�,�o�u�#�zq�����y��	����JK�E w�t�S�#�3���ck�,����ͧ��/���x���5a�'�Ǉ24.���nm?c��՝հ�����^Gq���c��D�{`�}�w�3M9�;�4�����H�`r�W�9����r����{�}��Q�ˬ�I7v�^�SU\0jR}T�VM��[��2ho5N�qPm�c�֣-	��ǭ�2�9���nU䵚����S���X���^�d��4n�nii������`ns��?#&�WEh�gnV��y���}�"�cG��%w<�-����8rX��3���kj.v�_F�6���s>��J���[z��]��9�*������8��j��["���nk��jrN�8Kwm��**;��g�gx]��^9���>��>��ڋ��v��/\r��}�)[�iY�z'B��H�ÄW쇽pnT�����h�u���H�����4��ò�ܼ�:��=b8�2��*�q�l�Z�8�Iim�+W��u�+j��>[[�N�����P�=��Vx:U}�=3�#��ݴe)��_9V�.�*3\ �+UB�T6�	�`%�n�5:J�+�`l�&��31S�r����b���:7R|�	������$o7��{^�̱���wK�|t$����Zo:�]���(}��:������%�=�r�dt�q(��un��	�}�1!%��k��t�_U^{����f˩��ʖv~�f/Ɉ(ž�{�&{I_`q'������K@���'DX��N�)�ٗ΂5��U�r�e���/������L\����y�qY�Y�M���l'��,��� W�g��xj�瓗Xq
{�4���b�{ѧ�i�7+H�|s��C1]�Jܑ\sZY��j��׏��Çc G�q�[��Q����u�q
�G�L�'�n�R�LO&�ǽ��?��q�6/�ݹዛ�,�e�e�y
��ce
}Z^�㘂�JZ�k{�ˠ�R�Zw�	�y���o\al�{[ΧrV�J)a�����ɘ��)Z��K���om�*�:;�w��xF+�Q��i��*���׸Fn��ә�����e�U��$ʾ�K��ڐ*�\��OM�`��
Ր^M�T�i�ʾ�v��YV;N��Ȇέ�fi+�=�n����{���X������0QXV\�2�֌ga΢���E�JjLҋ�iۗK�4_��$�0V��y�;��ƣ�ܔ���^���qpq%Ľ����h'z쮈Z]� �;��a�nV r�2-�j��i���H��oU����Z6�*�(JT�*��s�
U�Çh�x���%G������;�GvV�V�PW@��]�w4쌎�iN�2��l�/7yɛZ֮�^Ke � X�"RFb% UPXj`�HX� �	HX�!@�bX�$@PPX��	b�H�` SS)�,A*�,@̩
J�D�,*�B��H��(���owz�ާ���n���}|��'��1/o��&5|�b���)>q� eo�~�#S�u���0!�u{� ���a/w���n��<&��9X����7�B�WL�,��*��v.���]n\�����͍�H�;��%L��?6M�ug�+��v(*G�HK(Vݍ�����՛.��1X�E7z1k-K�y*vh�mvr����Σ�b���56%Ws��HLY�3�c?F������*	�/�c��K�⚳���`�k�yqP�;�T+!�Zǥ�R[�}�C�� ��t�8��G�B��,�Șd�7:���:z�n�bY�@�ujuuj^�k����t(\�&��s��2Ԗ�ԫ����cT���{�ɽ7�]I�9݃�XM�틹�������J��G��s���_�r�mD���<���h���˱޹��B�<�ћ�{G���<9|���q)g�2Z�R�a�zT �8�ǻNF�ڰ��,u,�8��-�Ҧ~�⫭���K�Ը�P0��Ǜ��EŐ͋&i�{=��s�����d�Nt��vc+�369ĝ���y�mR�hv.sj#of�R8(�8b��OE+�D}`������F�]�7a!�V��g��3SB�p=�DHI�qIYz�m�������8z�u�wN�6 �ވ"���q1X'[�9���z�hjɷ�MT�i�%���h�7��1R��L s�n��[�b�GTm���D���C~s]�(��m;&��}��Hl�ڴvьgM�=����%ub���v��J(r�y���(@����{1�C�Oom�
�MLEoE�%7-��WCv�������H�ih��f�a�G5���\��cKU�ݡ��g�8������g��n^I��_����v�<�#��������JF��t��*eY�'��fk܀v�\Y��}��A��%
��6�@�J)��o�eP��os��	5�jW|{�T!M������`�����~?F�J��j��w ��	c�Vz��8=t{|n���e }$zon���0	�>�sS��U�r���yj���j��s �e��5`Mw1 �FDm��*o�^H����uu�z'7X��i7j;��{�)F`�̊��mڃ;�Eh���s�~3�ue�^JB��n:E�f$����@{�K��:X8�Y��;O�VHZ(����
��$.4L����_1DJ�L�Z�c����<�V�:y�;Z��Ӥ�}�i��W��-b����"v]��sN����7K��� GY�go��Ѳ>G2�I�^E��9x��:�n��ǥd�2���Al�.����W4D��[G�������nh��*A��Ǐv9.���|�Oq�6��s�\)o{V�����OXu��[]]�������F�8��1�D9�)K���h�<�L�͚�K��1��3��38G12�}�J��<��;�^I��o�Qpmگ�P�W{��}R� �c�����RFt�(��B�m�Tȱ����ZLhJ�Cc>��3ٶ��H��S05܅��qӄE^�"���q��_Zf��6�f���f�k���; X��a>bO����������X�8!b
��K�h����i��O&U���2�d�/J/vc���f�F`�~������E�w�Yy�=�)���nX�3D�e���k41k���O,xW"�i����g�`->b����q������ ����]�
��%w�ү��}*4��r�5>�N{��<���������'�h��l��2P�ݯ��w}��r�B/J�g)j+���B��VfwZf�����=4��(�S�!L��^��ˣw�'�^���e:���UIO�ߵ�p�w;���ɝ�s�m&S�����{7�_����&S���L`��\'J��3���%�.��4����jM�$�Y΍���%��i<�x�w�i֦%����v���b�,��ۗM�t��FS]�9�|ޫ2��I�/�)�I=�#g�Z��뽋XB�ư`��^G�T���h,v�/h���ExEG�oɶ#K75a���uK����᪂�fJV����?�-�]��P����r�n�v�Օ�4���I��%>�G���[vq����R��ݱ�e�K�Ju�bX�.XL�%�H�"<��/���~�`ث6T���
}Hc(vZ���f`����m?������_;U�s�n�����B���ij��·s�Z����amv���tg����*�%��.��[�GV�E^�����IM9w�,ؗ�di���j��[2�tL��T4���n\��{CCU��K����^D��n�� �M}#@!`�������n�+Q��,��Ȣ��k�'�F���2$M� �n|2�A=�P�t������֪5W����Mq��|ѷ�nYB��;�cF݃�r_oL��M�'72�φ՜6���KjP�Sb�΂*
b����m`8 9��֊ǆ��о�l�k
]+�6%��#`f)fV�]��K{.i(�J�Eڐ�t�g���?}��K,�
@��X����AHb�b� RP�`R"P�DD�F �0"�,SI� 0�b ��1�R�|�]���Dd�Y"a����1�N����[mw��߃S�\5��^���������yt;Y�y'S<Lߨ,c�+}�mza��sss�Q��zJ����5����׎ٺ:��Q�i5 ��i��9����ŏ�Y�·�^�U
	~ٍ�����Zha�;ګ�g@QSY٫�{�xAHo�Ѹ���d��.�l{%��Q��͹L&=%%]Ѫ5\Ko��R�k��ÿsi�ILi��N�c<���'^��٫u;0$bf<�^��ٮ��4/�?~?����g�L�n�`������Y���F�P5:�{j�vM�I�G������_��Ջ�?�6�X+��f���ݑ�d���^Â�V0R55�و}�P����1{���0���kw�_9���Ii)�G��d'3i�N���q������ɤ�	��k>~�?��Y�������W�J��b�b����g��A��� ��B��}1�gmu�;>�=f9%:k�u��
�}��b�
��d���~�{\�==���V�ɖ�o�f亙B�皧la�^�<M��oӖ�G&�ē�m=�w���};�ھ����c�I���^���Qӛ���r�{azsY��˱�Z�� Oޝ��3lg�g��s��=��D�]|���
C�B��Aw���w\���6�S1�S�'N{��{'
윻�U�G�b�**ݯY�p�?n��h����&��8E1��P��7.�:��f	��J�?cp�b����s���V�¼8!b
��Z*
7;�����ji�)�%����a�^kS���\ݾܗ���衧u%�''-%9Ok^��2��mz��μ�?A�r��0A���������٨��S������X:�}ۅ�����7f�\7b��Q*X�<�4�u}%����s���X�{=F]�I��=�c.�1=���x��ާsʴ�W����(�3��dIL���Gs��2؊��^�{3m1�PێI옣Z��K���~��g;���wܼ�4��{%�Rq���������n�QlS����3Ub��-<�7"�ǂ'�à
�1�k>絊�c���lK��ݪu���s���:�n_z5�"$���f"��ɍ������--�2�m$��n�Q�b� /�M�g朓��QH����aW��;9�Q�dvB�-�"�v�Si�[6���-�?���~���+��0�C�f�٨��yx����N^h%���d��f%�
y���K:���u�T޺s(�㿈B
����#TEL�񬆬{ƞ���6��������d̒f��W��K�vc�C��󺦦�ə�*`���<MvOvu��������r�ft�;1�8���f7E�$!<�U�ܗ�(��۠��;��vw^��V�k���o[䖖����wyos��{�N���S�-�z�Qn+J�׸z�y5�j��8��.�f6�;�KV�36���\�tt$�9}�y�4�š��}�w[�\0~��Ex�g No�n����=;����s6�i=�8iǤ�j���%MM�m�{����wRSƤ˚����g�r��E�8����PB��Z5�}ٞ�|<ҭ�
�N��0�L�i�M꧕f;�om'[=�2������M�b}zs[��~�����N0���?��!aҭ�r�Ш<��8�Rg�e��k3���em�u��x��T�%��0s5n/��Gf,�ߝ�sUbm2�-�R&d�LgN\s�$�X���l�kp~�R��w�]6�&E�d��+��<�w#h�ˁz8X�ؾ�i3c��}h[��'�#��UėMrM�t�S|�Jo�r圚O'1<Onp����o�&�F�/����2�:t�7z�F7ɷ	�S�=�����G��d��hG��w<}[�e��n�źe�$�Ų'kti��w��N�j|�|�S�)���SΧ[�yʺ���%���c�"��u����U�l�x���>��9���&^�����)��x���P�X�N�������2�F?e�a��;)�:�J��l�}w,�}]k��pN�]�c7`�s$�/�yt?e,�
#8�+��md]c#�������t�ܒjVJ�ɖoYw���qل��t�lǧ��fN������㭧��m���nq1�ə(߷\���i�u:|�u�=�0��e�����n���6�tE�1~��x9�b��۩mۣ�s��[3M�K����Ġ�7�{/�k���P��P�ii�M�{ܛ��u�/����(������'Oz;<}���I}�q��d��.�`��N��烓�η<�巕��Y�[��췻�a%�>c|��> �!u�e���u������߭�:�=�W�s�h���n�:�o[<ƹ'q8v&3�:�ڦ�<c}ɍ��|%֤�o�)�=�&^L��4������؜JcؚN&_4��r�on�S»��S�{٢�4���]46���~�/���֊b�
��GMz~w�;�d��5�:a�x���F��b���4S�%3�-�7�0�d��s��w����r�<����I��V$��~����}�l�-9KV
Ē\���9rg0�{�Ңъ;D�V$�0�nE��<�n��N/{�9�L��.����Vt��t��ki�˗(e�$��u��3>��u��)~5�_n��Q�Vj�~�������AMN�K�HFLFO��;2��G��q%����9%�Ճw�z��p�^�=4P�
�N��tU��
��o�z�*~y�Y��԰���4�Վ�o2���}�X�I싖�x�'-�c}�}x�r��nOvOP�*hN���|�z����Ww��-=wڠ�O�Ô��ǻ��\�:�ou�I�ɯLcrO�\M&ܲ�#���{ի���7���o�an?���w�!�um��)�."�5�uZ\�⻢8!�T�v�i��Ã/bӁt�'�)'0!ef>��.xU&F����4@
�&��5�D�S�#���n���ڑ��d='	Σ�"��ZM����y*]����ö��+*7%�N��aK^�ֶ]��#2YT�;1 �|�Q���`���.��<�ȏuÁ�aU��Y�Q�v��ѝ���ݺ��Փ��;t�ʝ"|J��)�l����ӞB,.��o`!���̍ʺsj])&�		�5�I��EЕ�CM���݀���|���[��xW3]�S$kksV��˲Ah�E��Vt���r8)����+7=ߘ9W�ebYs)�]fU����J�$�RK��*�����y�H�W��#���C5_�$��δ;b��`�i*�.l���ѭ��Y������r�� S�tvd]ӹ�& >d*uIټ�˫�&�qI�Ri̑��1
�P�� S���`���0E # (� ��R%X�"X �0Ĥ�EH%$��)0��K�) P�"�����$ ��$B1u_}�'6��y�^Ϸ3�.� :F��n��N��_9p�L2�&4�̙�ž�`��\'���U�"����|T*���;~�����u29v��4�.1���+�O�6��T~_t*}��DT�Y��|�Evp���W:cx���9��5�n�o'ݼ���OfJz׻G���&6��7�<V�F؁1銡��K�0g�6c����ભj��Чo�:��h��[x����L��:*���a���;�@�޽�+M��v��5��	avĸI��dK�;ۗ��@ʠ�_�'K� N�+�}�)���X���I�v.d���`�ċ�i�d뷍������*<�'E8����x�D��Q\�.�1��H�\9z�*����CSU8�Ǝy����h�-<'3�VtJq�O�x�ϵF��v��n��z�7)�La�ItI��۴�N�LdX3f��Ut�`q�"G�k�����خ��U��=ә�a~?zp^�����|�&��˿l	����NN���r����1X������=X+�TT�b�+ƿ���d87ҳ��«�X�E?����	��'kFo�g��2�R˙��!_6���j4�
�o����(�λ�9���w8UBx�γ�5xb���Λ���wM��AL �U�� ��][4��9�mی�sV�OF�T{���I��D���M�b�Fd^��b0�J#��>~��ګEV��l�9o�^��&�Id߰c�o�\�Է(�L�%,���C��dG0�2�΁�tt���5���͛}s�lk�SN��yFnm�<4L�Ʈ����ࡦ0c�FΓK�P�nt��B�
���V*��8���\s��1\8jWޝ!�z��4���,W�TV��6�b���u����>�~"�M��d~�c�U�a�����V6T�l�*r]�.-}�7�|t��M����))�����ޝ��IĤ������1��ϹY{��'��nS�_\�O!�\��s�I��Y:�5�<�W8S��LPV���.����>VN=�yrOs^L�c.P�e��-kI��I��'?
�����5S�Y��1���"-u���ni&�ʚ�0�����}�|zor�-\�6�n}G�<ܜo�t���1��z�{3!O�v�us�ɇ����A���}T�A�_��LR��n�ͤ�]z~�ߝ���e̤�v��<�*Չu<M��\�'&�at1E+{�l<��T�I�P�b�ٸ��v&v���D?q�ET��"�!v�s�\����{=��q��u4�쒓8;{otFk���#�X�W����o�׃o�6jT����;F2cwL	��ѳ/���`s��p�Q��������/�����<������Kz��=cf�!���곽6*�k�=&o��v� #$s�"�m��]���6}��
G�=1�>���ƣN�����T�H�s��dԘ�;?�8˿>ny��`��٘�C��ʸx`���/��ID��{h�Xn�SV������,ZE�f��/����P�i��/Əb��[��G��1���2�P���1b~:.(F�1h\�K��5}��ȩ������bӕ�*�:�]c!�;��[�U�����D����)#Po��4?�)s�!0f.�����ݡ1�����n�rWc��#����{}Ʒξ~X>ȋ�����؄tL������\+���1c���������p����Jr�y4�۷��ԕU��s�����m=�<��X���k3�8�W���}Ok�t	���%K׊3�R�㴕��fr2x̺`����ɪ+�;���V�&*�Vz��A��H��>����p2�S�>>�#����Ѽ���c�G�[���U�� �����B���ZU��Hׄ�
�7"��U?^��Gl1X4X�����5wj��\�?MW��\�UF~��:u����|s����Z}�5��W'�mö:��c�u��W�W\1�מ�Yu��s��b#���>t���4^1<#!3�.��Kr��	�{����hO �FX�8K����b#2�lסc�W��z��f=�)�bk7F�m���=��9@��Ĉ�Ƹ�<U��ם�{�-��9�=��������Ѧ�t׬�4�i��u��;�R)i�N�I�����w�κ�8L��>�ԙ��/�����>���|蘨+{Pӓs;��/k��;O�x��rsK����n��u�s:��$��kEFjx��Y���^�]������c�F��U`��,�ǣ���x]�~���8J4�P�L�g{��s��:}�����c|�ZkriӤ��i+n���F1<M��1��&P�Ry|�U�GJ��ʼ�k�jM��{��ܕ}��j��ʇ4�h�l契YJ�9n�ۙ�d����^=�F�r��mbv��v��ҧϽ�ӉZ=f�{e�u��\6��놌>���%���9��0�穜O��zwZ�o}u��M��II��	\�&��w��1\�k3��&v�0=IL�q&�4����|�\�T�.�.���8�E�)霵3�͵�����h�8f$B�h՝��(������C�`���`�4�]�0״�ʫvz���>�E`�?*�@a��r�c8�k}k��{�q����i��Ytg��?�k?�#Ly�P��So]�K\�vb��N��2���v����(Qyïq欥�w�� Q����<4��~2Ds�8��t�Ob?\�����_T���)Ɏ5�����G�H�vv}9/����1z"*�4}�\�f!�Oؙ��^'��\����:��r�O"%�L���/����L4�����n}�|9E�˴,|����kg�a��3ӻ��!�O{\L'iO���×�4v�޼��^0�l�AαGH��`UeNnfH��n�:v�꼖����M!�ӎ�k��G���,R��ʗ�����GƁ[��`�����\1՘6��3�W��6�R�w�\p�3�ÓW�0��5w�"����#�v������{��m(��5�,�A���;��'s� �s�;��'0�8�J��rI-��b�z��wmt����Rm�k{��(��7�=N���5�+��kl<��M�S�nF�:D��{HN6>b�h��[,��Y��k1�q�.7�Vq �.�9�v�|�t�kw���K���;�{���u^�R��Mn��^�&9�v�g?]%)ԕ�Z(��o��8����}��AhF45�;6J�)AR��턪[i� T�&FW�ΰ���ɠ�݋�p�N	�U�5�'.�v���S�a�3T��J=�����(�U��㪥[*]�+p����`�JI���(����^bG�S��P�z1�h+�h*�˥��&���[6�7�^�JF����Z�u*|L�%��u4Tc�mq�eV��H䆊�w(>�6�Z܅N�ܥD��/'B%b�f�w����u��/��B$T"P�#IR)��AH��je����I�"X&��B�$DJ�R(�a��# �HaP�	3-`fbJ@�XD�Ref
���"��	���f��y'vd��![W��_�~A,g�H!�����ߵ�3S�j0��j��
��ɝ"2cg΋0D��[����_�=1������\܂!.vj\��l�l����"c�DI쯌X2g,�90����X�V���]x��	�a��5���o��N�L�x�roW�mӧg��u�_\����$SLԞr�ƦӮ�#�H��y�Ez�����FL9�ɯ��j���<<�����f�X� ~5P��,{M����`�&��s�Oߕf������>�'e}���[j�2���/�V7=��>�Uw�ǅ�'���.�<N�*^Vr�L~�����l1���
W��5-�鑛���ܡ��
��4�td��~N����f>j�:+¥������#VWx���!"��u�e��$�P��e�.�3gQh��$S���]�Xz6�2�B��|��`��o��>����+K�Y�l�v��,%a����ޫ�)z�N�f�Y+���� }O�l�%��C.��)���:\ڥK�	~�� �2/G����s�⭈�p��*����Q\ߴ��74�5�*��u����쭐6����+siK=9�}n�X�u��2鴗Uc��u�4���aܺK\b��|��ˋlm��F����0:��cÎ����05�%v�q)�
&7�c��:�	/J�X���?GfF	eg�i����V:l̃��, ��
��J,f�w�	N�����^����i��Rٱr�Jl�g.ѽ��3�;\6(yD�¸���9y�L���[N�k!<���>X����uOP�I1Ӫ�V(a��w܋wK��hu�5��`D���^��[[{���C�qb�I����=��+e�ٝ/q�qJf���{�q����zvcu���s��v�,��@Kn��O�ك��%��c��F��{N�_��u��m�K�[�pkx�痵�V�fuxj��H�m0g�����C�k@0=�J؄P�ʹܻ�t7���G�ЀN�t������׹�p����Z@�PQ�r:�:�:Pˢ�I��nJ[�N�پ��*�n��9���^�/�r��M�dq7��&���M=�9�FwxA�I�r��|�(7�kK���T�T��;kv���Kwhj=��Z��iq�s�~�
��{��q3��t��
J
~�R�q����@['�j��*���z���4�IX��Z�4�Y�!h���k��<��vFN�0��/��YMf�.T�f�р���X�u);�+�v��*^���Mk��{(L���L�Ǹ���4j�m����3k�㠌~}H����
H	1�.M���L�jZ�.׵��_\��;0&�q+N��7k��ܐ�u����>|��:�:��o�'
հ�O����[� �o���ǁҫw]��^�W}���!U�X��R�!ۡ���u��i�G8��Dg��S�	̾�����F���Zmm�%�>ؽ�{��1�m���j��q��V����6Q�D黡��VM�E�71x��4�;�^��)�<�E�;�*��O��J���	n F��᳨\��l�(�ȼ.(�}�5���=q��r��F��v2�¬�N�s=�]{��m���P��aH�]{�e(>������,�Ǆr�u�sI��E}�<�%�|V��6�ٍiՁ+�H������V�(�RX��f�dv;5��*~*�jgwQ�5Fѽ�+��5��@䈫G�+����f�� *���Ɓ�\틶�<���IQ���Z� �tح}9��S��Ym��F��S��1W�SOy��un�s���X�<�H%����\5ה��y=->��.��C�w1G�z���镾}�M���^�����ĤS���'���aЦ^�&���샽%5�!@p�B�սJ]��#���1�(�,��6��&���π��<:�\��J���{���;���ROYvN�+�px�'ɴ���r��,�O����c|��g�>c��?�T�$�UUUU~�&aT@H���誈	�޲�Q<��t�"�����c��>X>�Ft�(:S����v�F�EEV�
�$(��JF�>�I,eE�`�'��HD� b2�й�:�d[*��=WGhT�����h���`J>�+�F�ݭp�7����8_�vF��@�D{���w��d�*������4e]�=!s�(	�袀���(D$������������'�M?�����,̃�I�ઈ	����$A ce��`m� �C%���CY`':�j@$���&ziu -�i�����ȯU�4I_H�Y����" � l�f]M|�#Ʒ �'tHX@��
 `�V �@ID�>i�4Q�}ٍ���.X��LN�T@M!po@���%�</��[!�=�I�A{�˜l�HMơm����4���O/�{���7�L�2 (	n!!�X��C�W��xrM_j*I�Q}�@�$�!�CӦz��/��=E�b�V	�dSJ�e���f5�EQ5&�0��΄���Æ`��~#!���C�@�P��T@O@� �����Q,D���W�$ƫ��$��,���PAP�p�FH`tF�k���`Q�U$"#$���!�>��m�ӱ	��X���#0�B�Kܓ� )29��k��f�~e�3���Q٠j�Q"���OP�5�Z�� }��H�F&���>.�ڟ��;��zM����9����9�8<q�O��`S���J�?�"����'e��#`�޳$�q���G��*�	E��f����e���I�^ZR�v�C ;{�-�f�Q <z�P ���r� ����1��~@� ;�b<{��
`Ϡ+���G+
�_���6�[�Sv�OEK���H5�-���9��L���v�X
�Hy�:q]p,
#e0(�oa�kp���(	���HK�M%�~�B�k1p�0!f�]�)b�dA	ĐN8�@�c����H�
�P��