BZh91AY&SY���( E_�Pyg���g�����   `��  }C (!$�T�J~E<�j��m&G��=CFhOP�<�F@���TFF�A�a �   8i�F#	���12dhh���D�L�#  ��d�bA�T4         �M�4L&�P�=G���)�#!�G�|� �MI �@$� �-K���0 ,G�	)��d9��N}Fs��5�������T$$2���n���4��^ɹ0*կ��<�������x��̼i$�I�I,I'I$�$�����P�JRL�I+I'I�VK���>�[�pA�t4��ȗ/�� ��l���v!Sp���JSD��r�Q�yx��pG����߾?~|��a�BSj4�P��q���`��T��:��\�-�];�mf9@�!!�L3h����3��Ǝ,�0_��#�/�4�.r��Q�ɰ��K��u˽z��}2�)�O��UU̗ʜR=���s��̀9�wx�@9!�����4�~�DH��u T3��ݭC�Q�<�&����g3���]��g2Cz���2q��<�.z��'��}��s]����{W��Ib𶦭4h����CX���p�C�5n�M[$6��݀�ó<s�
��VuY����済��U�`l�$Acp䰳V�"��)���.Q�6d��Sw��w��u�(�H����ODMP��f�|�h���Ko2�6/n�&õ����0�lpjP��L]�mD^�oqWo �h|���2��ف8�y0Lf=�k���];�U,����!IMf�Zw#F�`$E�vy\+4�-N`�]��<ˈ21�;c��*q[H�/K3[��^�QX�n��||Xbbq\��jU��wuWz^���2q̒!�$IkZ*&����(�����{�N�$9s d���c�P!r�\ *�*�Ե  %E 
�_�j�,@*�� Z[�h`�^�*E����1ִf@!�I���;��ښ׿�����Xx*T7K}�;r�b�.Q�l��5�5�I�\3VwE�u�Y���l��X���=Su��w �	Fi��4-��D#�9!#�p��F�#�����<5(:e��J#�c��Bù!#���+�1A��� �j��DB�E��y��wQ�J�l���W*D�~,���}��r��� -BL�)�����nG����k84І�� ��򛂥:�>qj�6����^�������ѓ?"j�0i	R\9#�WM|��dɝ�؆&�ن�Y���P����f�B��t��bBD�m�����G��Y\V��s$
�$$x��h�9{��0��kEKfdi,�!H���+J�T�(�1 LL$���I�AK&@��H^�Vu�E��CU-(��
ayǻ�C�e�	dº�$��4-F	'
��H����<���z�@��S˷jBE��2�%r��l,��;�I�9��&]�K4�����h�*Գ]��BEn04�*������5%�3��q�m�wU�>��H4�f��$gḀ���e��sj���@�d�`d�Q�,?��H�
_� 