BZh91AY&SY<줜�ߔ`p���#ߠ����   bF^�|            |z�d�j�Y[m�,m�ԳKT��l�ĶU��eEj���l)[mP��V���ZVڶڕ�mMJ���mDڵ3M��cj̕��[u'eY��mGv��h�kZ�i�[&�*��Ii�D�[Mm�ڶƖj��Y[mj�Z�v�V�ji�Z-�kY�[m�`�nvwN��,v�   ��/}{�*��ԟ�ice�hV�r��;�S���T�n�N��6�W��Z�QR����m�lm�v�65��n��Y���v�f�L�P�km�����ta��-��s���U�}���������ά7UMָn[�;n��K�̻i��hWq`�v[s�J��wݎk� ۻt��Ti���mV6�����ֲ6[m^�U)T���J��nZ��U"nso��J�\��D
�ޟ{^�/l�']����������J�'��x� �������E(�ZO��P�`
���l���Xe2�[Z4�s�*U*�����ԥ*% }��� 
�*9�\��@>�����u��T����}���P
�E���P���W�z�U*��x��㪣���h꯾{�_M
)N��zU�
U�/���U4��3l6,��y�J*�������J�1w��@Om�}�ޥ*R�='��:�٪G�>w��J+{m缪�	���=z=B�nw�o	HT�k��kׯ%�"��ƺ������Y�I��ѳ�o�IP����:��i���zТ�m��x5EH�=��B�m-BT�9��*�m�E�7P�R�`۬:�;�[{�%U(*�{nhQT*�.�R��R�2T�&�J7�UUJ���4j�i����@��Ҩ*�G{\k�T�;u:B�(����T%��p�t4z�h �X@]v�  ��im2f����["���g�UT�N�� �=� �[��4�:� �p�p ��p �ڸ û��݀�F  ����4[fj�Vb����+UN��  >�^�(�4^�@{������  �W�� �^�O �� ��N� :�  <s͡��5n��i�b�o�UTUF�� ��@P�t -� m��� :<��/:�����]�������� 4{[ikMfm��ە\�Ufd_yUUR��{� 7r� ]ٛ���'  vR� ,L �ZE v�  '}
 y��t4��       ��S �JJ���h 4A��i�����      OC&��I  �     j��@��*�       ���
"b'����4ɠ�@� ��*�*h=L���� d��7������^>��7^{;�
��޿]�߾�����-�:T��
�u������y�<��� 
� EPT�P_O�}�*������/��W�_o�~����_��A}**�������D ~$�eQ���� �� S���ab?�(��TxX�Y#$�P��#��0��T�,FI0�����)TL,&DҠ��ab:,�����T�)&D��Y#��aD�I0��ad�,���2�D�׳�F�#J,#J��,���4��Q<*&�Dad�F�,&L(�Q=*I�!��0�T�*FL/�H¤�,,��!�"ad�)&I0�aR0�Q0�Q=.�"tX�$aD¤e��ab0��R\(��X�,FL*&H��=,0��T������aQ0��X�H��|S$p��XL*&!���TL*�0�Q:*F
I�A����T�)>,0��(�XQY#
��	�CⰢp�),&H�#	��0�*)dI�$¤aD��Y#$ad�
�
&#
��#
��H¢0�0�����0�XL,��D��0�QJX�,���0�aP�Q&�aQ8T�*FL,F$��0��R|TaR8Y#
��
I��aR0�Q0�*%,&HaD¤�����aRRFH��aD��X>)��I0��R0��T�,&
��$©IXL,��	��0�T�	�H��(�TRGe$¤ad�,��ʌ(�Y
#$xY#"aQ0�abvR0�H��L*&O
�����pÐ�Pad���#≅���p�*,#"ad0�F��aD
���¢ad�(>*I�JRC
C��L,$��O&�¢0�C��0�&�D��adL,I�H�I��,C$�TL,I�!��0�'
��D¤�Y#$ad�X�	�d�)&#
���������XO
��H��:,ad�$aa0��"ad��C��F�,���'
I��Y
�aa0��T�,���¢�0�XL,���0�Y#
�0���HR�&�
;*FaI&��I�R�¢L*I��aA�A�"0��(���0���0�ac�L*aL,°�)�XZVaf�0�,��)��0�,°�,°�,��+
��<8S��aXVa|+
°����,°�˅�S0�°�
�+0�,�ϊ��,�p���0��L)��afaf�p�0�+°�0�+
��/����af�aXS
Y�0��
°�0�K��Y��+
��0����S
�Y�af��Y�tY�aL,af�XVa]�aXY�aXV�0�ZY��Y0�aS
�
af�,°���Y0���0���0�,°�,��)��p�0�+0�
|Y��^
°�0�
��
��V�0���VJ��,��,��,°�ZY�0�L,�
0�
ag�aip�0�,��+
aL,��Y0���,��)���8SS�f0�zY��xQ<*'��0��,��H��X�)��{��?�N�����xz��`���?�HK���	ʗ	E��WR�鰕ڼ�����fm+�	D��co7[v�U��_��7Y��s��b{^l3�ˀ��UD�����*�0��[W��Ղ
!3G1ki]�Q݊M��U�mV&ئi��&�$"x�\cCk^�5x6
���s̗j��Z����3OQ����t�OR7�k�Io.յn�/%��i͛n�k��vf���y��SE)6�KdĶ���ǘdّ���%��Y���x�yj�:�֦eVD]�8q�u�Il��y�d�g2Pn���5 ӑ!�H��n+�R�mL�9i�@�gl�#l�%_���\�^�r�$m:���Xq-�J�c��!k�m<3*�ܪg&U܉s+#�+r�Y�����BX�21c1Gr�V�U��V��'/)f��,�?V^�L(\��ӨuԨ�i�n�::&lV��IU��������ڿne��Ii�J�		��ͣ�s"1��r�%"v�UXKB1,OU��vw/F^�|��M[L6Ff�v�%����6�-�)1�Y�+I�Vӹ����U�5��۳�pv�2�~j8Z�oN��⎭�=��fM� 4��E<uB�T�� �;nӇP��)��`��G2�V4��U6�ӳ�uq巘��c
:�"eR[w��S2�-E,;r���̫����D����+U�Utc%S:��)��.�ś�"�uxE�h�s]���nH f�y�VK�U�[A���2*���
��7/���w���^�!k�l7��k,�ֆa�WZs\�>�2�r�Ƃ9oR1�T/n̫U"r�y%�$F\�ۣ��eKR�d�%r�K+Z�#�k:w!�O�F!/Q	{�����n�[mf���^�FeD��nZ��8��3$���V�ed�0a6ُ�,-�"�U��%�8�+���&\���e��x�b޽&�HjB�ZjAZ���Xr��F$k6���	�bv���tv���˱D�kF�Cݮ��M��T0�"Ty��/(M8��&{B2��GQ��M۱�h2\swos$Ow%�WF�)6f"&'��0i����V:7��	l�1��-�,ʹ�x�4ʱmt�"�*Fk�r߮��2�15�!��eT8r��5�-H�8�D�1Uf�Cetն�ܢ��b҅���Hݜ�X�(nm�sb�UGa{��ީ%��+.�9s7Pp�݃���ی�Ȭ<�R�L�r��"���v��kZ�f��Q�+n���K%cy[�5��޳u�z��46��ln��(AY�F���d?9qͳnbz��K'��yb�ݦa�xC�-X��VJYHkXʸ�Q��-P���k.��jkq[�;tu�f;[L7E7��ӭ'�іr��w�"W�w�p�s[h�%���R�c�d3*��y�T%aҡ۔i��BRǭ[�UBoQgo.��;,��Gj�	��j��n����iB\�"E�j��u��թ��x���S� -&��B���D�M�/T���(��~U*4v�;�I�cE����(�.\U�U5"��mf9zh�l�A;a�ɥ^��`�)�71j�f�;5��4�ʣ�n�Ҋʼ9l=kp�n����.~[!aQa,яq��m�͹���BݱtFDz�N�e;ky�
�-�;{��Xf�{��m4rB���[L$�ωw*1N�+a8�8��%�J\J��?&4���&Y�MYWQZ�����
�m�X���,�ޒ��MnҢ���sm$�Mɖ���Í��sj�v�Si셔����.f�ڋ]d�FE�ˍ9�^S�2���&n2�[�;imcWkؼM�n�d��5�p������VV��Ա/I�^�S�ċ�IwYܐ������I8�D%�:�zޅ���(5��Y�c�B���)�L�ƴ�iʳZ.�=���ZoD���I�n������a{�P��3hۺHq��-~˲.�5�6�T:��V��Z9��xjC��_���6F76H�m�ӂ,�3v����[*-4A-س! �*�;%�97�+S�⤲m�%��˸%�vo/J��f�͓0�Қڻu3N=�)��ʌ<z�m)wtɩ�g(��͖�vYSmR�����仈H!�M�l��e���4s%��NŪ��.;���D���f^
�L���Ov+VGbaӁ�����i��1�nX(�)����Z�EQp��y�GR�HJ���W.����83(�P�Zt�6�7�[���r鴓.½v����=wxl�&b�)5��L��P��J([i��*�~Y����짎
K2n�H�SX��A�-]P��)Xn�*
��Z雯6�SR�i�+.ݘrC��&=�3o%�1���h�컨Fɶ����[7.&]�v�*.��oe�6�`:���,H�QaN�����^��:/rλV�9^&<
�BPl��T�$��7Ql�����l~�bBk2�D�n��l볡.�ٌ����=HE�I���c�[{��F8�U�쥷���!r�Ʊb�0�Um�DR�9���iI��S2�fD7�-f�&�p�6ũ���<�;�Y�yP����˄I��|��t�n���.��V�U�Zv��E���8ј�[8F�{lj�tM��-��p���m�y��qo䐤][�kqj��V�� ��Y:��+)F�yL����"Ym���xq���-���n�M�w�d;tsCj9�
�t%V�f7QHT�:�E@��ɉe�"y,2��L�p�c����[/t��j��y�U�QbsJ�gh�b��)��6�:��v���Sw�^xQ�1�i��l]�B��x�HB���Un�3�S��u�z�Y�����Y����W�v�ӱ$��]K.�Y/)����Sq\�U��(�J<v��t�ePU�������B��Yq�x�[uH�Q̣wna��;Z���7��4����T8UƐ/5��� R�u���gi�n�ۈŲ��n��
��d�˲IC�N�9JP��"�(H��n��!��:����j�2�A˻�e=����n4�5�S��U�؄
A�{j���e����^��ʳ�.��M�W��UUD)�U(]ɯ)��lb���2�٫#�t�ګ�	WJ�+.Z��jf�h��^<@�ܥ��"Rf�zS���ӆv��^5���ۼ�7v���Q)n�I<z
Q*˘��©����]]�����8��]D���L������KD���#yj֬S7/h��͢�ȕ�AI��8�L��i�NM#*�io�y{nT5z�m�dN�fU�P�mR�)�����x����ʶ1�a��b�+F�#"��:kNݭ�~�`�Zf�mc���M�<�0*�L��n1Ug6Q7�(�j�uڶ2A����(�Lu��jk��/H��+XT�*��x��!�mi��`�u-f,yjs��Ҕ�V����.<�a��y�pq�P���f2�T[[EJ��4,Ê,3iB�cm[�\�e��d�ř�&���b6Ԕ��d�4�&ͽS�;5uqC�3`���Rq�bfKT7(h�ufc
�#p%��%EY4Y���3�R�J*�^�S`��X�6M���:%-Q��iR�.����7Eȴ��n�$�n�s�C:5��X���WB��4Z5J֫����G"ɓqբ���UU9(M`��
sjQg���q�Î��̗�
t�.�A/-�X	���U pnP�3JZ��{Wm\X�S�����I[fe���Vر��7����n�i"X��߫3E�õyr��-��&���	$�ی�O"ڗa=��opm�w�Spƣ2�d3q!��hP��!T�Ͱ�8�WW�����f=��t醙:s\0*!�m;ݿ<���lFQ�1�r;Wo+q�h%��#���x黂d̗��n�3�o8���t���ɵ�v��أ����ꄬ�gf2�2���H1Ƣ��A�f�e�F��VBZ֕Ge�앴��5�u�.3!�Bm��"6�dۂ�6�L��u��:f�����*��qn���������{�w�JYQޔͥ�IX��^�'���i�B�h<���8�-������o����Z��u���Y��m[Kd�CJ"��7,���n�������b��b��Q�� �d���]���ʸt�0̦j�^n^-%.���k.1�l�V�Oɧ����a�@˼�b��&h�W�6�kԡf�ڭŒ��Kg ۷RQZ��hZsL�Tn�f�aб�n��wC��Z]*�f:���������.l����7Nj�%S�p*le���	cs5�"e�j�e���`l�r����93�d+F��p�m����4T�Km���Z�,I�2r�N���J#���f�I"�x��Q�5as�wl^�j�=�H=��I����"�m�T
�'f�Ҷ��>Yoi��7Cl��fX�c�t���4�c����*�+6ࡹ�����e�b��P���jUF%�(ltq�u�LI�Umm�ʕR�8��"\h[˵M�-d�zn� Fd�f��z-R�Pai�Z4�{4n%����[�T��f<�ȸ�"PV��]����2b�ܧ��okk��uNXJ�x�R�L-Jf�c�S�L13q�) ��k.J�$ywW����̭)d��&��e���)KyWo���Q�e���v*�ب��e]��3'%]J���b��A���z�j�r�;��ᕐkshT+�]Cc1P�H�#�i�c[n��A[�.������"��#�vRܭ��+X�ȓ���T.vB�ők�܋QN�V�ofٯ��PUU�lI���N�����JV� �4�cY�-f�6(j��[�Z-#8�Y�^V#�wB�G[B�����cQ�C8�ѐK�*Q[���A_�,�L��淓�.eZ�U��.fE�%E�S�5*���*�Z�ѪQ�lj�y��_���@���ʴ�#K3�Ϳ+��A
"�2�X��Ɲ��.�9WJl����7�L`���&��i�̎'Skk!8�mU��N+.1ykb_�f�-$Ff��h�m��`�[5GN�;�ܶ��52ʗ.F,,QVE��b����[{�n�$�LPՌB�
��Օ2UE1�m�b�NEZ������E��*]9��y���
�*:��bN���/i�U2*��E�B%�}fV�D�<�,̕���f���0�I�4^R-��^�M-pA���kYL�j����r���e0�Jn-ڵ� ~n���++)���',��m����g&8UX�!f=p����=���Z��uw���tU�,�q���q˶��N�����5$rPYn{ť阑����n�i�-�H�4�*�'V3�����^�L%�ZS������d�bƃ��@��F��4��Fr�V<x^3b]��}an�y��$����\�K$�T��H�f��ZT��R�Z[M2F�y,���r�W/42��A�\8A�wC��&UZ/ �8�б�M�=.��tC��G� �2�*��<���P�y͂�
6 �J��V���SP��j�䠚j��*�hn-Y���d�����4�1+Am�nEMi�Nm:����W�6�q�q��#s���:uV��{�uab�s����$��4[�iH,ɭ���Lf,W�Ƕ	jx�Y7�\q�؃��Z�bXT�
G�2cl6�fz� �1���ɫV�WaYBŻOiا�M���o89�u��
A:�N�M�؀�ޟPY»RP�b�C�������o
�
au��mp��(/x1���r�w��M��a+9C��b�!"���]����&�<oB�xJ��D��B� ��ᐈ�3lZ���Q�^��Z���B�~��XFV�-�� �0����Z�.`ӂ_����E'��}C�;Ʉ}�
�P�³C�X�n<A�=�u�2����.�u/QУ��chmPyb��i�	4]P@����ê���B�����x*?LT#+�lZ!Ղ?�
�m��,�`���3Ɏ�/(K��]��~6/`�BdT���o�C��A�;`�GT�t��X�g�,����a\�t�����	Av���#�D:C6�^��;^X+l9���Aa",��z�O�C7�X�����C@J�J���4,#��� �@�˸Rc��E�TV,�~�~��.�4|��c���Fily���AH=d8ů�/���X�-�D��)P� �~G�pW���7�:�#�X�!
�<�r�+��[�5b��c ����%�E��0s�v:�܃��$�f0Tb$7h�f?W�0��c pw��3`#A0J!41�0���kc�	d@C6���m����]�A�A���Y�R��*Og
\`�B�d!��,|เ�X;`���|/HοɄ�(�L!Af� Z�X#��pU�*| b��[�K�)A���w�<��H��r�����~|�V@z��q"$a;�U�[a���1����"�^�~�z����ަ2����^�۠V�to1������E���`�� ��GH5��T8h�¯��"!���� b
pjŦ0!d��7P�
X`w���*0� ����*a��VP��c���.�4�\�1�̈ ��h��N�
�
�^W�gz5w���$��-h�Æ�.�]�K��,�����1R�T,@��c�X�HraW	l~��Z98+��l�62��BpU�ubJH�Bu�S�T�f
��՞�pWP9A�ȫ��AI�/�_�s��@�0M���jA�;,^�/��7R,i!��8F-�$��1p���)�/?1��E�7�l�p�׃+z)X#�Q�_PF(\c^ Ƽ�Ǣ�C�W��c(.����	�f��6�&ñ���8s��m�~?{߯��C{����7��}3����'/�3�{�Å$wT�;�1ͽ��]=�B�&�����[�U2���`B��������y@�o�{2ss��/C�H=�:�f��y��E��1ԙ3������e]��v���v,�7j��9"����;��)1QS��H3��W�42�^KR7Y�ŗ8��y��~�f��u4Vwf���}P�@�;Y��R�oq[�V܂mH֯]�*f ����nd����¡�4A;�b��jm��K�r\�v�ڗF:졛[*�ګ�;�u��1�=�vºȒ�9�A��.�HcTpS,���s̉�J�okcj�P(�;ġMs��S��*(scvs��Iyڱs�YtTͳy-&,�U��g9n*���p��i܏W���5��We�����C
��ֹ�d佫�MId��Fm�u��t�a�i���Z�7-w���g>xreX�{1��GS��6jy�om�"���E��B���4w2`u��bL���ۧ��*��
Ӭ�ۜ�ձ��'�SmUfv;�	��6xu��-Q��J�8�;ŕ-�L����y��v
y&�r{}ŋ[�K���\��γ��쪡k(I;�[��F֙�Ź�o�۾�%����;�&�鑃}³^���V>T���{3}f�´�=7C3bs�'��Lf�3^v������3r���r����q��݃�3_������uJ����3�m��ѥ�H٤7nc��ӫl�������V��މ]�s]���{����Uz�t�3:��9�w���Qk�ϐ��g�yi՗��ȱת�'d4���ұ�����n�xTP��۴2����3	����=Eƕ������A�e���;V�TE����p K���L�u�h�K�JX�Q�gfb��]�܅��`�5��A�R�aمz�5�vj�{�ۼ�Ca���-�&u�0����CP.���+y�E�] ����}C�f�3���Y~��fLIE�]�AN9FK��;6�q��ʭ�ɷ���2�U�(��ݙ����M9G)�=֨]�Ɩ�Q�h��yu��*�i2��޽�c�:<�r碌[j�.��2	��wK6��K�t^d���R��p��1��T��I0M�[HX��;��Y��P��_v��St5+��׻�;p��Na�V��![�I�K+vh.)�	WK`������R��
;�O�l�8c����P�<��
�Ύ�q9R�V��z�W�k:�����̎���:*F銚(�y�_���]����ح]�5n��I��.O���hUe+���|�tT�o���-��e�d��֡�]6/��a+z�13�-	�q�5���+y�e
ɜ��JzR�r�u�%�_�T��4^Z���0�vi��6��Mf�7];���uJ�\{^s�ms^ZJ]M��j�ޕ!��w�=mU��͏���n�uw�7�����T�eH�+��YIr��J�=F��j�	�.���8r�}��}�뾙�BpoX���Vx�	^͌1�q�j�!��V'|\�(�u�uˉ���d�'�e9E����я�9�I�Npj�pZ�������S[Sj,�K��b䜤�q* ��%YT����j����ډhܘp6�ĹR��N�jY@�ou��6�ֲEپ��S�rOi���>Hn$NUE��j�����;mN}R�\��Ӹ�Y}for���8Z�޽\B�����N�=bwW&�_R���g7�b���m$�g��~'pJ\�\@o#wم�!w���/����vsоcw�Įcw[���y&�{����nu�w9�u��4�U]�p�E��w|��5�r�EV�T�w������&Z��.vQ�m�y������V�׮Ӭ�h������]�O�����q7�P��ȁ*�P�ܮv]�f�U��B�����̂��UG�wQӵh���*N7uׂ���F9u��M�J)���s�˵�A�c_��f<�=��2ژ�uW{.�T���7�u#v���3���d9�F��MAv2�����#���jVw��[��2��.y6���򞐷6�R�:�>ƟWi޼��C]7[�p;����{�*וI�,�auVx�����U1�����k�m%)���/6��*��j��z7�W�]�%Mkk0��0�0��� ��#l9��u�i�Ϲ��r�y�dc%����;b�,��R�s�l�ちfύ;��3%�-f�:|�em�����Y���nE���9�7I��G��E-�;,9��uE���!��Vn���w%Dj_[Ӕ��cV��r�=���
�����r�g��j-Im��Uǯ%��fF�U�Jd�"��^�Z�`�!�\�A�iv�=w3���X�@����8ܼ�	��z��ٗi�6[�0�T�=o�unX����ov"!o��	Afft �0�x����������6E!�5�v��U��fe�?\�uߍ�G��N���ME&�Y*c����6X]���UL�]�&�=��{d�k��ͬ�U�Ӣ�6^�ʫs���l�K\Ŝ�]��Jf�Q�7r�8��$c��(�"uq�K8���ڝ}i6o��GF�!7���gf������qx�uvh[gC��)�o�6M`��Xҷ���Cvs&Ɔ�.��h�|�r�n\��u�7��ջT.�
�����k�C1[�6����c�o!/�U����S�����yv{�X���t���$��}BWR�]mC���Pp[}�Pm���}crGv�XzCY�jEN�ݾ�Wk�K��`u���q;���
=��.;����^�5_G]�����`��NYR��ˈ��[s�E��]�'����b.0�G�,əu���9;�ّ�u��:�v6�GM1��bV��n����'�G1CFU=��9uU���w1>H�OzJ�{]�yi���>90L�v+N+6���4z�lZ7�]�*�v��1nf=��k�xb��c��t��<��j�&��l���iҤ0�z��v��s*r"��J� ���ݎ�?e�ȝ9j��ݪ��4���lF����,G�J1]?ݙK��Dj�_���9���P�%݊�P���(���p�*�5�g*Ъ3��Y�{Oe$�tMMmG\��j�,��vL�Ç �5{��y�%>W��1�{�[�Q�����t�_[��U��/Vcx���ݙ���Z̲��xn-ےu=�� ��쟨�ܡu�L�}B=.au5�ans���Y.�t�~�=�ynܹ�D)�j���Ƨ^�z�,dX���o�'ڐ�l�i��fV�"uY�~��So:�6�P����n��r�c�������\A�w�8nt���>�WF{m,�B<�"M�j�F�e8ە���yy�yi;;�F"���q�[jY�9�޾U8�I��x5ki�6���o;����[۷�nu�шѧiwY�Dr�����u8�hru�q�hKحs�[Aoen\*^��c��vc�����ʈ�O*%������y��a����t�Y�z��Z�������nX���R۸��ۋ�lעZM;q���A���Hh���~���#���9݈;x3W|�y�Qjʾ��(�<��w����NɆ�Y�3l��9�cR�>Z*e�\ְ�+&֫e�V�|T-��/�U4�uي�*ӥ7�.̒�����>%��em�W$���햜��0)��ǩi��pf_:�Kd�9}a��xUv\zq1˶;�/�Kȫ')�IU�:�j�2\���{��g��4Ty�~D_U^J�-%t��^����nMi�~�iL�œB���0�ɡ�`k���F�T�Om9��]��u�c��v�+f<�D�dLYB�(�6��CN��̻@�(nuݡe��2Us[r��Yoe��D1�8���we�Q��nU�H��wu�Z�,;�+{E-��+U�݆]n`�b����FZn��e�Dwn��sDn��Q�����u�)r��ei�{vVr��u��)Jث8U�&7�9ܷ"��v՞�j/�i,��_,��ȥu����{
��[�{�xvK���Eq���9�buɋA߮n�A5v�E�J<
�.7|(n+<̽��T�Y36z�k4��ۈy��&w5QF����|�?.JX/&Vp�k�����Mva]\]�gN��vNdC�:����w���N]V*X`�޺i����ٌ�����\���ڲ�l�9��9f�ۗt���Rj�[�}.�cGh�%u��V�.�S�o��*�VE��t�C8 �nY�.{�i��E.�����d|ֹd�"�On�>�L�duu�W������ٌi�uZRv��F#yTb3�ް_A)[��v��AB���I�k�+6���rw�o��_KFSʇ�b�BEڔ���tP��v�]1�,֦04eѴ�XBUfiO��b��FfC���wV.t�z��ce�{��cC��M��}SU"�Y�l39�g����*�<J�";��n����o�`q��ٻi���ggo�]F�^�檯(����oqhW9�g0s�Iu�́:��9pE�#�vK����U�|�\���\�����v�,�R���ey�z�2ݙz��-�q���ܳ�dp��euC{PZ�լBRV�a���km���:����Y{4`�P�R��q�8��(��wa��[Vc]@��5���A'��T���j��l]{X�ըT�KEMy���Ew�d껼���G�vվ�oLme������+.�p��W���Ƴ�]��S��v��[�ݐUkJth�m���]����Q��~����=��fgK�e�n�c����R��V��<�6����z+'fYT��R���>���<����2W2�#�&3���D��V�������{ri�8o���+6`��=|�u��A�x�o�A�5E\�3�����б�hr�kK�n �q�J�ǻ׷
��X�3a�x�:�L��+OB���:���3R���yc�X���p_#v��0�ʳ"��]ұE��cd*uS���y��wn��z���{�z��wu=T/�_����pf�@�n�5�tYI96(Ă=jF�:�K�ͤlS���*�t��-�YJ�S�P]�������"���k�坤ݷ�ع��n�p���u��
�AE
��qy��h�FU��y{C"�Χ���cpk���iHc����O��<��IOhv�3-��nj�3]��l�,�$`��$�mŹ�Q�Xଦ�c�;���H�yF�%�'�+i�{��P諘�X&����Sy}�{����ib�Aۊn�FӯW%��i�;P4���f��{�3W[��沕K�ꊧb��,�ᯨ�;b�y���z��."3�\�B�&�sᓪ�,�Ϫ�A�����t��EC����u�r|��� �)�yŐ���z�����kp1�,�!�;�R�K�ķ�q�hR��us]�[��u�n��n��8�[����Hy#W�^e���62ve�Fh���$�N��C�����BSh�΍Y�ǒ�͍\5A�����Ң�=E�a�-E�cݝ��^Mo;�+#�]6�"vr**sf�Gfgs굕6ZO��ir�ݹ��X������'��kmDTk-;��%�F`�,9ӯ����wu������6)Nz��]�oS켣�z�݉;
�!��(�8�VwN���2םN���͸s��T�_.�|��R�J59��4:�}�������p�{��usb���'+jΚ�5����e��8���o
�-�M���yبխ�����$�I$�I$��HуE� ��>=+��:S�׏Uj�t��^�+�=x�]�v�O�cת��ӎ=p�>cZ��קϟ;+�_��?)ǎ�ݫ
�U��z鮟�]�z��8�:=v�ǎ��>Uv����o�xq�_8v�ƪ�W㦽k���v|��>8�ׯO*�ztqӧOO<x���⪱X��v�Һc�n�=N;v����v��n�+����8��ON��]=0��G�|�Ӧ;v�٧N<cǊ��+����v��ǧ�+X�k��Wn8����mp���G�GJ����]=V8�];W8�U�Ǉi��ۍt�lq�=q�:q��:v�۷�������8���x�;qٮ;t����;|��קN�W�޵ӧO^��U�1���Ε��5ӵ+�x�v���׏�ۧ]>c���;t���׎;S�>v�]�v�ӧ��q맏^>x��U��b�q��q�����\q=|�>*���S�v�۷8��ҫ�N)ێ�x��Ҹ�ox�ګ��o�S��1�!� ���,�1XO�7�I����,����&�l���_�g!Zz�짗�2�H��t�F2��R���]�E~�Τ�&�ň�*�?�
dY�5����U��2KD#U5;BXHt���)�M�����-"�}��n�i�(�R�t��8�d�RDЭv4�Mi��A���~*P��n��m�E
��*�.�+�L��S��2�;n��&���<��H=d��=�N=V�k�fꎄ�U��;η`������]��`��B��'�����-�MY�3@ü�;U�*�Ū2�mB	�
�l��s0�,�I�8g-��an�F��b`������?ߕ���~�����`}�����=���h���UWC���=T<e���6�Kh|\���ѸQ1����V�ou��y���g1��<��%�בS#��i��\�-�6�Gm�]�#��m�o�v&���U��[ȮC�ՠ��Yt��{yt�j�x�9�S����H��ݣ�y�ē�)���fk�dw���jȵ��/%M�:7K��&2�9�/woK7�v�ˮ�[��R�KU��(�,�8�^	�T�ݱ�.�Ǧ��s"O
9����se$�]In�PB=�M�*Ŗ5I]4�xՇ�V+v����=�rq�T�~���C
��[���ͫ��4y}	:�ne�29�Nq]:����^<T�5�M��W+���֚��W|y1�$����/�ZQkUrcX˕�*̽U���ћT�ۗ�;��f�cP�QԔP�/0Fɧ��Ȫּczs��Zz�*:8&�4j���ۋ2fa>�ڝ��ٽ٘�T�R�]5�o*1-���8��a��U���D��\�����B�q�ݱu�k9Lq�A̪��U�&���;�n��K[6괓˸�����ee�o�7�:��l���
N븸���=��9+t5; ���9�����fG�B+|��Mq��vLp�~��y�߿g|�L<=0���0Ѧ�i��i��4�M4�M4�Ji��i���i�F�i�F�i��i�M4�M4��M4��M4ӳM4�O/��~�k�9�!U�2��v����+.�,��br�T��\y�w��5��u)���*j'��>-�2���n�Ol=Ç�_3/�}�ϻ��	�Ϯ��|�j܃*��]z���(�aSy��^4�o����)o*D��i�ֱy��胖+_^���$��e9���EW
�L�^��V��Fua(�{(�On�%�:n�pS�F������R�R,�Y��}T��'(.5�S9g_��I��j�v�M)�r����w�V�w�+e��Z�Ŕvɧ݉T���f-U�(�\Ц��;8iWĬxy��&��2�.Ĉ�W:8����um��o^J���!%*�\��j왈</���g���7K�<�1+��f��bun�$���]�k��zz���u��[{���t� ���SP�S&0��q�c�g���x!9n�\9���u2l.����1})���CkFc�Î���A�3���0mZ`����5�(���!{�}h���0�,Q
Wp�����$��z��dKK-����p�rj������"�Tw*��<*޳e��0R>"��oR$t*�AII��̡�('B����Pƽ���f��>�_���h�NT�T�)E���� ��!�����s`UK��9��)g`�α�XB]v9�;@����&��  �=4�O�4��i��i�iM4�M4�L4i��i���i�F�i�F�i��zh�M4�M4��Ni��iᦚi٦��.�=�+W�0Rv ��v��h<�B�~�(z�P�u8�"�@.�=�����]#O�!}�!A�u@_PD( ]���|��# �1]�{�%����y��a����o�w�Ӕ��-��F�[CH G���s#�uW��}z��Y�;'t�޵����ɍ����V�dz��!)c*L {�^��.��0��t�"�3|��1Q;}�>޻�-��{L����=��Y����6�=��`�z����zY2�e`��{���C6���(��	�w^P7���!�L��@r�BL�d��C�E:�ֆ�c��6�:���MyW�;;����K�G��7!X}�T�����fr��t�G�m�Z��� ,+xA���u��,�-��	@@y[+�J�+��C��r��t� !��0ABp��D�P.��yܡQ�66�����=�ĝy��C��;뺊��*��qs��1������جV��hS���Ռ��B�(?,jt(��0�����<�R� ��1��n�0x"���{�����00�*��������ZCl���+���c�Ú-u�n$��H�h�D�����;�l����Z�DEj����+sXFǼO��o3``>��C��_�x��ٚ*f�Z��зCU^�َ������8 ���u[�JUa��պ��,Y�����;$�S��͙kn_`�:�2]I����c
Ȍ`�}]�V� y����Zaƭn��]'�f�/�E���{ݻ�����:z���Y�V���$fu�A0�,�)-�L�Y�"�<E���l�T��4�`@ a���i�4�M4��M)��i��i��4�M4�O�4ᦚi�f�i��4�M4�M>4ӆ�i��i馚ti�)��+0!��	��,�nn�Œ�Ě���V(R�q��/%t���d���>u���H����0ޞ�=��j.������",�(�nw&f�t�� J��}��㱩�f��z�vT)=���.htXg�D:�$+:����rR�ܪ7�E<������S��z��v�))(����y��5��/��v�K��R*jځ����=�:�ęϙ|�
��uA╏n�]>�> ΎRuC�htk�
��39]ﳐ/=�i��#ܤo�o� �A��4�Ңd�ip���uW���ݻ��ĝ�k����n�U�q	�p��2����X������o��PTv�����}K��r������=�X���J�����\�a=r��Э�],]'�d���\�\�.n�fu�.��H�yԜ��P�k�p�̓�K:\f�ne�=�}g�J!\K=�ۺzƚ(4]��y��[�V,��S]�+�֬�c��E��֫�k\���M��y*�{��N.����������#�5Y�t� �B\�l뼾U��2�יH�f��� &�.A�&����̼f<H<���w�z�u�\��b5�ݪ�_8�q�3,�tr�ՈZ��#�#�U<����P�ʴ]:ESͥt�����]�:b/U�iu��~�L��%^��F���0�����?4�N�4�M4��M8i��i��iM4�M4�M4��i���i��xi�4�M4�M4Қi��i����08 �@)��������8e'��lU�Ҩ���t^�uK�-N��sM5:-x�$8��F�L�;���ΌZ|ξF�8ԦmT�1���]�-X��Ш�6��3����rek}�8�W0�i�u�K�����z��k���Au[H��˓��c�Ǝ�r=}� �ܻ�{�+E�x�$9�\>����׏l��S4���sު6wa�Ouӿ�;���fFƭefKꚀ�7=d<�
ncl�����o)��ܬ%3�?��R6�VgM��.��1n�ӭ�ÐfF6d�
�ZFc��-*mv���\�r�9g�o޳n[�� �Y�B�GQ�y�k�u\޵�jP��c��qfN�*ګ��ں�î�h{t��� F�Ȧu�&�:g���30\h.I7�"���a�������t^(�uqηQ�{ʄ�w�����n���Y��O����E�����6�JKY�u���r߫��L`+n�P^���g�#>��wv*VeE�r�I��8G�e��,�S�IX=s�ef�>��	��J!r�g	]7�aX�6�[:��k��ٚ)n�>�28��v�]ЮL�^y;�g$e�í�|g��k�J�J�qo@�����R�P���$*ڋ��y<��d)ΰ(4��񦝚i��vi��iᦚiѦ�i���i�4�M4��F�i���i��xi��4�M4�O�i��i��i�M �@����ءQS���`̼.�v��n�b
���z���"�c�/�-\ػK�3�1~�Ѽپ�%t=��Le�db����Z+#�Qep����e�33u�a����]<��C�)�ø@�����M��8\��]	gUF{�s.�β�<bU�E�Z8���(/�/����Agfu�;bJ��@�.q�r.)/w4WK�.a�+6^�v d��L�Q���]�޸��a八���sNMEm�y|�ߵ�Q�2U�~�f�%J�3�����AC�(���k�;������k�����tmU�g;Vk�B/3��D뤪ц�ZD�j]J�\�9�J���jI@���Ø9�M���(��7�03U-�-�K�\}�;;!{2�׮��1�!������9����եG��lb����`�yTǦ澷��M�����4Ӣ�>W�Ш�(/-���פfSxnGuim��[�٤�ǀ��Z좹�32������I
���,��}�n�{BC�%��pk�$��G:u��}���$vQ���W|��<�陕ݥ$��u�t�=Ž
�cZ<Ũ�{l��g�s���jLE���c�Զ����7ig:�r�����H�6��`�X��i��iᦚi٦�i�f�i��i��i��i�M4�M<4�M;4�Ni��i�ƍ4�M4�M0ҚiM��<g�[��	ؖ �.�O[5k5ǖDy��Vuc����nwqo2+4�\>u��ۧ/�{����?m���]��'x���G�.�,�|P���+j�hy�*��s[�P�o��9�Mo�Z܂�W��!ZG=�}�M��Ƥ�;���0V*'�0t�|Ǖn�W�	W\E��1��y��#�Io��l��Wd-O�I-
�Wք�N;tx��һ�������y�%J<�/7z�W�Y�aъ��sD+w�îo$6+���];��S*J0fP���֙N�h����Ge7D�󸂂:U79�Oml�˧qٵ��:�C�MV�#W{}D#-�ٰ����Xp-����v�|'��f[Ŵ1�(��|nN}B��:�W	�:�kc�v�1+�W1�*�uAt�S�7�WS/:�暳�n. �j��|T��5�0�#����;1Wf�}ҫ�7j��f�y�ŗ��:�3C��<�J���=U�W��ؐ��"Z�7#b��-���Ge�.�&�cb��T�N��Er��n��u<7�ŗ}�<��G���[����Pv�m�[�5���zc�����`�e�m&c������f�M��8$I�Y,�i�cDK1�d�F�NV��o�ձ�����SyΖ�EF��J��O�>0��Ni��i���iѦ�i��i���i��i��i�M4�M4��M:4�M:4�M4��M)��i��i��� r�P�Vh΂�gt��Ad<<5�(n�]�<	JO��>�2�䞾���ty�*>=ԋ�ҳN�+�����5��M��f��w*>bU��_X�{�����=:��u0��%��<���V{e��Q���n�h�[�)�x%gd���!ҫ:�aYJ����f
w�y��zc'�t@MXQ*@5�N��I��U�W�X�Fȝ�u���zV;��ku*|��eku�������=�g\l�v#�����4N;����"�ٻOnٱÚ�Jqv��m-J$�R^�D�,��Io)��QT�u�2��*8N�V/�,�5c��o��\T<Vs�TܝB�r�OH}cj��Qh��Z��{�UM�ɉ�ۮ��gl4W%��跓y�ٔ��[��[�::y�+�ӐIbm�J[b^E�A�W��#G��nWM���ŝ�آ6;�c,ur�zՉ^7�!C���^�v����w9v�nK}+݈s��\������i����k��KwY;���8�:��;�ӱܚ�֗}V_f��r��m�b���/MTy��e�x�����̸d�r����y5�>4b!̵Y/'Y���ĶF+��sk�.�mβ�י�C����JҪB�܇�B��/HV4st���=&ڼ�MwNI�x�,�n���}���i��iM4�M4�M0Қi��i��i�M4�N�4�M<4�Ni��i��p�M4ӳM4�O4ӆ�i��i�F�����כ��g�Ym]�B�/�so"X�"��	j�Y�e��F�yq>p��1v���u���S�\���h\�m�r��1�$DO�b�U�<#�gK�T��Z\�1��#x����;�1T��!���&"�.�8�Qy����bR&n�\͂���$�^�q[�o.s�bF�]�V�����Pp�����#�2�-�w�c63-�����"|z�^DeU*ֆH��T	�a��n���L�S[N�i��r�ގ�
o�l��EV=ܗ�-�1�&��¸!h��s(�gt��X�Ȥ6*�z���LT�ػr׹Ӧ�+{�x��&�[�y*f�ۻ�5���,l����;���: a��a+��Ʋle<'����R8R�!ד�:ĘO6�]5�}n,\��[1�[�d�Xv���wĮY#��	�����tX��ҦK4 m��`�R�m��y�K�1JYY��Nx�4AY�(��Ԇ���&�i�t�져�t�5����}�5�Q����n��`�� ��RݓVX��7��n�*jJrR��D���p�Yb�.�7W��f�η�bʮv$��,ۤ6u�Nᫎz��//�ӝ�V���_�D�|{3j_A[W��.�R��͵x��#8k�V�PƳ��nZ$�a�Σ�Z��_0��6ir�<��s�5-�P��2�^zw��uQw2�--Lj���h;Fn���(u��E�M�vaɓ�K̺�b7�{�6wx��en�WhY���خ�m�d�c]]�U[zk9q�22T���H�i�Ɏ�%[���e_[*4^Yu��A[��4s�;Z�z�P�녾�ūR��ӱ.�]?^��vV���Sm���sު�Qθ�ȁk[Z���a�ˬ�}����Ǳ
���Q�u
��*
:�mq]U(�Y�X�R�B���z�(_ds��v�����N���c�J��3�{X����$Q*��ʢs���WL���H��kI�+P�%F�v%���6'et��"���[���Rdfm���.���m�TWyM�6�]�O&��k���D[A-�-��,�ư^N3��QꡐfCA4)�b����%w\X&)�q�e[���n��5~۬���1ױӢ��G��;�5��o=�L���J��=bv�)���uX�lשe�1�m"�ꋁ<z�ޓghtٕ�w��v���5�W��ٗ�j�m(�@$/ߟ|�߯[�|�~߹�_���QU�俻������?Rp��?������~{���~�s���Ύ�g�A���5!��n���˼��^��ne�7WDTM��^����/d�L<����5���ʝ˺^s����y��&K���a�z�y�4��O�,��-�	�'�:;��w.�E�2��C�m���0e�Ъ�G�E�x��KS}���Sɽ��7#�h�Bj�5l�n]u�`�L��W�e�uKX��]+]�[Ǝ>�5y�Os�YzD�X${�&תЗ5b�wk�����:�^�;�����n�3�o��^�p�H杚�Vs�0�X��^�N��%Zoƶ�����gE[I��㾺���Jڭ���o#�{���m��o{����w�w���gh�4�]W��&��_��f��@�錇);���@�*ȫxsmK��o���3�5B��&4z�Uika��f��u�Y�+)8�=B��,łhp�W�.�ڵBR]�h=���T�+��
��D(d8���κ)�v��Ua�����+�[!6A�+�A��Ķ��l@޸m)ܶڶ��*����\%Q�q�d�%�FA樝u�)&����F�ֹ�t��q�(��S`��t�۪:3���C|����t�wsN���e̙T�_NΝ��wx�`BŎ0��S^8�ox�U]��J�۵q�q�n��U;xcǎ�q�q��O8��۷NΊ���DX@�8!cL�����e�ް���Tku4hљ)��IX���\%2�[Ǿ���u���6�aOp�j$+�E�T��E�z�Ķ����9ԝ�]w�ȧG����CM��>q�
)<��hk�E��э��^���3h���Z��4$���8ti���M�l#�k QCB �(DЎ�bh�ȶ.b�����
�hC�F�B�P�:Ѕ�F�h]�F���@�PPQl��7�q��b�(����b�`��Xh��AG|�����kQÁ�����M>�<��+����x�A��cCCE[F"��<g#LPb7X�G�:8A��=cx�Dko0scl�l`���clh��AC�JS���?0��]W*�ʗO��y6�������Fш��0p��yu�"�{x-�km��Iբ�c�lA��==>4��o%�W6�)c��1�^,LQ<�EZ�2B	p6��AVBm���JS����M4�b՞6
���4\+�#���͖����lQ���s�т�ΐ�<4��L4̝{��ܲ�V�d�Z�c�S]���MYR�/q\pᦘza��j=�}n��1A���8s�i�AS%�^�� �
�lZ�UL�h�`�(�jb�A���4D{��/�G{�sm44�|L���,!�91��[S����F�����O=�+���*ׄ�E�x�f��yp�I��@h p�D� ł)��0!kT�J�Yp�`1UF�J����q�����)���+����/������Z�Ƨ}�m\�9�EL	��YA>�H���Mb�;�3��Z��s��k����<>.]��d��FN[�&������ܶlS�O�"��U���@m����`}X��K����.3j�Ŭ5�oPå[�. ��܅��5m@� ;���U:�Z%��8)�����ibf�	��EVҬ�y����,��_1��|r]����zYiƽ�Z�ϋ̅��-�W��Lv2�0%��	&.4�3٢�/F%>���mHNlm�b����S%��^��k���kM^�Y�*jt�: ��[ġL 3�4&2���|7Ա%� +dm���3m�b@͠�aXw�P������.���z���������N5{t$���צ��ݿvb��$���֪�^��_LpΝٟ\i
Rv����k��sN�1��4� �1^�#���XڇI��Ò��4!���ú�S�y_v�=�M�o�e�Vҹ��^�s�6q���_>b�UL#^������쯼����!�@&`�Eq��+���ϕ��[ͪ�t*-+�G6v��c��e���x�|}�t�X���}s
�Y��٬���|\��1۝qԽB'�텆��[�sV����V$����)�t�@���
 ���VWJ:
ʻܙ�.͓rJ3N�,�\�{ ����hn��;F�t�1�K��z������|C#
��	D
~����>��L���7����d�Kk���C���}���Wo�Q��^)�Ә}��-�l�C�m�z�%��3.�E�92-m�2��W�~���<��p\�6�FV�;� ��*e��J���	�[-�͆i�N!�U���}k�Y����[Z�d���W�VH�rV��ѭb�V�"alت0�3�}s��;׮��}��Z��І�c���0���Wk�,�:��w3�$'Ռ��@�o��P�Y<�wr��f
x̔�����-�p�ΝYѺ��*u���n���Љ���ƙw?�����y�TI'C�'	�FK��Eao&9|�Pan^Q��0&����ޑ�T# 'S��Z��6�"�s�34��h/m���U[��A� x���f�N�+d_�� �[��.���۬?]wE�㘤�^��,��e�e���uy>�T}�~��@da��
�k���G���+�MH����v�bt�6��z(�p��1>��1*�%0m���v����b>���{��{Y�t�>�����?_���ᠴ�����׶�k��F��}`o���Ǽ��'_���$f'5��y�[�ER#SY���B���{�l /��g��sO�t�J|i��ͥ�%ml�27%�+.`��G~b�cA�a�}׫�<����)�=TX-uF�㪲���r]A�<�'��<�WގUTˮ=�ɿfy�]�ښ�Wn���8�gv�&랹��Åvuδ��*�}=L�d���gO�?�����t���x+-ztη� }�_S��]�%R*�]ܧm��vX�����F�d+�r�oJ圳UV�X����>����0�������F����i6{��P��S�z@uG���+B>ͷ�<�s�}���3J�#@���Y3j��l���������E�BC%V(}�G�����ٵ�i�T,��FV�Vm+��K țƤ{����U^����_W�� ��S�b�o�-ɺ�6��U_�1�X�P"gѶV�ZL�$Za;z�dc�+A�I�s���[����Eyp��y���t�'��������c��4���}����9ԕU�[  V*կ���,�Z�Z�"��x&�Pd?�@�-�x_\>\ҩ�������׳qI��	�*�c`,�}oc��5d'�OE,��ur�2�[#^ثإX�F-,)���	^ZIi� �4v3KF^J�	��9��}�|W�g�2Sz�T��,�~�v�{&��
��9��{�n�,y���<���EةF{j����w����R��.���B�kP�N��+j��AstayV�i�o����]^��x��-~�JB���S���"><�R�ܫR�S�Z҅��.v��LFCН���*Q_S��uH�e�Ph}o����0C~,_���hVP���5�_0�z��kjX^�q�m��%��p��M*��5�<=�v���fL��!�t,`�w�e��Y���~)��E�V���c����Y~�� ���c�Om�%�̵�Q}�tl��3O���L0�>sh�����,\�@s�+�Yw�P\+H]�T�����uf[�T~@e��uo
\a 抰ӱ2ԯ_��d;��D��	I�
�s��M����c"oI�������z�6��d�Tc�漓�����3��[�[x�a���e:x�2���z��Pi{�J�J���y�s5�kǭ�40*ߖ�����lMzt�݉��5Dk\��+2�V M�4!�r��-���%w%]�մ�|3L�p`�z���c��RaPG`��U�S����`l璳4���2�3UK<�L�(p�}*�=�6a���AF�.�xO]b�˯��zpY]�����,\jZ�����d���ڻ|1��c���|E��c Ay��fk7zT!�q��*����]fn"I��fR�U�������ſnK�y\�u]��cD�d*5�;8
.���uo�hY�KrJY�	���8����4�[�Է�<����V֓ F��k��t�U�����rE=����㊑��j�֦Y`5��ۛ3��pR*]'��M�
��V��J��� �VG��"=�b1�bҭ��5���C�r�ym��3��We{��w���p��\!%`FY����j���.����M�/�u0s\n��6���{[0����JB�M9��dm#��[Ϩ:@�T{��ٰt��X�Dm΃��r!;���j��zuuއ��R��� �S�)��F��R<E]a�7��"��];�Px�T.6��B����`*z�.��1�X`aaǽ��R	Q']�S�� �k������G@��pψ���䦢KZ���8�z�p�ͻ��pñ���Tj�B�>��]Fn�l�Y{x0���w�HƝl��]U�� �msX`7�3���.�)ذ��/fp����:��4��{V]quc��M�.�KwU2{Լ<t֓��ۀwf}9� ��s5�k֨{\
�G��D=��N����~�$�����$���J�ڧxжUG��6�ϒ��hɉJH�yc�����Z�R,��m��]� ��^2�ff�a�0�Mdv�ڨ�`0(��h��%�8���K}�Y4�^V��9i�b�����k�,�H H��!���S��f���fXK%�ɲv��Lmڂ�S��&H����l'���4�(b}�ڒ�[��^�ʱ�R��G�[�U�����}�ϲU}j8�R��7n]+91����r�|�w�a��d"�׌�~Wu��R�:%�\��l&���6��7^ݩ�M\���D���vEx�����@����߮�JO���گ��̥>h�>Y��L^��1��B��{�f6td�	ģ�܇���6���c��9��y��1{-)�^r�D}yϲ�{�\T��;)��.�%��x��Gb���+�u�1�C�IWbok7)��8�Fc�������$꬝�y�ٔ���8�tJÝ�3�QUßd��v���(E��0`}�s�dx7��m���lTX�fC�#[��8V�~bxl��5+�g�w����<�u��ξ�P˘�W���]���40��R����
�O�yU����B�J|�#0���3�>_8�|O�ב��̡�}��h�x�E�h���̋�-a���fN����p>����sr?��̛�G���l�?����2��*�X��n����f��)ϻ-h<���W0���f�/Z�,�tf���\L�uR��{UZ;4g�ի�	]ׅ�r��Ο˝�xĝ�T[��p��H
�ǧ_� "��>E��޽EyY�q�pL]���;_w'i��������?}�T�JAۛ��=����־]���	�/�q&)�ԁv#�I�$O_�S�~5k���4R3���� ~���K�<�@�:%tW3d!b���&���I�ñYݤ��;�sY��#�����^*��̰H���X�d�j�eK]YYDpmww3W��-@n�Q>�ɋ�-Z�ζ
�)R�&�8c�gKy�,
hcA"�(RŔ�:�Dz0!h |�j���8$$�f�Y��ςZ�J���ɹ�kì�Y��֨x�������@C-���dl��N�V��� ]�!e�}U��9KYG�DR�!rr��`M��qD�-;VT��t���Y>ѳ��f�n�M�ڍ��l�u��!5�E]p0���wu�S�ۃA�Ҋd�ݧ�3�����ȴ6�e�P���U{�\{����5I���#T�`>O�Y��d�,؀����B�Y�i]�h��egp��HX�`Ɗ
�Ax��V����6"�e��*ZH'Z)��U�Q��	��\��lG�,֙����1�+�9�P?��V�޼����$X�O����QQ�w#n�y����ѩ�|���/��6�D� ��2'
S@{��b�w��r�zb�h�W^��N��X��ӽYrOp=����3w˶��m�er/G%h�.�����ww�i��!�("$m�(L^t5�e1���V��/#�K�vi»��R�.*��꡶)�Ua���`�LvqWs��R���(`1����v���:L߉�u�,�P�8�1�=Z�,)�FX�K駙�w3�U��
O��ܻ�K=���%^;��g<��`�8��ت	�FCVE�rwrtI(dTy%3��8��0��~l-y�­D�%j;����'v�U���A5q ��Tx�Y�V��$ר�j�$"�ES�5�,7�!Q����}O���g�S3h�����إ`��4E�����j/��Trҭ��lI�i�vh���R�`ff�N�J��	�y��ИȰ-L���A8HK.͢o;Ui��ۻj*h��>��s��c�g���,X�Q���ڱ[1��|�~����ퟶFW��}��QώO&�[@�G}���` �;��nޡ�tr��QǠg՛S<&S���Oy|������`�����$X����}U#�����RZ���
��Ӎ������ֽ�ꯩ�����-����\�Z�o��-��(���ӈ�]��z:��n�a�˕/J��v�R'6�o7�^���#��ȼ��;�����5NZz�K�����ʥMG7Tkv�*����˫c$4���7��U`�qcʳ�R6�eR8�x��;X2���7��B��2�w��3W^Bk�vh�Ξ�����j4ސh7[��Ǯ�n˸�v�cz��,m����u�[Y1ѮS��۠�3˺i�"�G49Vz�oW9SMřO�g5�"jwoE����D���vF�����2��&��iEP"Oeԍ_&����:�E��t���&j���\��`�U0�1D��g���(��-(T�]�����m&�'E�d��;г������fu�P��K�MT� ��Ɉ>�P�A��[�tE�0��Ua4�nd��"��P��!GW�2���A�We���7��S�b-ז �W.λ�n�t���x�iGJ.�}�+$�5a�m%�*1%̬@�k�p�SH�ZKBq�㹜[[-����z�Ϫ�E�ye@�2%t�N,��cK՝�^�1w��3Nlᆑ��;͵-��;̊�kk	Qs٭eu������C���l��`̟�\ ��,k�"�@E�����XV��`�D�l`� ���V�'��
R1TB�PhR��k��i��f��zC<�x��^���Rte���W�*;+j�\߰��ᓌ����S!��<��YՃ+�u����s��e�Y'��d��>p���:K��oH��P,<D�3��QT����O��+�Sƍ�)�X�\-��Yɘ	���d[�q��j��j�j���Ap_K�m�)W�p��=�Z��0^6V��]�K�>��x�p%��WQ+;�Q9��sc���T����gG�����&u5��+M��vs=��3q%�s�*����V;�x\a��0U���wΕ����Z�׼:��Tj���6��ޝ]�/�SZ�]�+{���1Y!\�]Gn���D(��*�9T7�mmF䉮�\��b�Νm�/�_�*U\M�;�����Yy�����Ṩg:�;(��V�"j-b�v>�X�f�P<��بq|7���ܕ��O��q�X92�Q���;f�%��;�*�ܖ�K���^Y��}��*L�q�;[����Ɇ��G�0IX��[��>��y�A���A�Z��9H�.3,����]��Y�D:����KW_%�|�r2��ܑ�l���yk/�'$���[׍+�z�o�v�^+^5��bƂ,1chZE�7����9���u|?���URX'�F��lRiq0_N�r.���.m�j�������,[m��/}s��`�V�j)�*h.F�o7���׎q.㇝�L�U���0x0���O�U����8��V�STUxS�'[�j���l�,Z���?>?���O��R+բH�n�a�����P�QKQU,�ڈ��tttz~�Ɵ�bʽ�um&�=mM2u�"f5���1��ų�xwc���:f�i�[��o}u��W"�Tw��V�%���w�\��mYj�4��٧ƚhvvw�RQ�7�G1��<m�͂�5ͨ��9E?1��c3U�Vʿ�GGg���~�����4S�QELU��Z���䥕j�f�vtvzi��{����j�U�*ޯ&��<c�d���ɉ�)�h�uWx�MEO��AS��֊�K]��MME�_�g��W�
v���;�e�vۊ��œA��S����+c��s$.�>)�wW"��]��N7PK� `�y��<ζtF_�	h�L�ޱ��X������=��<g���&�����D�&��R�S��i�i����A��~Y�v��p75	q��c3g�s�U��5��P���o�\�?n��@* z�E]b��d�;�����6�����1^N��06N�;���n�W #B����,�_t�ˉ[qD�Q���� ���\�܉�br6�*׹8�M荟z~c:�΢���S�xeMv�͍����8�U��눉�ޟi��Ig�Z"��EX��)h
#wb�
�Gq�-<7z܆M>��M̱d�m�U�Ki�>�?s&͐-z� ��u!K��|L�v_;�sn�`\������|�t��hH�]9$p͗h5�0���㝙��3Q�m��jn�fH�n��3е�F�"�Q����X�/|(_V0�=qr��"�aγW��&��w}�@x���~��Z�$�aH�;�u;k�ê=YO�#;i˞�!t�Ʊ9�O��t�P���|!�>:t5�韾L�ewO�j�g���w  ¾g<LK��mo�[(��贮��U�PW�5J��-\��*�Bi]�l�9:�7L���ڳpiʃ�<�`�Ä�@a��B��[sy��N����%V����z��R��+3jF�֮K��ۛf���`W�-�B�jk-��t0�� Q�Y�����u랞;}��j��?+cg��r��<�d�/7�%�Iq]�=�k����[Q_��A�l���Ɉb�����^�a"f�z^K���G��2d�\����b��3p��yn��G��k���]��7������׳�p�j��ɰe��W��}+]I�&����3V���<i.��<E��\�q�xȶ�V����UV�=2lN���mѵWs=I�WB�Y��C�wnur<������F2}WB����LkAL�����D3+��/υ?��tJ�O�����r>Aj�����(���@��L�?=��M�uEݭ�z�|@VI��ܥ���6���*��a10���"'�G�=1|���PW�uǷ�Xˏw��S3Q��i�WA�L�:����MP+��L~�~p*��,��7v窏�>.�X���; F&�0�^M(��� ���~4(�צ$��-!�,^^^]"���d\0m�F�-����O=ql&�SK ��}F�D�oV�����t�1�|�OUmr�B���X)&�<ݫ��UNX�Jl6X���c�e�l�=�R�%�_P�ͩ:�]�2�6y����;*���H��2�N��[uN�p=�}����g=��s�!�U�'�Nj#ٯ(�y�(�6%:}Aݻ}r��=C�40�PA�0Og9�yz�=��۩��������I�����W˘��`�hY��C�N�����A�c�m�D~/i�k���F���9�.Ѣb��L��&�8��-�L23;� ]��k�0�S�O��o�A~5����dР��E�G�xvsOLc�X�]"Xq��!n�q�7�K���j��c�Y�2���C����όa�lx�V�f���X��=Z�]Ow���WF��ǜ��#�^=��k�zmLRq말�m]63��Z���;��i`˜��0���Ȁ��Sͥ��M�8�m��{\y�\Y���E���Ǡ!@�_c��|NI��b��Ф���8��W=f܉�83�k	,�<χ
NŶ��x���xR6ݷ��y�"�)Se�K�ml�t�Dbu`T{`_*[�S���.~�	q�|	�k���l!e��v�(Q̽�{����e�� �0rHXA�yn�8ޜ��`�qiĸ���J]Ԭ@���N=�[��f �b{S��ށ_a���W�%��Ɨ�<�8���Ύ�jm���Kށ����1���LE��`���g�C�:G��Vr��a��+�|�t�������um�y K82�fo^2�>�|Tw��Vn2��p�]<<4��O���i��D�W��b�~��}����hJT�|�jq�#x��Lt6GJ�����s,��Låk�KmV��{�9������~��>��uO�ǽ����.�gfa�_x^��p�H^���TZ���X�����@��L�
��aV���]�*�(x��fE�;@���<�ց�4�G�@tA��e�WF�@�8@ߋ�D�ｴ��>�w���Q�s>׃P�-iE���>��#��i]x;	�p����u�8�s�g?�	��ɩ�,{���p|���9���A��AR1�$�mb�����W�noc��F��5��;�K����t�T8���S���xjN��@icm��˸��:	l�X�5��ÏV���ˡU�}�I�h�򁫵Tl��r���?3P.'z'���;Ur�:Rch�X�� #C���!��Dp�7�MSw=�E6�vV0�Fd���~���k���Ј����T��C^��5�=�	�1���a�^y��wX���'{���'���}j�8��g���Ux<ưp���2=��@�Ȩ�^[!�G
�-�0|廝6�wOk��p�����V�������?�}$	�vv�,���q��|��ܪ��z%:w�>Ψ
`q�X�J��9��i��ؐ��i����%�f���A�sb����֍�׋Ĩ�R�^<w�N���'s�7�0�
 ���z�s�U�Φ^4�T���
���O/���O6�c�����ut����ݵq2�[�p� h��'�𑾁�0PPs(-.����ϑ��ܶ����z4���k?�����H�p+�}:6G���C�3����]/�_��GA��ek��Nd��{��}�QOܾ4"�Zc�S!�,��ǘM�I[C���E����ڬ)�4ǒ�mM�P-;�`��z�(�(T&�~5L��(l,)��V_��~���~Z���_�v���'���Ӡ��/��`���\��1���ݟ*���`�)|5�ՌxA��Hl��1.����t��g���H� 2}��P��k+��=�Lx5�v���^��(c�e*�e�L�|	`} �4>6���B��>��R:�D�z��ٛP9�|;)��ZXIF���>�	�&-�d{Ūj!�q��6��ʃq6���kx������&���C�ۧ��J�X�P�,���	O�R�@�Z�)��ؘ�YWQxH꫎f�%E�˳��ɄO����𤟖5d��5EȦ���������֘��p�E3[x�`��^2Ie������d<4�����`�i�-�R�z�H���y��(���jT�a}3��W���A:w�m��|�H�u4o;�"$=���n�o�=�j�v���)�7��I��u�c�iV��Vw_z��R�t��l��g1�osy(�;|��u���K�NJ�8�F_� ߕY��[B�?��Z�ԓV��3O�̋��o��@���v�z-�����t�^��E��:�[�Ž��kct7��я���_U�� 03g�����?|��&��l#��M7gF�D+T_�w�fW����vǩ����������/�Ӑ��1�����71ϻ{Ty����F1��IS�	��V�˓����TF��zr5���`A�\���IK��]!»!�xvJ�0vy�ޖ�
}���ފ�'�,�K��໻cf��?k��*nD�}��e�42�1Cr����կ��M���I�,���_��� ��_䬆�=噙�y�P�ݮ*�o���)�@�"�zK�.1�W������{ �|%�MɩLX�e7WOX�y;�Z顆-�Ǯy�R�4���gd[O��
�W��OL�#2#�N;6��~��:k�x&`���vm�u��>u�&�sW�>�7^�c:�,��,�,�f�q�{�\V:�����ش���b6:D��0m5�a��7P���{׊-����w?�:�N+n��m7�32�ew:zNڡ��qohǎe���Fp�:9,�l�����5r����1�Ǽ!�e1l���Mx����P��}�u^���v��zcɌ�!Õ�E=�9̧/�}{VJ�D���q�)ZXʄA��!CAH䈢�n��n� �4r)b�R�))R���k���be�����T�'��b�y�Q-����t�����G�[�~�P��X���dD��N�/c3p�X�K�f��_=�`ޔר{����˛���+����\��0���ɲ��M����a�C��=�E������V�����!)�q&a�ӿ�L����s4=:�x�:qr{�.���04vŰ�o(��t��&T���Ӭ%���=,��E��]w��S��ލo��y����^�\��{�����t��Qz����^-��sN4�7���c�k�ީ#�֎���g������ߘ������1���l�y��?k��V�M�����O�&�c��fP�z�%�-�%[�<(�sE��ݟ��?��]��6�Om?��̓�j{���Sqs���^7
�n�=3#b�����1�5���7���b�Fx��|f/q8 �߄�$L7*�'%0��RK�����|`���u��p��o��x��]-��7*#��m��͘壞 �u��b�j��aC�dz1�e�����Ȧֱ����W���>�ܬ7im}2�쳨���=�O{�*C"2���/e�X�U] ]��v�#:e�ڝ������D"-���/'J����m=�+�!}u�����C���pV(��Qi;H�\�v�si����1���Y��[�g�tW>l�~y|�I�)���,p�JTYJT�t�W������֮�p�o� ���;���W1������W�9?���#�S
v�����aY��Y�}����|p�fQ�ސ����X��|���W��Y\D �zfVD(����i&�z4�n�'�	���T~8,g�`�հ~?�W���L�acY����&��ʚ�U|j�>���U�2Ra=��\qr=׊�A���o�A�� �yF�&�A?=yɓ��%n���s���;��=��~ߣ�HQ�.��5�'�~8=��Z�n׫���}9z}�	�pT�7߼[C��i��D�v�v�償҇���;��cc��dr����<�mF���	�kh��ߛ������w��?\�k�ϟ�C-(Hp��8�ٷ�e�g�mVb��._��G�"/��l�}�Qs�2h�^��j�Ӑ G��o�|Pp�.9���|�W�8��O���wLO�]�"F�R.4�J�F��L1�A��9�s��^GDS>O[%��U|����v`5�)��r��V��̱w۴��-ٸ�J�EL���w��1����M��+��w������;w>���j�P�C7$���7]q�v��qN�Dm���%��/	{X
�!0N�Y��1���@d
�
�}\;^���rB��淃/�9T�ַ�>�9�}�ͨ�q�	#5}ٱm�sy]�����M�[{��_`?P��V4X7��#�e�|�xV��u�ӳ����@l	��S a����d�s^����Y����b�o�r�� L�(9��T�w֢�	���\���6��4Vd�w?��y�[ U&%B�*)���9>����PWBX�����v���x&-ǔ�� {0\j���O���CӢ�M����
C�ꕏ�᮲�C�Osb�u�ՊÉ��k���&.����:`�zU��Ϡ�����X�]�1l��E�xKwUQ��)��w�A�7�3@�~�a���>�9�ſPO���'��Ѹw�gr��_l�[A�d4���5qI5Oq@w�R�����p�#'��uƆ�����lX���	yO��T�`-�vj�M�1MN�h�l�J��,�l�����^p�BS�%5� ɘ0897�e�CTw��L��/u͸{�m,�0�{��7���a�w�+�XL�ܨ/�	��C6���`z��U'dczn��*��,r�\�ÅO�b�X}�;l�a���)��yy��&"��V�D��;���Cc�r�v2��� �yۣ�l��q.;�P�f�#2��S!���&q������!S��u��M���D^+��0����4C�����Q�f�����9Jn��P����Tq�����Q�+��,9���,pT٭vd���Me�T��^�.�<�|$ۇ����b�K2�R[�a�c(�rdK'�@X���6��)y`�B�� H%҆G�`�;��Ha�y��+��
Y۞s�_�� �S [F��j%���o���y�g�����&̱��Ŵ= ��YLe9�ӃL -��{�O�>5���\px9�����9�lQ��ڜ_�:�L"9�^�	|ǟ�M?nΧ7���}��`�`l0(����~W�����G��Ó�Uo��~��K�
���rً]W��2���|�_|
�\�/IB� V�� ��p����;����Y�@��p�bC���K>��q��+�{��pw�������g6��_i�\E��d��]u�,��&�(f��L��X���n4mp,�6Y�8�1���"E�A�}w�y�q;&R{]9ҟ{:�� !�ly������u��U��7�9Ndlz�[	�����l��f�o���5_8]��(�bHW���92m8����*��V�F����4����aZ�+���������wD
���^�EO:�ez*�x3C�uL��}�8ׇ(���������B4���<�<^�:o�t�x��0�9)<�({�y��~7��:������%�?W�>o���b^UP�:� ׿S � x{��;_xGuJ��W�VdN�/;\��ݝ�^4Q�u��E�+�Si>:.p��I�o��6����5g�+L��9�,M�uh�h�
�^Qȣ�v��7�H|�2�����y��c�`Q�F�d��/�\�R���Co�w��,�:�r�n�)��o��K�9q3}�gLYk:�>��1龺��	n�$9:��j�"����;4tC2�=q�����tf�F��`ݹ�ӯ�O���o�w���=��'z)LZ%;[��S/����:VD{L���������U��{�<�e�+�8�ꋯ�����Ro4�F���c�U�ovB̶n��s����3���U����1m4�y���[[�[w#<�,���m��a[f���"a�nw\<���7�W���n_;q�n�Z�k�����|�l3t��XN�<������7�cL.kUVl��1:������֏w&9-\*a��2y]��N4zri�e�ӌ�ޫsy����������GlD������[wf�ۇ���]����t���L����R��8�����û��$�����21ZOv�ݼs��ev��[0�p���\rn�7pTA\nnA߻T�}�] ��(v��e�7���} h+���V���Ac�1a��n��Sb�<m���.��j�ʳ�ShA�^�,>Fa�d챣� $@�x�F�1�v."!�,:�	�FA\T�:(�C�;��[a�8h�S�!$y�Ecmހ�e��"�W����繁�}g���0���{"��� qW=�3�q��X+mŸY�8�z��hg��Y�MM�{s˄s��Q���@iu}K*�ҥ;�۩�Y7��C{IrN�uGu$�fv!c��'r�K�}�
4w���<U����6��"ٚ�G����_�g:�-4;�6K�ȍ*�q.�M� �'#kBIPwƩf�uƎ#��e��Xض�W3����;��˲`!��鎵��2�Sl��Pn�r��}�P�AQ����]5��ԝ0�{x1�벑6�*JNÊ��d�͌S���Q_::����Ik7D#QKq�ܶ�a��3���6{�fw��SLu���*�\����Gw;yd\�Z�^%�'{��0��O�کx.Z�o-R9�&�r�����c�/���r�#H�����T�lي�K�2z�;��9���%�M̾��z�4�l�#��豎�9X�[@�j�k<���#��V��puM���d绱"�Ro�!�	s���+U$/�����f�D4���<�O=���\�=w�:'k�eF�=}:�H�S�����T�w&U��xڄ�d����ޮ�����ՙ��E�����j���M�7�e��]4�L�R�fu��T�4S����'$���B�A�E��4X!��
�N�ǯ��<p���i뇮��\t�]'�T�|��:N=qۦ�tt�q�qۧǊ�^'EW�p���N|�yז��i���b�_�Sc�� �	O��uٮR����v�R��u?\� ���h����r<�x�1��� �&�����u�L�^�F�xza��-���𶣛`��p�E3Tq����Z.�����nժ�?
~~|i���m��}�s����i��DMy�TB���\[*�˔�[*�pã��0�}j�����ضڵ���i�
)����1SA�[�%��Ҵ��|i��<��rJ�b��]�9U4E�N�SI>cD{=��y4�>��il��:um*�}�QQs�"���5P5m��ޅU���|��ӣ��L=g���I���R�ub���`*���h���K� ��a��[il�-Z����8��&�E��;�����\�-[VZ�覝��hv����oV�{����n^-Vƒ*����\��M����h)�X�!�8&(����������S����D��N�=Ty'G''W�D�/e�du^+/���Y�gZ�����b6Y��w#��j��i���B��#��F�Q®��~�"rpB�,�X X!|J�
Y$=�����~�y*��ξ�W�9�#��@v¤U��(\czY��T��|�+��ЃF�F��ޯ߮hh�;�t���P7��y�*�G����c~;�M�Tz�M�̙��ؼݙ���F��"i��?$^|�=~l\y)ά�@<0*�0װ��Q��UN�\d.���\t2ZG��P��CH	������4�_X��zE�P�t{���:�</*.�+��o��W8�/��ǐk\��'yh��X�����"�`���}��L�'ё����$��Y��7�l'�!�����~9�&�����vJ�5j��/ߟ~��̃Z �_h�A�s|��X����S�/\�ڽw�Z�g�&^ߧ��!��c}-%?{�����>�b���ԭ�#�w��_���E[,�lp�b�� ���%��� f�υ��`W"H߫SS�[�'*ls�B?�;0��x@o3T<>˻.m��+|��2�|C�����9~��1i&8��I�y^Z���f�[���4�����3���xr�C���dC�z���z��~��W������ي9r.��ةW>f���"j���=�˫+s�s��y�ʲ$�m(�U�J®U%��Qz����ӆ��[\��k�=��QYAK���g�v	�!�}^�ڿ���0�%�Wt�ϣ��m��y��L�y�ޭzu��=�]�n��T��A��V�� �B���� ��E8P~Q��)d%*"�'� ���  �܍�C��[�o?><�gX�~˹<z�&�0��qM�.��s����4��/��x���q��SXw��ʭ�4k�?[�2�tSPϷ����cl	��2���P%l(y��1��x���)CA�;��=��S�`鬨��!�f�1S����Rcc��@�S�Z@�x�{�:-�����ܤ�7�g��E
��K�0�<�b��?�ৠ�{�XPĤ�Ԗ�M�c]��,���۳R��9�&����}I�0%D`&[� Ӂ�Q��ǯ�
��)�3[������A/�#��R�6#0���T�ûZ皇;2�������F��Lư���7>AoX�]C8Uި3L܃S&���x�@��=p�f ���CAQl�3� �p]�:�0�����G���nN�M[ t,ā��0�`m�3����)��}� $u���9@�kf���o9c�gkş]� �����%�x|�n��������;�~��ƗB���Y�~�9�<|�V�V:�C`7]�ճ��ɯf�7���U�������y��������c�xF?jÉ|sH��ޔN� ����F pܶ�V��z�m�/5�/��U��������t�H)�[	�􀚮�}�V~X�M��[U[�n	(�o�7Dw~��w�B�g�~�\@�K�T��d�W*��J}����+��V�꜓)�*me$�n��L�9^Z��<���}�s:s�z�3���=���ܼ�D��`(�N!	D �����,$��7<���������}�/��<��Hk��� �1`~�E$=�*�~��!b�����_��2�hHM�Uy�Q/H���m��Β��?��$z�"�F��Љ�ÀVjc��b@�дG��?����P5�����b�c��1~��y���Wt8��1��Ե��0ٲ¿K4�p��
�
�kU��]MHgl�Z�be��n��&���;I���2�߇nӸ���J�@��F����~�3�i�����X��}Ňw�����
�R����Z)���`�"�VO ���1c_�m*�i�˫n6��'D
ki�!�µ�H~P��yO�*���\�r롎�8��#d9q�8�/;!�.|25���mғ��2h�>m��2�Ps�n�~��NS�"ª�1hКF�2����s�,m)����p��FĂW�x�8�
b�߁6*�Q��C��t��-����zu>��1�1�6c;������k���;r�����z�°�!��/��ƈ_�����պH��Cq���x���$���\����	��pB�a��Pd�	�\�O���˟��¥˸gKHgfM���9�\�d�8����@�L�D��+ޭOK����V�ȯ.���VWq랂����P�U|C�Fu�OϤ��};OAԻl�bl#"n��`���}G��5Kz�����v�n�-��� ��<�w�����V� ��RB�)"��A*|�\A"�����<=�` ��h]ղ��GkC=����#\d���W�{�DRR�QG$<0��(s�dA���[�����,"��i5��5З�]B�W�te�<�����`n��Y���Q8:���8��G��sd_�G���
��X�Ͱ��o
��@���
�ܫdl����)��������1<��;>�߆R�Ysh�N-sRvN5��|5�fN�O�ۑ� :���N�'w��)�ͼP�=����o\PQS����p����fO������� "λ�|��Ʌ�'�n(��ZU��@�����~A�1���=����Ȟ� p-Q[)��AtM?���D#�6��SCOE��ƕ���8>�k�=R���1-�ܲ0w����T�w�?5�1��� ��ܰ��m�=��gam���vOC.�Y�i�1i�ɕ��n��l���x�H�p�OHB���	���;]=�p[�0�6lc�A�v�W'�m��^���Zư��ui�v-�*#��l��T�7�+����f��H &��8��~�9�k��>�ts%\!4��mdu����O�]��Wǟ���M��|��.FM���bg,���+�W5�L��Y��?��|�!�+��� �	{Հ!k �G� s�GDA.�<͵2=�"1*1'[ɭ-��R�'�7�Ve��#�k�"��.�%l�B��̼�pX��p#ϯ=�λ���H� e�p��K %A�� `��pH�R��Y�����Ͽ{���'����W��V0-��-�?�d<[N.�H����\M��K|��K4���1{o��ņA�"��p�@�ֲG�l��,y��?�W�7��G�><S	��ޭ؎h�/P��v�W"vc���"�L0~�� �������a`V�Ϲ��ڵ��U@�Hc����M��n=r$��0= K��^��@��H�e���/�Sv���7� `;ͨ`�+b�C�1=����A��hh��}�-�EW����ǨC�>� �,��_̚�����M����=�fg��<� ��d�.<qE{|�f,3xn�s���)��=v����=�MV�̠'��%�|H:s�D�+|��g�@���Z��ng��VM���^���tN�|���[�\x1|��8���D��x/��J�>M|���V�� ��Ռ� x�o�h�2�/2�����%�ߍ/���,@���B������P�+�J�(a՝?	.'�dCQ�l��Z�;�f7qw�3��������c��OB�����%��`�� ��s�W��L7��爮7�_[j���.e�'�v:ѦH�����,Z��wz+��m��א��vH�F�b�u����S�1
��O�r�B0��AA�R@A Ozvy�=��nn�u�~�&��rn^P��P�ƻ"DѴ�P�fwc����-�$'�K$%)	J"�",��
��� ��ޮÝO/���S��ۀ!�i�7޻c�_�,b��P������X^�ҐT۸��
J�}��������݀a�0�oj�n�U�����wE3rC�	�U8��կnb�����0��^C�]E�w����>�p�"�:����2co�
�j�q�ڟr�"���d���,��qY��ȼH�ڝ��J̈́���p_ɒ@t��.n�f�%s��vS�C���Fk�3��~αz�����z����o��FFH�ό9���:�o\����6�dj/�����M��:a�1��(=O����_�hI�f���(�TQ~����c�@��( ��@�~���T� 01 s篺H�)��f9�{*Su�2[it��"Ǚ���wc��2`ۃOg1�Mm%��_��ȗ6\{Z�h��<�9H�ou�8W�)+�.׹`�����b)4������g}�	>�9g�$�E�Vvy�B`����ؾT+z
pE�.{�y����;Ov���ׂ���Æ��`#l�35a��<�X3@~�O�Ϟ�
~��M�5���u=�K����@� ���Ks����d�����>�����a����f��N���^�Sk&����v�Ӏꚥ��dz��
7�\U�R��7�:���΋�l����v�Qu�㳵ҩm�O*�v��W1$b�:��D,)k���RE:s�`�X�*�_��3$¤��K"�NBJYJQ#*D�R( q�~=�:;}��L��;6ޟ�@j�z������בx���]�0������w,��P�C/9���U�Ʀ{zc��x���w=>���\�9�c�(��B'fU�\[�h�&oLy��K�-"XW�#/���#?��t
�n1�������x�:����*ײ�����n�#��']A�&��eH����1�>ۜTe�l��XH��@�@}�f���9��/:�X̌�LI�>�E4��qѫS�L����0�[��w,�t���A����j�3���Nv�a���!ǫ�MÇ�R�,löu<Kd����y���A��!Ƨ�t{��ω��W�̇sw����4?�=�ڪD������pr��Ĭ��b讀p:AS;�"e��K�2�S�.{�&�yn�� ������5V7��fX�$~��넢w���>:a��Bo� �\�{X�c�2����YHׄ����9�0W�]� �6^[5vV0��/&���k1�k�K;Y��l�}�ï��C\����@��]����uO1.���9 >�ݻ#�r&"��2�ڎjS��]N���+4�pt�9��ݪb��\�ؖr9gMz	aR]�ø�%h�\�l=��v�ٿY�@Â��k��ֱ�s�V1u{HNt�,Cn��o3)jh�1jɮ����;��o���R��TpH u.	����ua�H)d�K"A�?6����	=5˦���(ϥȁ�+�i;!�y�,+�AOADW>�M�Y��oq����x+|k;�J���������3��qA�g���x7�@!����R�qwVjw��0�335�9���^���(8$�8g�	+�a�gU:� EL��	y�W`K6���4���6��[�DHN�Գ���==?e?v�h.��z�����r��PX��G@�i��ސ��C;�H��S���,b����C��w*���� �9x2����ֆi_���f{f���@�d�`��G��}�/���5��g%X�O��A,��&�zǮy���/�$�01�i�VȄ�X��lN/���ܙ���2k{�3�;�6��!��	�>��,���-�7;{@���B�#����r�2WWI�O���;Q��[����C�vd�<�-9tXٲl����
\r�������à�Y�{��_|t�<�*o�K��T�����V� D������\z�ag`Y�F����,��1�����7��F��c��uE�9�<�J� X�g�W_+_θ3�ȨAyF���.�e�k�=ׯi�Ng����o��tj�m�.C��u٬�_A�:u�k��@�Qaz�!9b�QN'�3B��_e��q0���t%]a���bl���Mpk����z��mu~띌ރQ��y��a���w.u�t}D@����*,H��"B�!K�T�J�$�2��s9=�������c� w�N�_TS�#>�a���2�1'=��vۜ���ʚ��V����E��� ��A�My-�ϗP!tSM�Zh�I�=��M��#ӠgM�ćBϰ�siV�]���È7����U��:@�T�>,V1��?������*μ��y��lk]K樑�=s���5�]���~��yˣ?/��`����d�1�5�K���(l��|�V��<��nk�[pn�N�l��f�{��ː��E/��!����^d䧤�[?}�܀�"o�j��ۂ�����Pf����@1n���UІ�0,�$Ⅸ����hY���+��v��{*�t�+Ox&�KSE�`��X����f����� ��}�a�ug䴌1[�h���!�C�L��ޮ=� ��?	{��rs�8�.�cK��ssPH�e�H���饀�k�[O�١�ڱ���.kUڨ�C�fO��M�c�ʢ�?��)�@�R*�����c"Z�Y�괧���['��&}���wN�^����;6�xK ��]�Q�ϫP_�����;��B�t�������'( ��*�����W�Xyt����/��陊�9�%Qo�+1��:M"&��o#o��c��**z��[p�m��mfM��̺�wlb��\��^�Q�{�lu(��S���o�+���Z�HA�}�V�$�?������lG�0H��� pJ���xx�����l[�7x+��OT�;6?|�?��"X��'(zx�P��V6=�8hkoP99�k�LvEv�6�#���Q�:��L$(�0������Q`|�,<�&%P/��_N�widZ+�۴�34���|(P�.���ky���<��Q,����4�}�	��:㰚���#�O�T�����,���ěҸ�U!�Ļ�y�Os�������}m��J�x���!�ZdLto9�*/[Pˀ�{%��0r����A�{T�l�g!�G6Q��0�p���>$o��O¢���هzh@���ƁR��Q|��\C�c@N��1���
OM�[j7o��w�$�Àd�gV��-�ݻ/&��9���V��@��U��c�B?U����v�'��љ�ƶ4�0jy����6}��!w�V\"�b��Qvl&���!=ϭ��Y�8N.�~?��7���k|��5��>����B�����9/m��[�=�'�G2^��آ�^�cKe8A�2��5k��}�<�5F�o����}���H��W{1p��� {��y�W7H���{'sڮ�c�s�f�w�J^�T��Y��u�J��I��9�e��G�vsgG�<��ӫ�H�t�tx/+/V���7kN:J.���nE���8C���ʗ�!�9�Ed�%nŝݠ�T�dȻ�u��S\��tr��ա�nNݫ �����S�H���gJ=RN}�����љ��P:��qr�Eu�3z/U�n������Ȗ��1��V����{�)r��-'�,�'i`"]�mw&ۘh6:�֚���d�������J�K�)
	��k�{���� ܛol�����ruF�ƺ��ՌlL���V͍5U{�0�L���o"!f7^q����6���#��v2ﲚ��.�{��՛�
U+�;��7��j�	��,֍Ͼ�\�#|8���h�d\y;E"9��{zꅩ8�%�T�Ѭ�݊;j߳�4�{�6F��c.�#���fn�FU�������+y��E)�/6侺ȶ
0uA>��ꝵ$��T7"2ȷ{j;V>��nԁ�U���dr�)%�;DN#F��-4Z��D�׏Qʬ� ����U�0Ε�_b�(!Wk)�K�3quثh0^�ɗ��]�A�.�Ȟ�S�ݜ�q��`��^�vgS����z��2�K
ګ	��c�-��k�0S��HY[C'V�(�X6b�8@��~
��.�h��d@�t�a��׸AcA�1��4%�ׯ���� �"%|����ם�'�1����#��g����n��U7��}s�V6VJ�Ƒ}��}"�n�(��)�o"�c�]k�����wG �CwM8í�G�\h)�:���L�M��U�7/i2N���2�W���N����j��)\�kN�O���H���j92���,ڮ�J��C��i�j��<d�����w6�CkUt�Ӧ���r�_s��y
䃗�����c5ESa�egTВ�L�akz����աR��=�S�nIy��@�<��I9�u���t2a,�K%;�-����y��e٧:T�D����sT�2�U���T�5tܽ���ܼI�.���G�t�>���H3f���{�$%�XzQ�׭��ː<C)��7*SɗyV��j�V�o��c�C���C�s�����0�Y���\8�T�%�B��5cDM�N�O:o=��:�9/(�.w\�	�b�y��VTR���9f���*�p��A)�^�R�ٹ���4Փ���̘��M��GGA��"ݳ�u�;ݻM�N�c'+h9�x�7������<�8<�O|�Ҫ���q�� 0@�,h�c�`P��p�lv�c�;ۛǽ����b;�[�%�:�u㚨����9�(������~ӣ����O�����xp��<Ω��l��15E5W9�W8�Z��F��gƞ��w��^��>I�Na���6��:��	HD4Q�=�8~��᧯�s���Kn��RI�����W"�˅�)�X�S6h�.���A��ya�=��;�lR�4Uc���UmKR[jե�����`z���DU3^�a�Yl,���KQn�ᦚi�=�gu)�Pr�Dg6���YV���xS��h�;aڝ��gK���CU�yb�Z�E��f|`�Z{�
V���8�)
��JOv�b;��4�d�p��}���h__:��&������0^��ԗYw�:���8e#�_�~hIZ�yr�kU>�NSf���b����d�Ie���Pڊw����� ��HR��KR������k����{o�a�>�jO���"6���M��ة������Ok����b�n��-�g���'�~v��v`r&�9#sUyO��g��%_�y�6�p�η*�<^:�-M��ɸ^^�w�ş��ϑI�I�?�=�%�S?����vS��ȾU!���y�>�B�Б��N�xZ��~�0�j�l6;0+�Y�;K�jz,n��:�÷���s*��-�ˉ��B�z��������F�_�ec��@{�+�T[&��H�O@,��a>����}�;�k��-�Y'��2\u�Vū�c[���ƀ]5JS��T*D�0�<��[Ц���-�Wϸ��;	��ul�&~���'�
��g��	!����f���ޞ�9?�Gw,��h���{e���p��5@x/G�N#��eF��[����H������_�րGW:���A�K�U��������X��J/(2ƵD��3� ���j��Xg���w0~`���Q��g�����r�[��n$c�L�8y�t�'e����~0����dqda��[�HP:f��Y�p�׃;���[���3y�GR5�X�v��|�������WZ��t<�`X�)�>ܸ�}�yPN���ɻk������G����1��C({�5٫^�ז���ﯳ�:����,��*�(�B��  pxx`+���7]����� <`��?�ta����덯�K�M�C�j�b�F<��@�Ŷb�qa���ё!�;'�ؖJ�M�� H"�����B�?v@J�f��m�~�Q�aD�6��t�}on��{����;Y��e��S.{�M��m�.�`2\A�	q�N�*��0��Z�%Z����	;��0&`W���_�����
ot�t��l7������uxg�+�n�/}���;wMU�������(��~.-��|k�wO�Љ �b`s@�d<�g��*���.��gcin��^���&���<������z���������<��k����q1�_F��w��Ȏ[�[��~����F��=���m	��	
��Hg,2u�w~m<3f:y���U/�tu����Xd�x[�`=wAnϝ���X�c8���=���m�1v���d�4I����^y���!� ���6�ގk܊c�*�y�e)֜)���A�g�d�K7��bu�B���`�������ua�-�����*xH5�j �ȍ�V���<��G5I����K⳪쪘�����+f�ԕ}��L�Ӓ�<b�!.���Z������6'ަO��,��$/�A�l��e��ؘlR�u���oh�oPV�)�r�x?�_�v�c]>�M;��&hn��T�K�������� ����=x��Ӌ{�\�_:���Q$��$JTOh�,D�$�$R��!JI�Ig�u�3z��d��?:=���N/� ����G~�����}��S�#F����r����?uȝ����c~~�0spG�I�L�g�"���o-�@K��!���:�z��� `A����%�4n_�7b�<�����%P���Q`M~J����� ȶJ�m�ӊ���e�~�csCuo.�����0�1�J�Cϵ]Bs ;��q�h0"A��>�]}�v�c���}K�O�VE0����Lj�ͯH�������Z�O��_"�aC�;c��$����w��a������	�XG*�o˶�JU�\�(E]���gp�ܡ���
)����q/��÷K�P~|X�cv����ڧ��חӫ����^�d8��pNc�[_��E
݋>���Tl����	c�V�庅6��C<vvR�`�1X����;wf�X�aofְ�=P��?�6�w��Hf�f���cj�D�ݻ�˦�3pZ�YZ���Q��nGA3�45�u���'��0��;��O@|(�~ =����vB�̹g�-U�E4Y���]_Y�ך��6�'qTΣ�]⦊ؒK��s%�S4YS{k�q�T�[uAX���ם�A����������IF�uG.��3��*���2O�S;���v�wY3��+�� x���+	��0B�{�`z8���կ������ƫ�a��a�����.�@;��m���?�5�Y�y�<=Zfy������0?�����^�*�^@��-"�izQ�̑�˸:�	�m�mٙ�<�z��X�f׹6��b�G0���8~~O-�V�����1祄^ o�|�t���ݞ�teヰ[o�!٨!���C�$:x����}H�`~B�)�Y7�r �.f��$�TonJ�~�X~��!�_|��[�
�I;���#&ȑ��c'�ݞ��y;�5u�`Iu��hʑ��:�}`�L�	�Dk��"s�4
�~A;���|O:;����}�~g�=�x��g�Iv�@9O` ҺO�E4s�ywΧ���e:m��T�F��ÄL[.{��Z3���s���&����]~ ��w����Â��Rn4��y����ה[�,_r����P�c���?�G3�xj��z���Y!&@��x��{��;'��;��n�!��G��ES�&{g��Å�|��^�g��Nِ^�3Ե*�~V�����C�:���U���#�u��U���%�誉����݋{��W����@z`R���/4��O$�ܘVT}���R�W=�L����:�,���N���V�0�����n�]W0�Q������r��,�)G*p�J�XR��'%�����������s��={ۗ�_߶iD�}�S��Z~oB�����O7��~;�͇�>�7�Cp�-��j+�b��Ә��a��C��0ڋi�0r�&B�I��*9�[�6+,կ��f��H����@�^]�WX�~�8B@ՙQO����pS��|��Do�����~��2��R�̹־l��)帾�G�3���e�~wq�+�g�]��\���{|432,0�1he��8��ݯ^�o;%�j�a���&���9���WC�w�u�ϸ�xp�O>���(ֆ� �c�C�C(6>,f���'���~��B��������:臜�G9N�M��~����gOID�*��%�$���e�00�6,)$�5"1����̲̚�oם�{27���qg�S֨���]�����&�ν�9|�W�T�4=����Τ^:y��=�2�j���%�	P��>*-��);�/Cx�튄�A�8/��{4����@zn�C@��:��#?j��!5x���4�'�/�W�3:xHÎh8רu�ahœP��']^���V���4�������U���q��Zk/�Vfn�M��f�w�m�9CAY�`�ὴ�P�P���C�X�b�εÄ�o[,��j:;��.Vų�,H�k�W:�C�,J���o�;�>�3�ſ��*)d��,)QO��:*?����?}��y��t��S'��� M����KC`�/��o)M�<�:!:���΍�v����^�����,R�N+Ӑ����!���0��?%���iJ^灇�R'7/�AÀ�C�{�*�7��X����*)�O��g�OE�p��;���.C�	U�j��gn�|�7��߈�
��L�i�L���E��#"��K��qJ	�t������l�(����*`C�<R*�
ǿv�'����r���VQx�7�Cw�>i��ؔ�I\!��'������1y�lJuh&��{k˯,_nN�-ٷ����̹��c��wS�ɷQ���t��n���<n��������/��}���Sb�a��;jٶ���F��zr`��s�O3��	��[�k�Gs޾ |b��
��O19y��u����	�;����,t��ޜc\����@���z5�:=�t l��H֘ݐ�;������M�8օ\�����W}�Ec�X]��Ok��A� �1Z�X1��I��ϯ�v��N�-/0�p��h?��{r��}���`eb��wAבr\Yyb���"��0�����sn���
��f�དྷ�6Ժ]%��s�rެ����|�v��V�v�-��!w=sO��o�x����l�V2{�"�c�`���%jە�ƹ��P��`���`��`�!�%�x�����CA�;3{`-��)ܪ.N��Q����P%���Ť'�x��y��^q(���;׀�|��g�>�iy�������������s��'�V@K˖ 2]:� ���/���>/�'�/%��_�[Y�ķ�s�Y��=^�^f�Ju�
)���3�UI��Ҙ0~02�z`��r؞�=s�l0,d}�w��Jm�3>�_*�
G�ѝ����7�n����͐�	���#��c->��@���$v��B��f�Gt�V06��j��� �E~�����	��_[���Ά&l�1���ܱ7�F(^`Xa���Ǆ��/��u���Q� ���ʎcv2!��}�l|�6�ըs��<��ԸϓE�;x@��a�zi �3i	v7��s陳����&��g�[y��_�9�[�y��Å�z6=	��S�+���?A��O~����	GnvS#���381�ͥW������5�N��C��Α�o(6	��j�c���8���&�>>�{*�Ϸ��(Rºgڂ	�a|�T���|e~��V��OaW$3�ؼ��'qnCa1�x)�Ҥ��a���K-����XT4���CҭjǎbA�o}��G�gp�܂� j��l�w��V�jj�f�o�oג��QԬv�~�/��)e,�����IÑΫ��\/������u���a���V��� ��Ĭ�?\(:�u�m�!��h�񒾘��iĄ��j��Q}�:��$�[:�t2� @`�3��/���2�����ފk =�)� w8���G�h��ڹ�ژ�;t���M./x���ۀAO�=(�`3m_V���{_ꀫ#��'�?"q��砊w����ֺ�A���Ҡ3+���;�R��}�>�YCvS��Y��y�S�+��$n]�^�ˀ�an		��v��&(8���<1k��v<�!��P׹�.j�ZsG����0R�1oZ_(�_L��oQ���.bMO�L��nA9GAF�-/�5Q��@�%�2�:b�SU��N��~�z�h@� �Rk�aϾv�mh$�缙/���� �o}`n�����z�=���֣QI��{M�nYo��hl�]��`y��s��q�b��\�8��f�ǱO��Iz�H��JE���ȅR�Y'�L@�(`ż!ݛ`P�a	\ՀAo�X_Z����ɞ��P��դ���Y��&����#YC߉�G��x�`��?����`�1�o��Q�� ��f�-4]�>��u�̺�Y[2����a#J��ւŸ�:��~��e�h[K��m���&�7��#�P�V�{s�����:N�x�9�l��t�S���Gv��YͰ������������䆯�0q��\���p�-,�)e.���0�+i\	S�=�>���9�� �>��/��������+�4����V5s�yw=��؎��o>ok����0׫V]��C��{�z�TJ3�9�3n��S7a���P*���G�y%>���w��P�>a��� ���y�t��
e�4��>���nT��"yk����;�S�0�o��]"�_��I�;��hA��L6݌�0�=l_pnR�)l����!��cݐ�R�Y{լ)�nC��=��:����#� ]cNT�1̢k�̽#�}�3����tݏW�E��wm�}n*�7��BuG�w����l��e��uP���̎����z��3EF6��aH����X���zޱ~���47�._�"-�Z1�i�r�S�:��a�ƷF�	�!�E(���_L���Fd[�u���<����L���)���?N�����z�?��]"l��
:ؼ~5���o��O�0�K�CdCS���8�6�A���?��}_i���{P���@�bc���@M����)�_)j
p�)F�J��F�w5Lh$K���<�J�w/��g���u�X�ǿY��ipz���.N;���r����'�������h�~l(jx�Bxo���b�C���upy��0��kC��>9�]�[��1�S���5g^�IN�9Y��/���)J�RҩiT�=���}��|�<ߡ����=#�}�Ι��ֳ�C	��6z< �wu�pm��ͧ*F'�������,�N/��F��_wJa#��i�D������|畾G�}�L����G>U�w�g���D�8�����Á�1TP�*�M�E}D�V=�������,������Ƭ��0p��s�4ɤGF3c��5�Q��?!�w���ݹ�S{*�l�o�:׀h�?|��<��ߢ4��G���f}��B�V�����c����U����S'F���J��������S�M8���T��(��\��;�`��0V�D\2f��/�23]-���	�:Y���T:5��� 4��H�]�+ք�>{z��c�=Y�2R٣��gep�����Eev��es�����DcG=IÓ�_1��>�����¯=��˶)�z�p��G��sAm1�J���3��\UR,
�Y��݈�S
T��ZO׎�#� ޝ���]��&�����/>�ɦ��غ�
C���_�������(�TĨ����������ڤ�&�5��:�;�s*aŗ����d齎������Q�]k�T�,ڷz�z��k�����SG'�J7p����'�[�E�SY7ijt�|F�{���EM�"�Q��e����E�t�uk��K�V�%Ci��phq�孴��7}���ы��+nԽ���A�S�^�k*���ٛ1��B.��ݔ�p��fZ��p�ֹ����A�����]���C���B��H(�
���{�k�n�/Y̤��o5wj̀�閡[��O�;�ߏnWkT�b�ު�:���.<w�n���y��7����En�4UN�|r�r���k�4r�u�e���-��.���4�se��h<��q]˩�)pZ��^�y�ر)�o�ܣ��sr��Ϋv�&��A&�6���.�oS[j�;xhm�Ǡ�
G��U�-'3oh�{Os��-0����A�.W�*��j����{Pu`��Y����]2^�#�5»T�twr�;s���?��-�n�D����$L���'07˫K�T������N����$��Oq�����=}jB3E�6�ޅ�I�����C,�m��F���R�v\hê)FL���![J��nt��}Xo��2@�JK���ؒ�G��>��
P��,��k��:��`�(��@��s��L�z8ga���"y��ѢXHdt9aa�8����0
�����v������>}l;ŽDOv<�~M�ȸnP�3 �;e�`���-ȨhLPX�B/q�,ꪣ|-�m�vTo��%j&vleP�W-��J����S�}#��U���˫�n�ۛb]Ypcunaŷ;���ry�dخ�L�;���[�2+�y�·uV�up���O�kⷲS�T���ШΎ�a�V*��y�^|��i��&@�Ue�1�"�UBV�٦���@�:(�LD�S�yx��0�\�oJ}�oU��{hl�ٓu��v��ɺO��{}�9s��.�[c��Y�?�@v���mG���K�U��7e���8L�����6+黐N�ۦw�(���c�V8g^ot� ��&ػ�6�TT�4�UEIТ�=�n�k�K)���9�|)uf���v:�vK�9u,B�N
�d.��	�orm�X���E�ɵ��X������]pi��qy�T�[�K�e���̺ܧ�����+����>q��`�yʩ�0>l�9en٤�Ҙ:�XN�������}�N]Z���ٝ�N���<Y���7q���t*J�4���}��S��=��V4ݜz��r��o7�)��)�!��Vnf��ewc���ts\�r������M�i�%���ٽ���� �A�, 0!��Ҽz�W��8����]�t������=z�N+�n��Z��OU^+���8�ӷ'o^�x���_U�������u��uOW��%Ҵ�$J*ZT-��u��`�5#�E�F�O$�/����g�X�kT%4u��A���O�>����Z-�d�ݣ��MR��HҜ1��i���[b�lr�,r��(�;���z)ã=a�;CI�%^6��H��WI�'�5H�h"B��A��{>>0����Y�r�j[�NT
��*�)����x�X �采��'Ԗ�je��Ų�Ô�'*-�ʒ�e8va�a������[ai*�jK�"�Y'V���4�M0�4�=Hw\���^�=A����'p���et''͠���v����r�%4|�RP��:�x�(4|��+��
�L� �r:��{�ַ\M�(U���zϑu	� �5+6�t���tPM#,�y��̣:�����,��+�Eb����;�u�r��>�wo,��r��4��@`C��П��-rp�-+�x+�[��>�>�|)��@����n�����|�_�(���� ��W�u~+�A���o��������6��R��y���57���#��;���[ORD������;�����_q�����B~a�́�,s�۾���ƽ�ʭ������m��C���F���=�����r�7��,��X��w.>����5˿�����otv9c?0�����7�_��g�8�Ts���SX����nKQ�i����]�S��ѩ�:�n�b�����5�Q0���iD�YD��=
����b��Uj�)��DD�m��c"ԉi�%��.���,{c#�v4��a�C����\��zޙs�Hf�����Y�'�"c���A~l���6Ů
�jr��-�*4t����S��X�@��Q@�-�}�t1�0ν���8t���by��1�1���l{��&ߖ(�[�� ;k�����
�W}~��bY�B�{TO�����q��������>y�X�1�gHږf(喾�n�������~��3!�&�!������sA��,}o��{�;����G�ʄ(f	SteR�J�+)��Gdh�ҕq`�Ev��ڟb�6V�t�|R�:�_kaP۠�,���$�z�͏�����E]Ҫ��f��u�"�t����U@ݛ�,�-��m���|z�߾�tlk�򾡆	�b�,r�>�+��a��{?.��H��j(Ȁ�@��	��81iP���Q��r�i�&r|���o��VOZ��_WKw�cM���.���@��A���1�V�@&���vmL*�i�U=�p�RX��k��`SxLlohcm���ϰ��C����`Z~߉u�� �-r���:	L��Taݨ�ޘ���L?jF�����ֈ��T[}���
1,��Mu�|�w��Ӥ^l�bw����ViV�Ϛ��J��1��rD��q\�[+ l�x�CvSHԋ��ilGv{�X���^���e"�����V��5i���Tl�~�	��	�d��fn_�sc<e�iv��a���a��6T����F�Ee)�5�� mE����O���ٖX�!�]��m�-�����_@hV@|�}&��1���uϻ��X��dG\�i;bBx��T��sQ-<�6�i�{!k��-"G��3��4��g�H1 s��K?�tp�عe	9�(ent<�K��Ù�-��!0L|�	ϓ }��_�!���ȃ7\����sjFO?
��&U4���7�fCNO*N�hcW��c�gY���8tLr�*���s.�L1
�ן���ƨ��}[[�8P��,a��]��\��$f��ir���1�V.�p^��D�o�]g�7cU[�b�L9���ğ\��c��Wc*��p���)�~?�/� �,�)�NNrp���~f}�����v}��qh��v��|�l$i�/R��9h�R*��%�U�6>�j�O��!�Ŗ9&=\�KHYo�����5�K:�NСP7�XǮr����^�fΓ|����f��8n���oک�Ȟ�*���D,$N�H�Ϡ4f��S�7��$/.W�=�#pp�<i��/�l���zO<�G�I9�ġ���>iJ��Sm1��=�l�|%�Le�H~eq��G�=5ݼ��И��G��3������/9f]ԟ���`�%
����5�ڲ`�(].�'�cu�$	,�o�+�Ե�}�s
�C	Tk�{�%�s�w�jj�_�X��2�� 6P.X:0���Ϥ�}�O+y������C_%@��z�SPb���p�*����QJ	y �CK
��x���]�5O�-��c��������j��Z����)�Ccf3�}�zSXx��a��0�ڍӽ�»ƢE52c�Z�o���]hVg�����5��S�c�xpW�}�jI��V�^gr��n�ы�r�2Q��ޏ����¬��V6���p�Ŧ�+`�c[�zww�<�%WyU5a��D�r�-���:Zu���}�ў�oS�uw��'^$��e�(7��כ�}/�?��-)C�s?w�>�?^Wa�[�C�8-��'�-����BO�O�+��� �A�;�����[���3��W��l���n��X�y�QM���wO��P�vF��;��F��U�PT0�z�ΠuD�D�P5�Ֆ>D�1@t>���������5��^�)���Gce���=L�y5����ڂ�qgז���G�c;K~S�|�gp�[�lC��*��8ɸ,8w�H���S	�md��a�C�f�x�Tظ�p9�F�0�O9;M<0���zM�׳�w@���!���Ʊ�	�����q^D��uA^ �v���cw;���F8��3�B^X�d��r�lcVE���1�cjzb؝�i�]�g��̡�D����t��>���n��/�0P���6�x5xcY�̨p�]���L�7�o�7��yx���f @ǉ�H�����U�����q�W��|�-�Y��ӈt_L=��͞�<5��za��9S��U���c ��r}3�P�c��~�qP�c$E~����}n���b���7ou���.v[6�D遑�JX&e�p����(�i��+	��D6x�rܹ�l�Iň����XѶ��($u��7HF*�f�|��ޔ�㼷��N�8�o����O������WL1������� ���� ���ȡe�� > H@�ӄ$��޷ݴ��r�Y�� ��(�.iję��!X��P�/"�C��x�8O�K�v�c\ {��؀n��u$d��� ��0��vS�-����P����[�ު����<0��T�F�gd&D��X�`q\mNT��b��}����g�k���?�f;$Kn�|Ǿ��M��`�3�V�}�*�������:�培�DUUb���6��p���	
,P^5�c�"�~���,r�U2hN��{���*��&���a��.[�:��q��[���}��B���5sh֭���ʭ�������u�ʚm�m�X����ڃ[P@SP����p�V��TH'��P66�i31M���/{�AOJ$	�}l�m����z�#��<�ݰĘ:O�ٴ?#>ft|%A ��w�+Y�xVN��"�*@��zu˭ԍ��{<g��Wr�Ϟ�A���@=)�c��^}�-xLߛh���-�[P%��e50��=Ѱ���P v�H��4_K*��}����$Se�����E��ʷ>��h�ʯƸ鑥y���f�q=��P�1U����	pX=�($ݗr�u�z���:ss����N�tW��ȏ]��3n�H������_l�kF(s�F�T�%����0�}�lwd��%y�-�����U�)��B(t�t���o����c��&�Fg�V�&z���$JvT�	��\sʱW�{0b�����}}e�n񭃉�;���D*��y�b��"&
8���F�� �9��]X���t\�E����⚙�k�Gd*��64/UXha~1ڨ<3d7@v�7%��:˝�͝�]=�c�G�B���6,��g^�!㌡�}�|�)�7坮�A�igԡ��d����ȓӚz���^ۢc:�O�@��h���X�O��_��-�c�)�C� �;%œ}_p@�Hp3��b|�� �@Mǆ@]\��E���otzj�g*2|	D� Zo[6�_�D��a���D�E��P���?[n�B�h*�*s�U�Y/N:k��7�Ēx��cc_���vA/��gH9��_������'�Uth�4���yT>T%��\f�K��~���:�o��1��N44�C���N����<1ڝ����+��E?^}�E��	��w�6�.&�i���i��U��_]���f�k�7��W:�_7]T���V{�|��hP�ڭq�W��f�&�5cd���i}wT�b0�[X� }����LW	�8��,b�C\y�{�'�X�F�	�> @�>�x��������PXF�E�HA_\�����~Ρ{WՄi��#�^��B��N%��J��(g������O�y�%Hf��j��
"��p�i�Z��6	�ή���es���i�����ք�	~j���x{��JǬ)�.�?�t?��.cHl�|Ѻ˾^����>hRL5da�[)���*�As}��F4������,��f�U9k��X��fm|�O�;����.��XLl���򨧗�P����c�iO0���:�4f�լ3���*�l�u�N0cV�M�z�u��$:�o�./�H\��bH�ѽ�-od<�ӝBE\���5��*���EX
��:XH�eW$����@^>�d�^���� z��}�:F�<{VX�uO'cX*�LȈ/`k�3b�W�/0]5�������p�:=zC�u�5�
�ۊ)��9O$�=���6�^���WSv���]m���.�h���"%���,|�`_�SE���Byq&/o�Q}���ò�UFX��m⾋D��S���)��%�,�ne�a]Z�s9ջ�� o��:�\�vx.J�,婛�v�!y�j�{�d�uG��;8�//���.�B�[�c�������-vbn�קS�Y�0g��� �3꽜]�#����c2��?�Ғ��s�w�?�:J+����T��e7b`죃�?|��|N�����{ןB�ݏA�~a���LiA�KHAѬI��dy�����7�`1�O'/n79�qp��7��[,`qB":�p
�Y�|��%2��P��z�����%��ơ�e���4]7NgJcM>G��k�u��� r� QW_t��_W���^hT�1���P�hF�=j�zc�|1|U(��oU����'��5=�7�k��2!'�=`W�-�Y��� ���^q��ת�UҶ����,]ķ=��]8��͹ph�f��Z�y��m��޽��ABv,�C�}���B
�Z�>C�O�+?��� ��w�������6t�sՏ�$��Wj�{Z����eà�����P�醆�zǟpe�[�M���)��9�2���w�O3Swü_S�!GN0���e��KK���gO���htL �w��_w
�afJ�m�����j�P��S�럓PXv5F7������~+�Z��3�,�����t��N�fa��1��N���/���͘G1��9���͕ȴ����&��lQ(K�E�x�o�C,W�.ݛT�ו�Į���Ȼ��N���ս��u>2����8�ܧ1ڰ�v��Պb�gyoq���`X(P�E���e�ﾯ~s�;���)ꊢ�j����¼�,̩�7���f-=K��>!��7X�5dTR��;���g�|/��?\�/w�9<-��q�}�
?�0�ߪ����A	t���]����Lg[��l���.&��U�L�7�oj�����.�8��kb?+"
�_�$(��}�-ֆ`�;������H�*C�Q3�Z��V�A�����U�W����*��⦗h�}��Μ���Ɠ<̥��Ã������XCW(:5�Re��!��%��K��n�+3'�9J���xT�(�pb�C�{�C��b� �W�"F"頯�z�Ǝz�N@w����fn��ڰ���}uo��5S����B這a7T6:8�7�C�0$�k�cY=��;�[&�65��	j�`��+Ź���ȭ�d�*������Pv��ӠKV�pK*!�[�"��o~J����~Y1c��K�*O���'�e[j�SS�h�šv��پ,m�ڡ�޺�=�U�>ZA~�TM����r-l��iy��.�3���hz~�u�]{չ�&*y��O*��-��c���Yֲ�r:�&�>C���!�v�˛F��8�1�E1Bm���j���OujN}7�^X��,;��+�����J��18.�������T'Gk$�����#͜`�����6��E�ykz+_�Z�u̖�����Fm�*�h?�O} �g�h4z{��_9�OηN���Y�����=@ALMѬ��������X���n.'m��Z�ǫL��s\��Z@n�L@�-���}Y%�e)��S���e��F�;}"����9b�u��ގ��_]�~�Bv�&����LTƁ.�fC�/"�d��qˡs�=��`"�/��V��!���+h�nM���C@�� 	�ޝ�qN_C��0�ϟ͕q�zYV!�9P�x��0x�{�:��k\n	Ȃ5�c[�(��E�<�ϖ�ŷl�>S�y_v�B��9����	����<G��+$B�U�&�����wlxu	��q����2��Y=��ލC��������cc�XV�$Q��%���^��8�?1�5o�������r��qKC=��n��{���X���\�s����t��Q5/]�� P����P�t���{�������ݙ����ʐ��zx1N��n�x�}����[����GTFd��i�(������U����`�]f,NX�Cu�׏q��9SƯ��f��/E�c��i
�����U"}���Ɇ��˱�uy�Dw�+X�l��˰c�Vz�r�Kk��Z��C��2q,�L�������{q��n,��)�3�,���U��C��9�9���k�f��9�Դ='x�ۈ�n�G{�y��#���,�}X�M��btk���&Kh�՞K��GK&��.k�.�T�������.��r�r�VgJZ[4��T2�Gw!	�U�FLqS�����	ӂ_[���K��8F����f�6/+�b�����P��ij��8��U�G �U�|Q9*�,���J�c�gmsYѫ] �\�%JT��Si�
�Nrͻ�U�u_g7���V(8�fL���k�41��*��ē����XMWہT��m�;�(Z��<��̰�kB}J��B��Z�W���1�����6�74<�v;U���
��A6���JS�

�gb�3���jUfA�ڊn
n��d,
��IB��P�E���IT��3{5櫖�ֻ�֤��֙���"�ʷ(��n��f����L�-8uo:����%�Q�H���U�9�a����Z��Ҵ%�:Ъc��)�!�haQ�T5���X��gp�l"	����A���0h�U�>���
�*Y�b��|�S��Sz4i`��x��8��%�÷0/
��� �#�0 �!�%�;C� ��o��$
�Ew笏���z��Fo�&��-�]��Σ�k��捔ˣ�̜�T����pt�����ʌM�n�71�2��Utr7ԷPf�7�]=�0WT��T����Wqah_!�LTԗ[U��g����+^��Y����u4����c�*	�j{�����`�-�2�n:4���1ņG-��S�.X��;[���h��O��YƝ�m�l�f#�X"�Eݭ[���2��,U�Yևf:���:HZ�۸5�U��s�3�����T���n#�t��TY<�<-�j3�Ó�ӊ�����u7K�t�j�7��J�����BrI1�mܫn�e�^~[����5|'oq؍ �UJ�c�����Uތ-������OQn�<:}�c�÷�v�9"��^f�ʮ�&eKa���M;�Cs��I��u2�/{r���1h��CDz���Z����{K_'���|�ɤr��U"]M�+f`V͕չ�x��ob�_��J[`�e+B�u����.�JTK���\-_VM<�pp{��蚺�;k&�;�a�Yؓ">��j����7��sA^]o��Gӻ��,hCF �C,@��Â��vЕ�a[ӻEJ�{���{ ��y/�/&���rJe��il�i�}|)ن��a��}8j�����Z�gU��d�:)�M4����;�R�����7��HR����Ɵ|}I�(���A��9��.��4����L��O�>=>4��}KVh��	�|K�u)�WO 6��wg��<0��0��!�=H�}C�Ĝ�H�JYh��p�G�i���M�_pP�d��`�S��:)�N�0�N��=I�M��>G������r�I�Q�N���<?����>C�>�S�:�(��d<�buS�8EJ�J]�:�AH��D�{O{���oW�w���۽����2�Η��Ф���_u�x��ke˜���:��u8���a���q�� @�ng�C��Z�����]�ĵz.9`��=v��|S�0�,3x<xԦd�;]��/�w��	�j�	e�+�s���I_ʃV[g�����m���ݗ�P�Ⱥ�'n��)�f�;��gXmn��4Żτ�.��(�z��OM�#3�6nϮ k�_1��V`���h��<��;/ۧA�����}�����R~�C:�����{��-� ��~�����Ս��bԍ���VQ�I��aٞ�� >���]�(GB/@.�c�3� �h�A��w蚪��˭����􆚞��Pk��8}F}!�3pW2���3�]խv��)=s��X��ek�Q��@s%>��_��Y'���:o�\�<��>V���}�~������1��!�ff��tj�8�����aj	+��_�dܙ�߻ ����ŋ<oKҔv���{�����ginJ ,Yv:�v3�e�c0����Gtiz����������츎���7e�2Xe\cxzY���Ie�����]����p`���ƼO��,|�U�%��0|#6��V�$�E�y��C2��Ɋ��jrR,��ږ�g��c����O�;-���j�:��κ'1i��E�o,�tE�nrBҌ��탚A�K7����U���B�C����ƀ;����g���,�zޱ���7\�R[�A�����UkH	Ex7�j�N���ݛ"�$�t`�zW�7�����$H������*Ρ�زF��$ư`���'�^��3=3��q�1�V����!
�I�?�F��u}�`a�=�i�C��2�����m)^g\�K���v6n�.�mh�' �o-�yD���� �g@���'��A~7Zc����C�S�[�=�7N"|�.����bA7���_Y��iFiߨ�j�#3�9�ߠ������5K�>��_)�)���r؛uX	���l�����K��K��!���� 2�����%�c�S,�c��1��8�>4�f*?b�|Ԯ�O{���ik�Ț��)��f���R���~t��Vo�������%��{aׯZi�z��N�\�4�d��e�?oy�i��6�d�N��j�	�;v�F7����r\zS�h��-##dHȄ�,��2������;CV,���:���\K�J�%���4<���44G���k�'~6>�>>D%ë��a�[o�+����nᠣ��ʹ+Y����j�����z6�VC�B
���;U.K�0�;j�h��"�P��v��"����wU���<���i���jL���͸+x�ɛ�n�θ�F�w���4��4%�A{xH�X!�!�A�f�b�X�.m��Ԃ������,�������UxՕ���������a�ڨ���b��;�h�j^L	:�f⊉�a�1m���sqd��]=�*:CO�b��������7 ��:�ׇ,�˾���݇�����)ƚ��Q���Ia���s��a!d��Y����g�>�z9f����"���X�b�������U�)�����t�;�0�cTc/�f:�ˈe(�W�s��6 G}`��i��0Sץ�Dd��r�r��g?�y�u�4Ξ��K�g# r����@�ܝ�p�;�Z�� ��=���%1�1���d�ua���gO7;�鲁~���_'��a����H�V�@�a�n|a>�lk�����=��*�l����Z��ס�7(M��-/����������A��ȧt{�O�C�ĎVf�]�o�3R���|9Y�ߖ�\^�c���c}(�*�֨�9� ��o�u�|�lY׵��NE�@��\`?/<�P�d�mx��2.� �f{�f+��]u��g�r0����Y^ޔ3��ue��JW�,�U���O|\����ׇDˏ��Ũ������y�$�����9h��*���m��(Qvn!��|�pm�W(�2��F����_c�t��-�\���\��wp�Ê�ƒ��ll[� ksCh�TSr�d��`&KjDۭZ���m�V�+�Q�v����Ra���?�	�M�ޚh�5�{���2��j�v/�,�YP�U���-{x�����}۬66(�)Jg��*uAPܦ�O��Sx�;���atݗ����U�K�y��ZfX��QM��r�0/��]ǟUH��@�Ƒo������kQ�l���!�_�YP�A���y�
��'=�VƇa�b����hw�ߺ=��M3'�� �%��9�[�p82���|Pɽ�8=\��9Am]�X�=�����E��hA�1��YnRp0�3�7��v� �M�`-ݺ뤷��yP�����F��u#u��صE^���u���Ϗc�����P��7��9y�B�b��ޘj���;���Ό�&]��躚�����p�j�@�`�4l?>�e���Ζ��V����ɫj�G%�uFu�Ú��Oc-�>f�1�{�R0a��1�Li�~�P6s�~�|���^qΌF3�[Q�����%���K�U+z�Л ��o)�;]4X1����.�����Wx�9wX��T"#I�_�s&��1�y���׽����E�+Cx&�*9��0�0�T��s1�E(7źm��8S�	�Wi��ڬ����!�7�<� wp80xp�=Z��up�hsO?�U��|�z�r^�w,'�_H�Nn�{�'�T9*n��L>RB�w��]oG�z>��r�H�l�����SΝ���s��pD[F�T?8NK�ޙD�Z�*�w�x;>Lkt�+��:�}j�[ DCzi�h@2��8\W�T�>�=�w{o�b��m^�mg_�->I��}��˘
�v{�����F�ރ�ߟ��y�,�|�cjg��Jɹ���(0��+_^��p�N�V��!G��*��� q��G�C3�N%�(+��(�3w��K�N����$��ҿ*�Ֆ����aW05=˅��nb&���5��wk��o�Ss�s ͭA<1eIeS%�"tgN4�~�Y��`�hN^�{�
��>V�Ɏ�����{L��6����S�{:E6��ǻ]9&���h�[ymxϳ3�����8~���`|���/�u��+^�G2Y�+6�Ռ5�\\�^��ΰƕ�x��q{CK����e�k4V�f��j��<���>�t��� \���.]������J=�2�Ru��ܗ�W^:�镡E��뎰ż0C�c�;z;ȞWk9�L:�HD�㴆�B�����&b��)/rY���d��/��/9[ՠ�gfJq��]-!��b��i=xtGml˹��i�ˣ��P'�X����Ѽ�����}�w}���"��8�m��M�o�"�q�[�=ve�E��;1��@�b*���vfvq���2�ˇ.Z���zk�|a�#�p6G<qz���P�_���1�`����Xg�TV�243c���|d�,���vG5bC�_䬇������<�zඳ
�R�7��cJ�e0`2����g�}�q�:��kЀI1��M�`����9����-�ov����-�\ftX�='�j���n1��l�T%V�O�S�h����a7�\��Wa=��̺���L���/FD�|��J}�A�=� �B�ܼ��1����*z�˦g����y��9�<)cC�@�D�ҁ�� ��}��|~�1����k�;9Ew��e�8�\��ޙW����o0�&"Zj���=}@��|� �n�MQ�-�'�n�����3Z4�X:d��=Y�.8[�f����%RɚwG��ڣ}��v��\�%��[i�@������"�0�#�e�=����l�	��9�����k�1�+���P�8��7����=R���uI��L�$��\�t��a�����m�-�Ş��2d�>�-Q~�V��t[#�9�-�˝�>h����ky��0*���C_T�O��]ŭ�S�Saz�Xj�ٱ>ȌD�O�U�]�s��/�	���[���n)Z�_0�J��N<z�A ����d*�B�FfTş �� /� >O9b��j߮tA��t@����䪔�^	�vg���S��� �U �v7�XSP��xy¡��C+L�3=LV_=��k�co3濼ϐ&�.|`lk���N���޿�Ӭմ.�������0yDL��$���ه�������}�/�U�4�k��q���O�$�l�JΠ�B�֑�I���P�$X�s�-��@ff�+� /��>��@�^`��?v�X�v�̶r�U�vU��QM��O��]�J�yhuj�/=�ИD��J,�?�gW�vKA��<0!n�����~�8�A�����9���Xs�\H��hgǒ����:��U<q�w<�X�j�؞�n�2&���F�Ҭ�e���d]���$<�'b��S��kr������)���l�dG8w|N����P��S����C�	q��,q#��u�
�Ȇ#��,���F�H"C3��q��3�hs��LƧ�o<�dl�{:�� 1E�B���'�
ӈ��{�l�(���Qm�Ə2>Li`+�
Zo��	��f�<�{�p�6E>�g-�5ɲ�nt+kbE�I����s�q��ʛ�Y�]5��\7�s�A(�$4����׆	A�C�[�'ِ�Pٵ�[t6N�t���2g:���l6����%g�թ�&�4�߀�� q� ��gp��d�]q�����ք�\YR$�	�$N*}��M�d����aY�gsk���4�/x<�L��Z��������n0 C'L���Ѯ֘���#���W��v�V�]��}����2f1p8�i�N�Q���zym��m�e�Ȝ�Z�!��nLM�����V��� �^с���Zeڊ�p�/4�r��w���r��i��@D�j����5UG��h3��)Y9:�O�v�"�Rf�ͦ*n��w�j��f��%-���� Y�h�ۆ�tqi��]��a7s�;�TΟ9����|�����Y��m�.�+N����pPNW�Ou�YU\�^D�7�ޡ���Ur��sE�V^��C���Y��.(ױF��agP�\Oq���6BT��og�=�*�)��/�I���C�����w�Xg_k������ܠ(���E]�����s��Hv��Z�����hG���������t��]� {H�\����E���K�²�r�Ugd�$��XkF��J2��Ƨ=�ʊ��ۓ���$cu<֊����9]uAN��Rs�WyV���_'�F���?�>`x �!���XW�].��t���q/��25�=0����b�r���wΒ,]\,��pC�uh�>_��s�Yܘ�0�p�L���S3�ݛ'�P
��[q�n�m���#o�6�r+9�wݭ�X��T�2�RZ�rK�����V��m˫ݞy�a&���>�6��]��6��5Y�z{���ɫ��m>�{����g �E�3�v~��\p�G	��f7�l��Lp�T��h����ha����:^����j�v�vSZ�z�<��3��Q$�MZǄn���pd+�Z��۬Gj��)l���� �����r�
�se�PG0];���F�8��o �n��k��ڱ��
�mۆ�n�$!�x�]4#�ʘ��[�*k�sM�i�+z#osq����?�;y��m��;�2֧�$M�ry�Z%ݼ`s-K�n���O|��Iw|�v�X#��(TH�u���uͬ�}���q�⢙����&���]��@r���f��
�1@
&ލiv܈���Js%���Z��t#��wƴ��JY�B�6f.�.�L�8aݻ��z����?�� 	 S�; ��7��itO\ >	TC�iOP
���F�TEu;Ơ�W;{vCE��#sF>MU�B��q\����
�f����;�{�V�!��"񷃙S�.C����Y0�{Z�@�����m�90)[�gaP4]}ݱq�o
L��;.ooc�{⛄������l
!�Z��G�,�⧷hخꜬl�x��e���Q�{Q�� �#+ж<�a���(��=kc��8���R�FL��k֢�W �ǎҲC�x������[�ggi�^��f�4z�p�$Nf�����dl`}v������w�S�(��.^���2��#Q��үv�*�l
�����38�wǧ�����z��k�d�P�lv���������o�d�eՁRvR��֚�F����GF>�!A���@LjmwHû!�� �,��&��`{��C��vS�0b����p�f��[A���$�J�v2lx�
bs�t��rT�b��1��Q͗nErZ�r�ȍ�s���3h��UW����T���vj��ܶ;��UvF���D�ژUQ���^=����x��0���.�c�t*�K�Z�ou��W\�P,Y�m"�k��ru��J��ǩ;{u�w\�y]��o���*��ߊ7@�C���ce(�v�t��/=Z�e�̓�U����e�n����OM��Bjs��4h�Y��hAv�F��S0�Z&#��V;��-�Y6]<��<�'2��[(��¹�C���s�b=8cNW#&+��z�ǘI�ؘ19�}��tM��Р�w�OUlw��G���mu�ֻ��{G8�43k�-��'p�\�&�ی1�7�ݡ��t�hy�5�S��Q�i��6�s���Ff3y6Q�ڹ��8�u�v�P�c�b{,�by�S��Ԫ���eZ�FVc�B	YS�6,��1IF��c�@��*�eA��oq�d�E���Z&d�Y�\ZF+ye�o`�ӪS�$�]�t���i�l�(tѤ[��w����ު��<������`�p;윲��j���i��a�q����vz'���3y8Rh��ʴE���9��T۹��z�k�k�n;�W{�ܻq\�d>���< �#�ע��H�����f_/�Eﳟ�o7���F ���u�(QL�-�%=}�P�G�,P��(1w�C{�K�ᣋbPc[�Ì�#�ޱ�w*R����g�!�4�f�d`�5h��`K|ɟ=RI�-��S���w)Gָ9��gݻ���Ǻ�WPt��3mF���ݾ2�!pS<��4R��)pqM�_VAq`cmQ�N�͹��M^KY2�cNe�Qk�Q�,M�u.sc�.�]e5gqY׏��Zir�J�W��n�ܾ��#lod���K)-\�|���7I�iZ��}�KΧr�-�9�Mӵ��T��4'GN��bF𹚱p��}u�^��c��:YZq��G�������ҵ�	�\��_N=gSp�&Uu�TaE�z���dwM����t�F��XR:��[q��[,��4�u�,�J��L��]u��QoE��X��n����6�w�3w^��Ů����ܲ�r�|�%�^�r�~���R��:�gm*���UuW�MIڨ�����.&���K���0�����c��vJ��
9C#�S�
�W�N�5r��p��!��F̴l�n��ڏ{��8u-6�GWw��[nnG����m�(��l���u@�j'�O���\f�s�����z:pֿ��w��T�+W�~�#L)'�Dw�îg7xY�1��8 �U��.�S�6=���((h��Z�:qۊ��;c�x�;z��㉏:c����\z�]�|�:Uq뎞�:k�:U1��8�]<qҺv�O�x�]1ۅXA�, m��:��B���LX�²�z��r��,l9I�E5D�R�,�{��UB �R꣤�T����� ҞetP��4#��r�J�S������O��2��_�&��<B�B��+�_ķ���p�M4�����z� Ҝ�����	ԣ�<G]j�Jp�M4�O��}KfXy*�Oru'$
����{0�O~���NXuS�?(�������u�4��y-	g��i�}	�$˕9V�}dՈꤪ�܇E:4���>O���=��	���)��G$+^A�(;�� �<;4��O�X��#�R6�u�P=�r��P�ҾetR`��ᦟnH��;�jK[m����=�k��4P&�i�.�9)���J�=����ּ�Xe�S��]��t3����+h�ܧ���>]G�Z�Um�s��6*�ɤ7����6	}�����81��`��c�W���u=����X��s��@
@@(���}0�X�J6��	>(,�/�C;���y}������d @8�J�1R]���,�d��N�	�c��sd�����\�=��7�`�����9��'��2��H�Z�B�V#��g>o2I����:�|�֘�ܐ�%�5��&yvځ~־m�������4��kL�Gov㫫)d��L�e�Ģ��l2��&��	�!<zl�Jb�:���k��w���uu{Q��{0��j0�z]�3K�uS KCΣ��{)Z�h��[fzh�F�ӆ�Pӏ�x�4�/[ג糰_���<���D�\�0�o`�����O���^`c�9� �U��su��tG�'K^w�(OG�~w~�{���H�q��^�#y����W��4�mz�O�H��o�" �Y���1�;�cd��oEj�F����ֹ��Y�В̾�rί{g������֟E��.n��o)w����6�@��NY�t�Ȉ�̑���aY�:֬��͉	ܴ�:}�Y�S�Y�0\{$��w!bd���c�8�Ū���8ހooe��E�J��N9F�I��R�j
��]I���~ �<A��H�8����WV�P�����@J�����g'ȣ+�<� ���kw	t��70ūUf�Y��|��oG`�NM���*�s��ggw@���F3P��{��ޜ��" �7��5�x@�l�r�#�=k��:��F�v67��%�-$Z8F+�{L>;��3�.Eʀ�~YY05e^Nk>ֽ��p:����) �kZc��tb:�>`~����&�֖�+RG�f���sz0k{��!<�v�!�Kq}�<�Uٍ��.�Y�Q�� �Iuw��0y��� �{��J��W��i��u&Wո�̔Ը��^$�Z����j�e�r&�P�0(7[x�L��݉��a���L�	�5�;�I�?x(c����� Sڧ&H���A�f��K�3��צ��o�W�x�]�+,Ӿ�W�T
�L<�5�YVc���j���gP]⟥���G#z��Z��P�9���]��Rn{w����m���|?w�U��O=��w�f�"��t3P�.�+d.-nFV	��:6��uk�ɝϫ�\�E�*q3S��9���}XqwmV2��vŽz�'��p> P `?ӥwun��|?i���̭�l����Q�5nƫ�A�H����MD�<ѹk_:FB���WE������/ ��ͪmO,�}�r�n�<B�:R6��k�����ݳ�{������j��r��wݤ�ؔ7�M�1���]�]�Y���եJ+��w�����n'���C�{��=�0N/�lߍ�T,��5���*(��{��󞊴�ޕ
�l�]���	촁v݆�O����9Q��B{���:rZ�r�<��oH�4����"������j��f �4���mB#yL�<�h�y�ɍ'+�볓�Ji�����<��
i�$�_�9m(�}��8�k���h8�AڋA�)ʼ�X� /�䯹|C�F���?3_�Qͽx{�H��.��<9�^��!�U�t`k�uAgQ��x���FT><;��w��Δ����^
�6��grk����pt\��	�{�����Ҹ��qDhf�]Pl<r��F1Zk��᣾�>s�(�W+��U�e��I�]���e�i$ksz�0R/ך�}|���0��VN(��%�g�k;�����B\�7���� o9b+FE��jћ��7��f�F[:@v�́�\�e\^����Ƣf�U���Q�,b����C�{���, �!��]����'���x"오�Q(z��a㑲���x7����.�x	���icѫ셚�������Q�{%�n�=�e*F�\g�;!�
��#�^3o>L�I�[E��8ϙ�D)����3��s{m���]f��s>]nэ	��b4j�$��n�V���kvv�s{��j�iJX`R|� Le�b:ʫ@�_�~L����r\xW��ߩ�Xh(1���'��y�ݺ��+�i�"t�Yۍڷ���w�;!����NF��K���1��kB�'L�QGP��[�r����5�<���$(��M��~U����h�U���]��mbw��v\i��vu�6�yƍ���w�|��iQ����@�1?@sT���v��՜�;n�n����Z��c�nb�u"�ָ8uɕ�������B|��M���"�5Є,P�W�Ξ�x�|�~ym��|	ii/�⭭D�����8Ѿ����zh�ڞ�:��=���`f�1�gtu�}Ƨ��7���q��wӭ�o4�{�k��үv�r�+��['�4���jk�^�_N�z��3�y�=;�Knz���@6ⳬ�^ST<���{��=}�L2���dU�9�mV��y�k��y�n�yM�S*�12}[��p�����2́BB�f+��9qQ��UMk��ܦ�I� $�?Jz�����]�+=2�Y�$/��͠)j�]`�6ϋ��acu�*B�: �j���	Mn_Y�P�|���Q9�.���jg��r� �j���X���k@��^Yt�+O���Y4z���f��ڼ�W.�_^#nE��MD'�-D�V��3��' ��]�K�^�� L���i���a�ԥ�G�J9B��RqƶZ��)+ܻ�?ֳ�~b��Is
�� �����G}��/��t%�����J�1��2��rh�b�f
 >�s��k~��һ[�[鸩�EN��R�ho���kB[�c#��,T�ѵ��Xr�;�劮X�",�Ü�}�� $@�0`>yT!2湭���ʯf����h6dY�\���>>6���{���-���8w��}�����-�ˣ_��@>���n�B��kq���_��M]�{Y��E�'��n���=�)?���6��wl�dG��5,�y�)eR��sqk#쑑p5�Y=�+M�s�ޞY����(B7��Ãb�N�a_|5���s�:^�?��xJ�>��겟ŗ[�dvޟu/�����ŴRDށ�܇5l0L���r�F/	�7�a�]%f�p�ц��p�/l5�P�ӯ��{�����j+App;o0Z�#zb: y�k�_Cw; f���gD�,���P��03 b�[z��#0���7L��a��q�r#X�+�D��![�9��ӯ
�p��ޗ����{�.����R�F��4o@�ց�cMf��Bx�6��X3��ꢘ=-1����?��!J�X9�%e�}6T�:�����j��7�y���w��Z& t>~ii���F]0�A���o��d�$�������a��p72�U������)�Ý�Tyу�?)�_��p��o�W��� � � w�][�'�fDYSb��8��,�1��Ńy�X�k�]�.���d�jg0ۚ;¦9O�m]��$��3��!�4d���Y�A|:R[]*]�q����s9-¦�G���U@�q�4)�s
='^rLf��*�$�K[:]��WK݂�����fvN�F���v��)ўg��n����_AX�fؐ�w0_c�C�M5	Mp0X��2k\K�E�q:V��\�[= v���_`�
��g_U�M�t�k���u�l����ӵTC������e ���ANb�)ٲxuX�3�q�qG^n���v�nq�.E����wq�ZKGgwl�ɞ��ԿE�8�����5� �\��U��E��P'����Ձ� ��"��Ѿl��GKB�n[o�
�Л���l׹�τGi��ۮ��æ�z�݆�}�96���5��K��\�Z���淍(l��|��앎��B1���\✸f|[��黓�f�Zh�;,H;�0c�ظ���Ao��dU��p���W.�o"�͹�ff��/]l
�2�Uv�>�AU�_Q���Q��8�b �Q3U�o��5���wuݛW b�w%�pv���q��v��T�oxs�}��,"����don?=��sx�xzU��(Ŧ�||\l���Ɵ��Ʈ��{z��Ð�����_�w'��s�ϞߵF����``�љ�j�ߥֺ5�[1��^��1m�.�7�`,R�t��U�1`'T�R`��m��؋�)���4��{��hsE�.���[�x�aDlUԳ�׍EՉ�'���.��} O�M�� ���O����wS�0걼I��C/F�n�Jݠi��@�/:.�"�H����9�^jr���]:guP��3C?� ���[n�$�w�-jCӆ]5a���R9���+k��oSzn��jCZ`
 DZ�U��3}n�[{o&&]�U��D�j;F��漏3�����0�)�48}�+�]���̭s��`���q|�f�^����KN#po8�
��y��"�h��y�н��\y�ܨ`^]���龫��O�ޮ�Ū�v/EV�P~b�y5�%-��,/��8	��/k5s�%��a��j��r�D;'?������i����L�J���� �F�8P��B�f���.���?��`� Xw�`/[�%��q�ͻ�H��:�Hnr`����t�"������q,�cc��ʆS�3R��eWǕ=��5�^.��8b�q4DsʃҔh�4�h�����N�{ �.��:��]G�AH"�;`:�q��-�L����K�Y��*�tp�5�_�����8ޭ��0�q�y��f?+WISoq�W�8�YW۸gPF������@�jɰ�Ѓ}/��%3��ͺ�������wĠ���5��6 ]=ywH���L�R�F�_k��2��;[��%��ʀ��}Z��e�7�'TE��3J��T�u��7�G��2�A�3�8�2+�� l��+���e�����N�t�3�+ӗƠ��[7��^�ٽ�+Ѹ�@Dq>�j�cKλUӶ��Gj���l7x(��<'�K��;�@�W����k��M��ƭ�#FUm���I�%�(-��Z���5woM'�S8���/'[�֕~��� �����מ?`�'�}{x7��&q�'Yf��0����)��?ehH���'��('�4A����{�k����
�՝�m��Q���u�p�֠����Ʀ�ϸ	�{F�������đ�kڈoH���7�W���
_K�k,u�>uL���kgr���g��5��כ�0I��N�uE�O%��=s�i�m��r'dKeR$Pf��⭞��L`5���3R9t
,���O�V
���o�"��]�t4+ͽ����#R�w�ݶ��ޠ4FFUۥ|�՝J&]B��l�l�>�̽[yr�l�V��� g�0�`}���+.���~�j���[W�
���Xz���f�āʵOh�����=�� ^��^�S�Mï�6Q�\�,�I�rh�텧Ay���<������Q�d`�����6�=Q������ l�Ѥ_\R�>�@v�D���!��Ɗ�NI�ݭ����pa��%�3�s��R|6��+ ���xP����w)F��}a�hwSy+�K(Y��:��v���{$��r�w\����a�;"�ħZv.��ʭ��.�&����X!�N��;�Z�����>U�U�|�}��)�x�_�ne,]&�-cuVg]�ů�oD8\��fU��(>��yUv�8tm���ʋ.Y �+n�%/^c�t۫�]�,f,�lB���l��"KQ|oM���"K�2�2�UU6�{��N��W(q:ж�J�g�v�e��*ռ�l#���D���0�ܼ��������Ꮦ��R�����QVb��|�0u��g�Y�&����� <3Y5ysl"�`����e��"\�c1lVЭƞr��;~�! �5��Kx`�]dc��M2�ԣgU_e蓰�X�V�Cs�J�y�ڗ�LJ�KT�{;�b�m���B���������Ba�r�Ý�s����rm��&n>hq���NΧj��
����sMv�i��!�uv��&�bc麃���Ėd=���{�r��PU�::�{�A�aЙ��q����#z̋O��ڙ����Y�8���S����P� �zZ4vV�p�=��G�T�S�n;ڽEҵ�+7�8Q�ѱ��9�Z%9���F�3o�URrf�,q�c�BX��8���'�:9<B�1�P2�����,*�v���ߍ�#<|�tD4O�A�;��:	"�ń'm�����QZ �}=�Զ��f���5�7��5���;3�w`�(11��Z�8wgv�$�Y(U>9mz���5+pڐ>ӱ��iՇQ��Ɉު9���_V�:��u��s=b\Z�s��n�y�^�E��)a�aP���2��-���w��i���1҅Х�f�M}vܨ{�8e��n>����އ�R��p��ٽ���-����j�]K���n��.⃴����j+MEj����h���+�j��K�:���{��	��%�<��t��:��c���ݱb����N��9n�7�pM��jtk��4�1a�O��;�3�k��Yw�5�b������3�b�ZT}O���in*\A���ʫ;�	Ʈ��qI�l���#FP�Ծ��U�9d��`��KwθT{���H�Qw���pp/^�dά�O\z�(��#��rtC�n�M�%�&NA�y�8u�^WM}L\k���ٴ�m�Wv�]�J8�\S���W4�P�톅*62W[A�`�c����8ɫ\����t=����Z��,�<_m�ʡ�8�bI�'Ӄ�Մ���9���v���}G"�Ϧ�����cwG�}�����K�cR-�˗��kI��j�SL�sTN58wm��{�N0]�m���ϟwtP �,A� � G8p�c� !,h�n�cM ��x+ߞvtx��v��̣K��(�{g/T�9I:0����>B��eM����ÕY�Ui�I݇k�,NE<4�M4�寨ʖ�h�U���^� �%��؊S�Fa��=Jz�II��J�R�%r��:��[V�Ԕ�F�a���>z�{����^#OQ��)�1� �瘮0`�M4��2�XuIlL�'*����X�G�#judwT��4����Y���9]�v-Dҝ_.J�C��/%i����}Y��8�vu_�9aԴ��x���r������7!iO�ó���O���S��$�t�p��)�4����"��yh@SO�䇈�"����" �>p��I���ԗt�<y�Ug	p.�n̘j�����(f�yδ�Q���(�v�W'�v�z�����y�TĔ�䥱�p`��:n-b=U���kN����|�xKCz7��-�hz$�A�7��?�/�����M�`�'4��Wk��~�<�S7�Xʹ��d�q3� K���ϋSw�i�6��
�0 ����OJΦŀP��0?�,��g�Y�{͸�l���%H���p�{��V 9�A�P�x]�8��-�	�r�Re�{�5�����Foh���bʠ0,�D{�kEwD�g�;�1��ӗ/��
D�5_L8�ͪ�5M"�<��u��Wu�O��p^��o^[N���~�g<� ݵ���{ ���:��<Zh�;��n����ۙڛ[��� �8bSDNfx>d6��u�ɹ��E=�L���Ft���n��і:�Gr4�WfVu���ULi��{M�X����6�.mTD�dx��c���uS�z����uVE>S�!��W�	#����/m�k��v
&[�v2�%�#0k���.P�y3-Hh:�tm㚦
��+=�ɑ�O�N��J�FW74~��4X$�B�BX��C�E�.��Z5v]�6�s��*`���r������J�M������p��ƍ��	�81��$����= � ��1��9�}�dS}��4m������t���[5��c�1gm<كV���I��]O�[�DXe��V����%�����[*{q���s��+m]� _��B+�~�s��y�83�qZ��Ah��:�O�"�2-�kqg�ulj�8�np�� w��Z��a�y���6�tS��A���WvL6$����
O�k�� /-�����[M�s8�a�8i��l�\�h�Us��ܦ���3�^/V]^��H+`���d�{�F��Q�Ιԋ��<:�B�>�f���mc�r	��
$����:�ƶil��o�8i�.�cXўUס���8V�U�V��<B��Vg�/��D��L	����������\�5��w����]����]\�����*/���@���a��w�/e�<v�{->�;�C䣭{$dY���t����
�V��|��3W��xj��{Jnt�R&�w�;��`�f݊T=r����������S�\�f�k�����h@�N;�5�DUI�.�45���N���лw񌛔�ȱ��V����G��B��#�A��k]<Ł���+ǅN�:q�O)y�99^W:��NAFCC�?�% � ,� � ��W�#����?`a��M;�u�׸D���|��a����'d5�Y�������e�J)��w[8�RDx�/�;\��(I����2�K�!�,�J�yז��36C�h1Ť���1+�
`,�E0IDU���]���Z��L�X�BS�/��)�:����T(tvN�8�S5�#����Z�V�J�Er���u�)����x�m�n�٪s�8��m��%R��_{�ŐvZ�f�X�j� ��s(8Xz@��'�@!�^�޶��0[��ѩ>a^�Δ�����5� 3x&wT`�hkx��n
�˥l��Ų���b�Y{3�26{Ima�x���X@�	���	�Otu*�i�1@40��;����fr�{���s;������rZ�+��.���M���gt�KHм�۝n��6yE�r�g���h	1S����̝�;v��5���I-Iy�kn�l��wn���R8�xQtJ�l;��0���������\�8i⨷:�Z>
�=������T�Q����+�1�^��> ��ܔ�W�|���;׽�>�ms�;W�z9*v6o�/N�Xсx՟������w�3�MI=<^Y�@��vPM�<�E�0��t_.��Wx҆G3�1��`�)�ڛ0����M�� �o0ݯ8�2(�+��;��	��w�����z�N�,������ƩZ��&�9 \�����"��M��wZuox�Va#�%�Ek�<Á�������ވ�XD��K⺎��f,_�zj��q��!�]c�Eg���Zc��n��5�5�y��SW,*��L��@
𭕖�v[�u��מ���*>6b����D�ޞ@j
07��*9.�|��~@{�9�J=�bw0��
t����m�hH��)�@���m��涺�5��3aR�)^�z�%�.��v\ϯ���UW}Wݭ/����ۦ���g��n;�o��c����}9=�g����E��|����r^�(�Ty�C�\����k�.*c����NA���*p%�3)�9u.���U0EX^z���R��՟c<��:����g^��\ֆꓗ2��r>��1��/��$^�4�Di�&9��JE/sKq|���t8@�N���-?)���^-c��}���o�����*��ۛJS��]���PM�r� M]�Kgk��ͭ�;ۊ�!�f.�D��E��+F@O=�ݨ����ZO����Qٸw2�B)i�m0Pg��-�n@
���9W�}���k���`�3r-T��t%��]Õ��_͗{ ��wv�����ym�ju����"(P�����e���cU7��Ff����5h�b4	����+�n*��Ve�c� �M�¯��-`�@7j`&��<�4%�a��#����)^Cky�v�7����2.7K^y��w;r�����5Y��F��A�ԙo1�̡y���z��63p�$��ꃊN�w�����V�}��e3�~ѭ���"�M�k76��'���ݵ,�)��{TH6p6���0��᫵�Xx��e��j`)�ou�|���闎�6>�ɨ���&��I�{%�x%��*���oS}\�v1
�C�=K[��Hr{7�R���#]}b̋��xZ�� Ѐ�H@^8w�Sw���\�B!*41������n\����r��Q���Vj ��كo7`�#����,`/R��y����q��v�T�O�bg�"�u׃�s��&`���+Z���ݩQqI�G���AE�wS<l�xsP*0=MfBM�e᪒�{����fL
��;�l����Ⱦ�x�q�ˋ}���U@4�v�1��_���y�u��o�9d����x=��w[Bs�b��Iy�ܶ�[a?�k���?l
��:�w�6;�����M�5WJl�>�u*��ȉޘ��}�P��@���������d[Ȣb\�ڀ9���lJ��v�=�vx6��#�Ц�K��;�U� ����1�?]�,�u �2yvHY��CV���`P��:�D�"#74��@�@�ݮ��I���a����r3 �6 ��i�1��HQbOR1��(�Ω.*��wTMoX8�HQB��d�Ax͚�>F�#(�q��'�����!`$�ݯ����
�6�L���G��v�ە�澙l�oݱ����?���AĩUc#������۱h�z��ӛ�`��P���������w��Q[����B;$�h�ӌ�ㆅ?�3��\����Ͻ��]��+�
�t�]�W@ɹ�2ɍ"�����"@d@$�
Y>ݟP�{��,	�A�6^�����X{'n����+�� �R��U����}����&3��xY�J�lP��B��K=��'��'9��Ʉ�׀�5��{!�=��f�X�����{;���M"�ne7j��J��5���E�����u�~�T�����B�ѕVHNs���o1r��*J��,��H�vY�@k�펺��%(���$+�Y*	���<�@�mH0
�LZ�u���j�v-52*�:l�cz�狩|�v:���q�]9�C���"R]=�!G=[���mEF���C6�wG��^���O����������P���Jc�J!�-P�p�M���;;[���̪,x�c���)�!�� rW�`^mk�銙i��s�~�K�5Sy��A긓��T��ɳ�|4!�dG��]3A�Yg��3"�P���R>��a�ֹ�'kBA�/u�i!�����xNr�o�*�)n�5�H��^�N�g�(l�e���/~ʲ�X����.����#�a�7s���;w\8Te����U
����,0[��p<��� ���Or���Y7�|��
�/�pr�M[옿uo��N[w��ziH�Nu��u쁒3�K���G�;6��.���w+c�t6�B�Σ	�E�hi{�{0�]\��ۛ�;�U��]��@윜}5y.����q��y����= �f<cpW)����>6���Kv�9�.�����SU��T$��5t��n�o 2��{�C�|�������N�N��#��\�	J	>��
$6��ޏ8�SD���u�ͭ[�c`40�ְ�N�{~��0O����[�cr�N
��E���&�eQOȚ_����/@�	���W�����_�v\	�k2�=��sU���{��F)Ћ���l[����\����j �=r ��7<D�>Dr��zw-mF�9�14n���jZ�t�#5dS�NG=��]����1"����{3G+ݾ??z[G�)T�=����3S,`��B��H%���.F5�te�W`�������z�W���[Z-|�]�UfL�]9�l�������ëej�ǝ[K=���Y�D���Hp���|� �0��W˨�H��l������5]�}���>���w���/.byR[����^J�W�s����-����x�Hm���S(�{}����yqՓ�f=[O4��zBO����ֱ�@��UP�@eRjyss�Y�&�vq��f����1�t���˨_NOu܃��5l�&C,��rjp�ݳ��-���{3�EX�=�7`�����s�Ԫ�.�Rp7n���{����'_�	�-� #�@���OT���{���-5�,wvК��e��u��^2Vٽ�Bgݜ W/��p2y�
�3D�ʧ���YOT��=�o����_"Q���p.�rzrR�l�	���۟s�;� $@�oQ}��pɂ�z�¦4�>�(%��c�cC@_���,���"��`���9�4�t\�nm:��:�wH�- ��*�Ϙō�cadp�����f�"4ҝ������ΪuC=�+��#k�ф���D��ed��mY�H���0M1 �Rm�N��{1�pة�+F<j֢,,�鬭��z5Ү<�gu�o+['�[�}����o]nٟ����Ŀ���p��w�ns�ً֣�E�,k1��܌5�:�Z��@�8�]س�z���O=�.U������S����1-��l�p	p7\��0=�U[��[m::�-�a���_������%�-xeۋӒ9xך�ئ�y�B�t���Qk�7���BoK�{���!u	0z�e�S&���L�X9������p)v�4�A`�>)����Qk`n�J��<M�죾��5�p�T	Vm������e�4!��=5%�X6Uf�Y�`^xY�`8a�E \��IR�weW��3��FC�MeS�Fn�)��7`̟P��d k��j�\lddwV�aŐj9��*{5�m���]�>�ȉ��5#a��l�q�;p��ݫ���{3v��#0f{m��D?Z������k�"�� R���� ��{���O:�#We~n�7�sse���vm�`�SP�I\"K�ۇC�[��Q`��X�������UZڌ�k%�f6Ş�l�IvE�y-�Xu��rxk��nt�2���ZwƔ�gE�r�6^^+v�8��^����뇜�͜��H{9�WM/���q�8��Iq8nG�3��2���=�六I�7�j�{P��˕s�U}:ָ������ac�G�l���[�BF&p<�.�mgc���T�q�u�.�o��0�#|��g[�;TYYu}V�7��au�C�q�}\���e�}�z�짍o�j3�6�gR��6t�,��к[J�F�l��`&���}��"�U����+�Tf�F�EF�G��[������tQ�3�S�Y�RXb!��\��XWhm+��-�����i:{���zp�W�)�SB��֜m�雡Yc5��~��uE$h襋����5�b���������f_M��qi�MI��^ɐ��.����j9��f��_�1��s��S����|,����Ӌ��l8�ؖ.IV&e�VN,6,�+[�xҙ�ּ�]����\�i�e뵕!]*K�p��@ξi�u��,�L��hK�τ�V���;�.�����̶m����mq�]��t��C���� N�N"ɹ��2��ANuI���`��'���-^���o�c��;�h4,X^U��1�b���v ��b1'�qX�7�X��bac�!�@*6��1T(��	�:x��~�_ h��0�X�u��8��������0]��L�~~b��W��4r8V�D�w�ׄƚ��`��T�`2Fd`3E���b��@I���4��\1������v�a��c��k�*���R��K�/��%!�˭����"���2ꉗ	����ҭ`���#EU0����Vhξ5}m`��r�{z�����Y�*jU�Na�v敜��㏡�g'(ņ��
����%<M��5y���~G��L���{�%��N˵[AJ�6k�Lv�s?G��LJ5$��N�#���	T�N�n�asm�kR=Ժ�N�ˮ�"��:�q�#�m
b>���9VkZ��e�+�Z�!��7�w\�wj�m�����o���A�6�p޶J��n?\xD�Z��&�MNܮ����y�Dy�b0�r�amtx6%u������U�]v^
M)J
X��FNfn�j��k��uW�4��w���{�.����X�$�j^�f��Z2�+X�H;����T'N[�R=����6MЧ�%�v���jp��.���(n"눥���ǴZ����1����z���v53+�<��Z���,�EN����$����$)wi���/ː}���i��uY�/�SzJ}#����{&�rwt���>v�v��;v������:v��Gn�:t�U���o:c�<N;=<;v�:t��<q�ON;q�n�k��z��]�};�Uc4����@D�RO
pR����QLt��΍�"���x��+:��o������h~Hz� R��
O�
B�`��������d��H��RU�|GU;�׮��rZ�PҕAa��Ɵ����Z�e��B��@h��ri�j$��f�|i���T�[������͕�8 �<A��M>2�\��vKR����@�t#�9R�P�&�p5vxa�#)/܌�uP��uRw]��U�wV�
p��L4���S-���喹b-OrrJ�[^�<����R��zxzi�_#�jK|��e����!IM3-�A@{u�Փ�x��c,��짇�ǆ�ת}G������T�RҔ���@rZJC��
 ��N�<��"�ob����0M V:�h���*�bm�¹�s�̘P��\�^����YԵLvGn�M�8$�P(��P�x8�W
<9��]�Ve�I��A�oPᢀ�@�ł��"�7u%a���@? ?"��hg�|�����*挥��ʷ"�� V�DvW�FG:)��'V�C]��)s5}�ہ� ��7e.�i7��0�?/��fs��73����&����׹�ٮ�A(�5vy��cM�X��6�ɚ����36k�u����ˇ�N��f���&��*U�(��2B=p�9�3����6�Z|!�a�6� l
7�Go}��t	omI�p-�X���<�4�����W]�V����|&3�fi(���쬕A)�=&+o���o��l�g�4Zi�����F.��"�͜A�����*�k8��#�˩�lM���.�鲧�fUl+14�� ;8��=�g���v��ZFh:g)
��-3�0�K�+'�%n4q�Mw9�x��Q����D����>m|��p����4?Yk��Vķ[�G��<̳�e(͍���eS�k�ՕÐ�v�]�|2���2[��\S9��6]�n��9ܙi����gV�Ң��4jcZ�[=��P��������եMȲ\=�:�tѾ=5ac^8��{�#� ��� �C �)���+;<q�>z�qA�Pb3똀7'���Q�QFU)��x6����E�Vz��q���|��lP�13Ǫ�@T�`ڈ��ݻ��/~2�I�6�̫���~�[��W� i���v�1�_z��jA�t�T��Y!]�����ȩk���o�μw��L��gk�%�C��9]�O�b��5�r:��ޤB�;��`ޣN��}>)�y�aQ�ٺ˸�܎�,k؍AV�|,t�̞����,!��I���ཀྵ�|�lWu�ӱ݁-���<��H$5�)���;����Nޠ����q� �ƃK{"�L��R*�h��ӻ�q]W��A�ٯ��;�ƨ�h��`0Kn��#�#��t�t>W����M�l99��,����D?yN�	J���|vК0u��F7ЩD<�ڌ���k/"<��i�DU~�Ӯ�M�w�.B�]�y�����i>��d�Z��B�K����<���"?�{�eW�����F�mɓq0����.�Ν3��MnP��Tފ&���V�j��Qv�ۚ��Wt�rC!����|p0`*�dNtv�	̯�iX���PX��@tE�����{�vG�~�������o3��l�G�S ��@ʸ�diM0�J��}��ĺR76v�*��A�"�E�o5�ؐ���#P=ZmM��f���T�h^��vH@B�sdP�`/̯�&�ׯ^���_�鹅�+̫c
���<�w�m<��4�@��l���Ǟ�H�0&v<;�6����	ɼ��i����MI5g�g0�3�0f�
����-6�HBݑo�[�Q-
��/���uk�hJ�F��W�c������*�6�@��DMn�j��{�8�������w�uY���.Q����B�i�D��^:�sz}��(ˁv�B)tyxwl% %<v����"��9l�.�xg���9V����J�p/��H]�Y-��F�2����ʦS3շd�BK�ٳ�/�9�Q�9in^�;�u��=��Α%����Z&���R�xkk5��S1>M�$"k�4�m^��S�l�vZ�J�,�d�;׶���՗��@�IUrۈ*�T-P�irզ"�j��#��,A�#��@����v]{�?_�Uh
������@1�R y4@�{:��"��_'縫����xi�N������d

Y��Cf�9a�q�;,��ܑ�����^�{�����z�wcFP��fn-ڶ���;�hy�5�/V�xZ�F@{\�O���v�Rd�V�Zۚ"�Y��D�M�w�V������w�~dfc/f�@~�#�lB�ʡ;�`A�q���X̌��Nt���G��x5�p���W�H���Eٟv?�&���Ä��ud�I� �3�Z�E��9�- ���q3t>7�n�tDW���>��wC��_�N=�|Oo���{"L��@@}�U�]�w�CLs���iAj�3p��x��s�����_O��?�6`�z0��^Q�뉹������Eɲ�V˶z4S{8F���1��x�
�u5�3��~���'u��N���$�"����W3B��mǋ�{�t$�B��H��ÊY�m@�\�qP+�.8�@�[b0(Q{x_>�)c���kն��n椅����]���'{<�u��]՞�o�b��#ƖU�`�@b#�L�p�[����	x�rr�l���8J��<� ����W(�~S���J��z�+���:�S��\��Vc���Ԁ���o6b1��g-ޅ���}L�cre5-����e*���qV�x�34	Mp�uև��۹���Z[Ŧ[��k��h��Gk&��UTX=<������������Y�Q���n]��WkKB��ݑ�Z���A�s�q
��7-�N4��mEi�.�L�{KN�܀_�S�K��ِկo��r��5����vM�;9�p��C�a��g��wW7`�i���y�;f�u��n�r׵[�����~ ��IqVfs�����,�c#�p捀?���+�A�B�񪧾�<��?<� So)��|��]�T�K��<!ܥ'�ݢ��I�A�	m�>�3<���7��d0�8�3H��`1��43N���rcT�c�����9��hx�{u���Z
��5�T|�u8i̤qHi�
��ѷ�{� X#��(V�q��G�r��ͭy����1�9�]M�W�\z��/�μǳ2�-׼`45�\5��c��hbWu��@� y�����kp&�����c��byxRx��(�!ش�]��k���T�-խ����[Բ���{M ��W���?s9���o�w�����bT�u���Yr�x�ھqT�(�r 8�M�P�/�F(�1��P�I|1�0�l+v�,�������������=�?p�=Gm�W]X�/���7������w���@zC��sbG�|�}����N*>!)\N�\���v2���۴	ɛ�w�lp5�x1P�&yx�k�fljK��	;��|o�l  Q���͚o{4.��]��^7@;�LUq8\�縱)�M��3�����|�q���wǦ����p0�E�ꇉRB�w�"&��b�dnhB齂<T���T�oV����x��0�+9]8�ш`��mu:K�{�^H|ƀ]B��H�7��;k5�0C����e�^�c��ns�3!ܳ׸Sב�2�JKG�P��y�U	8�/o���=� vh�mU;������Z�A�S����,�>CC�Ue�'���a�u�o1n�U�U��Ȧ�zʷ��e�C�e5CF�;�y��D���1*ꫜ���r/����1<{����<zC.�D-2.:+���mp�i�^U��H�l0����/B���x}�5�8c��8j�լˍ��UWoZمo�a'��ʇ5�xd�	=tⱧ,N���`0m� sP��o�ͤ�ݠ^�fm�����&�|;>�\zr�	J����}�қ�q��%��B����)&�ѻ�cD��[�v[SG�+���\���n��cU8,��M��\��*{��{kj��WH�U��o`gd�H�T���ލ�&|CE���ZF�u��l6��6���X�2�{ݒ�{��nԥtU�`ȫ�˼��t�6U�[���6���5�״�i3(dꊗ�Nm�t	����(i�h��-�a�H{�n��V�3�G�tT�����#������|�-�� > m�`���rZ����%�vOn��{M]�E�B���� E�+E�{O���������`��l�UX�,C  � %��<�s�7.���J���ט�J�y�4���Rt������7���,Uvq�l_b|v'D�ͷףd�~=I�S��-��T厺���??w�����&�ݴ_�Ui�?�����qƐ)����P���^g�y��O9������}'�o���6۔��.�����]�;�OwA�0�-��WSs�xЃ�@���~<�<y��d^��p�6i\�=� q�*�iطi�ᣁ.Ȭ���'4���'�S�㌆���7�}��:��ݖpL��c*�wM܊�v�+ ��ܦ� �1�k���Ȟ,Ѽ�]�]�hv"��p��w�+5u�bI�����l�z�i߸�3=�͍-B��KP%oA���LȮ]!-���~Ɯрn"�>롋�֬�]1XZެ�ҿ�L"/j �{=>�둸ztE�j���>�X�D��R�<9V�om��B]���8��@��Į�����&����}<*R����s��Y͐���Cg�o7b���} dȻm$��/J����z�U?��"���5X�)|�(�[��eor�!ey޸�d�$�Ӳ�랪��T5K�GM�7�E�2H����P$�����iλ�����b<$�Ǽ���#nN������&����l�B�"�t3B�EcB�,x�O*�W�]�Χ|�����G� �ָ�ͫ�`�����F�����K�@d��fa.�`]��/k$�Ḣ)��]nqŸt1�W�z�����d��g�� <Q�
U���`��[�J�uMT���aA`�.��F�@CXŁ;����U|���ٻԫ�m�4�?���h�Y�W�� R��5S@J��
Z��-�cC�gC��#uz��wj��?MN�]:3p	�0�T#Od��6#���{!R�-m]�}ܧ���N �`�`�L�]�7���W���R��	k�[�*l�àZ}[��[-�C��TT%t�C�D	����3�=��׭��!���p!'��}5����̔ ��;O|���'�8O"�p���P�A� �,W��ז����K�$1�+E�-<w^U;A���ns�n��T����=1��,����˥��w�����)O+~��*��ߝ�L,�"��9��7#���-rA���6��I,"\W���G�b��g������r�Z��?rk=3��p���z.���Y� �"�9��h_u�Ne��t��y�P�*��U_x��y7��f�7���}s��{�:t�������-S�����c����]>��&@����.�i _��ͻćN[M�gJ,9�1ehZqac̈́p^��i|="$	]ѹZg���@4�u9=����QXI��:�@+4�g3�6�ǣ8ȹ��3^ ��A�9^��ap�vr��c/�ݷ��!��:��`l��K�C��Q�N����i	�g�u�h�p52 ��ao6)?�4UWq5"���k����aaG��:��k<ڣ٤G�I�˩�lR�I�%-���09�<	D�D�[+�1�/!A�x�T����V�Df�Dr��3D�~VyL��F^�+"����;��י���]����
A1�x:�\T �=�o��qQ����H0���L���	��B58�*njmn�'j��d�7I2omV�TͰ�����Z@��u	��2���ܛ��<F	:�mRx��
tjf.�]V��E�0��j�n���G�Hn��*��S9��R�P�1Q����-D쬴��#��#��%��v��妮�Y��4�HfW��;���:��6��kI؅^&z��RVu*Hb�;u��WbCzV2�+M5�,��J�K��1��/�X�]�+�u��D���N��o<�Al����D�w/(p���QCt#=�5�-w���S�H������"N�&uX��Ғ:���[+���+!��L��n*.�)\s��M��ȞnV��ә�/�l�V��S���0���ջ����ຣ����\pfv]GU�����NoN�=��Xe,٩�I�"o�f�T��./N3MAQ]j�T�`!���u�к�>�o���7:���v��������q�{�0_;���j�V������F�R���Q�S��ܹ�7�t�"���\Hӷv[J�=ײ��,or��CS�8����l�.+w\�z��ѕ��E�r_fV�L�����"�)8wN(9Z�e��U4�4^1F���β��Դ��#�*���Y�).k����u�)�i]r�9zi����F�h'`�dۮot��k�堋��w��ܱ��g���r貛	�G��]�����^sL����G��
\8 a�<�0\Vb�:l
�w�xk�^��pU�����߸=,����D�ct`�OW����
C�
�����,H<��~8��eg���>d��W���%�U����_�`�XϦ�u�\/>7�Eu���n6�g*�J/�VNa�9u�[�xZ��jv�5�jYs.i��5�0�����yy�W]Ɛll!�<Q��	
��ľf��XTs���4�]�,�{ک�S��1���|�&�=��W4������KLgm������<�ܻY3��ĳD�I��L� ���!ժ&�g*��
�S��)9#��v��@ټ|S:�v��ϥ�� ��'�d��1߆gh��V���9	���1}ݯ2�cW,�J�W�.]r/Ko�%i��Z�X�a}Uݛ�Y�}R��VJJ��i����l洮���U�#����V��H��_D8k�i����XH�G�)��W#��˦\�̨�X�湺���ق�#o*M���A�/\�O�^R��l�`��c�.�=�jg`��Ӯ���L�&MV��"�k�g=�whS��!nFp��l��!��ba�~��4�ٽ�/��KV[-g�96�"�*�뵓f�>hj�SԊ�jL|+*�)�5�#����嵮���is��q�xH�Ub�~U��qwBy��w35��ƫ�>ٕ�ow����s��M����B(Pap��cE�P��5b�sa�����^��.��=I������ �e�gU�Y|�?(ꖖҝ�zi�ϫ��VY-�ӕe���b
R����+�Ԅ`�a��}2Ť�KI��ub���F��4Pr^�PD)N�;0��ŦYŵ�<���j�N���aJR�}�>�����S��OM0��Ke�Y�WL&*X�(}I���J�ᇇ�a�(��V[Ib�&��4P{�@x������,�KiN�=4�M>>��Dx�%��Pwi�ˠ��T����3�GT�z��Ƙ|2ʤU�����}�!T��Qch���"B�.��N��jZ�Jt~�Ɵ���
���T�,TS4M�L%rj�*������KX�QR�TD��� _� �I �<~ʹ[�CnX��9������/vv�J��������&aG�9�5Is��:ܭ5V�[-Ԇޒ�N�<���$��N��wp�v������ݙ5��~ϩt잷�e���W�TOG!�m�3.q����?������*@���;l�q�}Y*��=��Ʒ�u��8��s���rk����W�χv{����=��{<o�Em8��2ifZl��b��7�w=�X��͡�����M�PN"�������ѯ�:��A�N9�dB�>�U�~�C6���oP֩��ʠC�;7�l�x�ڤ�NX�gzՑ���ƃ��5܀��LB�U�Ub-�8,Z%gu�)�[�A"��5f��p;{D��w��R��n���aZ��[���^�����f]J���JO��,|v��O��'�%�&���*��I�b����%���X�)�j��#���v�����r�I�a���z^0q�bEr�,�d�a���"8��~��s/e}3{�xut�5!E��*a���>tk:�и��T:hb��t+����9�����3;#��`��� A%�A����\���T�dl٥�XE2����_�ֹ�����M�.�Ȝ�l�&������G�����`/����]t�? NgWG��ݟ|}�.���
q?|�2���������*�^�/	͡�CQ���%�mɍ��{VO0��\�M�qa��n���S�aos��M,E�hP֤9����ǌ�b[�ms����#�4����a�C;:}<5������0v f2�{fJ�[�>��L�U�"�ۨ�^�<�1;
1�eaFT��uj.;v��&S��Nr��r��o_nK�{.�f��!8
�ww^�Ou��_Sk:�E�nݜ�r}�r0n�f�m�u���� ��簽ڻj�w�s#c���D���Zr��!S���;���D�7%��"��\�R�軌�#ohjD�S����n�`;�j���e@ɽݜ]����kvl�X�4�\fϜ.�������������oeO�Хc�ߛW�
]*���rs.�B
���1s�p�=Pܣ���Out�,���{i��ݱCc��v*��/f���-��1�H�c7�K���K(����'_r�H�*�R.�U���ug�����#���y[�  ��e:
����C�jI~�ޡ�� ����@��L��t���bwcD֌����]���G�M��K�N �<�@y��}����0��qu�,3��JXWT[+�G��=I4�m��;[���&���6�z�C��_#Cb�aE�ݻ�qѹ,_p�����N���!��xC�:�� r�;Q7�KdZ��<�t�l�J��Y_`|�p�jC���w�3	t��ɮ��ͼ�T�9�L��"�6�Q�S���@woS v������/�b��z�`���S8����!f��ಝ��i��F({ ������[aҽ�~9i�\�:f�Y���O�+-�K?^A9o0��t���Ewv,gs�͉z���WK�=H����ZCf�(���	�_i<����UG�j|(�nou
Ǽtg���z�M��ن��D�v���^wu$���Z��siV��s5�!ԣf]�wN������kδLb�K����sBL�V_a��6�>;�#yu��`�;�t!����:S�%�1W�S���89�Z��!���&hx
�&�+M��̤�ؽ����mm�~�v��ԏ=��E�xW�9څs�Q0�"��,�]G����޻�@!�����TYin��m-����B�E��2�gX��ʷ=�R`�Yk{ݰ���0�GVx�O@a�l�Z�t�M۲�o_��J]��Ew�T�*����Dٳ���Yac\�Μ��h�{6�rY���p�FT?^kl��iպѨ.e�C�9�1��g�����p*���1q[��j�Vۥ���3����4V�76�M��t(ʎ�Ν�#������/Xwi�[��5�d�>�`�TH�g`����5w�l��cOp´���g�RB��Ʋ%��ʮ͚�6*��;�Qf��8+���5@d��*iloK�ܗuS�l�Q:�Z����}�`������g5���z몄o�C�1�&~�x��7�l�r��M*wu�N��;����GV]TC+Ï�Q���u���&�s'���ej�:;��=�xy��3���\��5z��m� ��A��ٻ2j�����Tݯ�������p��]��f\�񈺧���D��/)�6DN�k�iL�j�Y�%S�y�YU=ÌUzX̭V�>�mF����.�{U1�X	�dQ�\�3t��
|�qM57�Y�]�Ex����].��Lc�TS�=Z�����v�4�k���a��ݢi�ҕZ퐺�˱��x�0Ȑ+�/�0pO�xMīA��<g_"0lwV7�:�@��{Qw�Uă�Zu�T��f�p�����,������.�tPK����R������`6��iL[pÙ�j%�����FC�$�� �P��������]�-����Efn_W'ضة#�v ������/�";L���ov���2����-"�o�f�٣/�in�a�@����B��m����D�W5���&�+��/�T��eţ<�C�4�.{B�m��;C�WUvq�^��+�\�z��b�GԂ֐Gp��5�,x�.*���NY<���ڹ$�x���%!�k��lx�]��b��2V�w�����S7VR����@���[����v"�Mp"n~Y ���-ۮ�)�k� lh�p��8Gji�)�0��}}K�y�}it�Y�r�+R�@r�a�_5J+*C=cҬ��ۡ������� �X*6+��<qN���p�nbZ���:K_�儌t�6t�"6�Է�����57��<��Q����C7n��Nբ)%'tG'k���o "g��>-�⩜V��ڋP5�sp�z{jp�Fj7Z����'m����g���2��ش����US�-1�����w� �	�`b� �G�%M �Z�c ?L �zv0�xM��83{�w�X�	�iJA5�VX�ޑ�n�,���b�%9W�&��Z9��� ��X�~x�En��IU���k�PO%�44�`���n��U��`<#ʮ<���3d��٬}�t�����|'�ƖS�&��vXv�ٰ��S/����zݬ��B36���C6��n<u��F��R�ŉ�W;xN�EB��Ʌ�.�X^ �J���0:&��sUw��^���5����1�k(�f������\��B�v���5���엝@�@� H���2%���W��Ť����sUU��'9c`*	Z�wq�amL�t��E��'��G+<gԽy=��~�e|�����o�M5UB�K7"TL�]��K����<��9����W F�&�����Mƭ%�� DӇ�f��[Ҏ���� F�<ہ��z��2�n�ӛDγE_Ojgݦ����_s�k��)�Ց��Ֆс�ϚmQ���`���L�f�GC͓K�6�`�Cԫ-�Xiע,&8&�O�d���ɥ�i<F\��j��}��7m�6 Lʜ�������7 )��ݜr>qqְ]���O0ʻ]�2�4�]�B�:�(_��[��3��Ӻx8�N5ڔ����].�IpiI�ҝ��Vq%v����t9W�� ����S��Y�W:�m^�Ʈ�����ӽ���2`<�:m
�U͕�jfv���St�~k�f�c���"�6i(q�[��CZ�f�g�J�R�T�beU	��b��D�+X&����-b8�IVn�v�s��Qʘw9�gw�9�-���e���hZqT�]�C���[��;���O�,b�Q4������9�ܭè��ـ�K��K�����=h6�ꌝV��0�h�u�n�����΀�o�PȴH��Z�U���,��AzW�u��m�s6[l��nb�7���ǚ��Ơ6��. ��MFǱѾ�*a��Z�W��傗��n�
�8UW`����X��G;y��T���} �9��<�
���Y�8��6v�]�Mr��y�`���\�%�\��`�m������p�f����=�8x�/����2�,ˉ�Gk
�pr�j9�X3	z{X�D�L�\�	&D���̋{�&��O�	u�3��2�[r���s�i�A�� �����Zf��tG��f��Kw��il�M�lS3�ə���co�V��δ��Z�	�^��v�$�������	|UQ���+p�xH��k��'�>]�����lK�e�v��gk"��w0|ds"���(m�����ZeN>k�-Y:��u�[���mm�ѓV3tk����c�7�L]B��&��ܡR�Tcη�q�3*L#7)���sŰ:U�t9û�n�%�#Vǁ��H3jChv]����U��4I�˫�D��kԗp�Ytr�mc�r4ѐ}�S��N����[���۬w��C���={���}��*J7!A��n3{�^E����Oe��f��ǬZ�W=��mY�r����� 05������h���}��@�e� �g�2���L{8��j���ˌ�����VN�/�	*z�0a�����{=15Uv�l{4�Gs����å�	��L�d�AT�n�M�ԓ���L��3��<98���E�C[T��IU��3�ܩ���]q���x�����ŀ�/��.�����ҷ��|)�~��yJ{��l�뺥������=^�0릷��U@����<����޻�B&��qc�ex��W����@�ב��k�,IK�0~�կl�-�3�垾Er�t���H0�B�}܋)��k6Ug�ܘ��J�Rn�3a��J:�o��Y�
�Iw��Zh۽�/����c�֏K���m�]np�(uNօ+醻}sy��2�KzU��<|�n��֝���r����҈�.��Ӫ{v�p���ىw��Ȭ�ڈ�=�Tf�
�L�a��#��FW0*�i�]�_^�/��(�[Ƥ����+�(4�!�ռ����?����g��c�۫�ӽ`��J&�~���4�i�H;.w������;���U)��OYҍ)-��Y�++st���������_jeS��|7��R��ϸ���z)�%�I>�q��1qZ�&j:AU��m��M�06̋���v�آ�YNN�zZr�DKM����m�0��#��I�����xqO�o@�F<C��[X�̸����}�,�,M�7�`��7Dk5v�k({��b���,]S ��TSOtnؙ[�'/3��b 	�!a��|]��;�~������������?�T �
�+��QA������D�����u*H���x���t=�;	�D�PY
!!Ad$()$����IP�����:���Ē �wd�8
I!AH���DPX��
�I�"��Dw�HDPXB((HPP���B�'�p�(,"I ��!�}ЈPPB���@��PPB���PT��!AD��@r(,��"
$�Aa ���PP������J
�κ�)��R�KPX
AP�PX����DNRX
(,E��PY�i)"��J$�
$����]�AAP(,AA`�PXIAREIA0�	pP,���@ (QĪ.��x��<w&|�w�PF�H$P�$�}&����N���O��?�������;�	�����?��S��?�����7���?s���B���O�?�?_���~�T���G  
���W���	�0���_د���)��ETW�ϟ��������N���G���?�@��&�}��ٯ�?0pP��$ZE�$X�V�bE�X�Z�@�E��Re �ZZE�VH�X�i �Z�$�R�Y�i�f��	�d�i�f�V�Z"Qb��Y�hV�f@)��i�a�d��bQb�V�i��U�%F$dX`V�bE�E�E�@(V X�fE�@(V$Y$ZE�YVRE�% ZE�E�Y�iH( ��E�ZE���� �Y�b��b@%�f�E� &��Y	E�@%�`	@�	FE�@�E�YB��` dX!X� "E�V�e�`	$X$XV$Y!P�bE��E� &@!	VHYdZ�A�A�dY!Y HV$Y$�b !�iaR�eY�ZE�I�b��@�Zb�Zi$U�E�ZPB�D��A�DAJ�P�P��$�[T!h��	B�"��(%
ċ
c��3e�����QA�I$E�H�	�"��G�~��'_��~ߺ�R��?��~��_���������U�x����7��>�S�����n����ǐ����>�?������>>�����2��+�/�S��t�s�����*�(�~�� ��	U�$������:_ q;�g�$��M�~���>I�:�TV��~�?o���ꊨ���BO�a=�_��������s�~	��}��)��W ���}?�~��TUE~�}��ߣʙ)?���?��N���q?A���/^��>�$=�wo�ETW�]��,u��y:#���6{�3���a����� AE����I���T�����<��S)�������1AY&SYC$e��_�rY��=�ݰ?���aL�}�<�UT�DD�R� E@UP�P�TP(�� ����z�UT
H�(��
�*T�IT%�R�6�l�7wIURH	
���*J��J%j���ٔH�$�()Im�� �Uۀ �\̴h+Z�ر�Y��F��!���B�� �5�F�[�IL�J ���Es3f�e�� ����2�����m�B�� 5a ���m�5�@H(&��٨)e1�b2�
AB��M2��d*�T
Z��U%k+(�UƴЩ	�X�6�*6�j-jbU!U%(+�#\P�Mh4�35f��ֶ���al5�ִi��R�f���e�UTD�KngY��k*VƲ�R��ɬ�,m�٬��X*�jR���jP��U(�*�Fۀ���d 6�l ��6� 1(M�����X�T"�-�Vي�)��	��X  ��64$�MJ��
Mm h�� �4*��P��(%HA� #� U,��Հ(-f��fŔ��� 6�Q�mm4�ES64 6�
��[���VZ�+m�l�B�ن@�l�i3k-d�U�# ;�  �  �  5= �JRj���@MF&�@ EO�0�T��0d2i�L`��)&M'�M���~�R?Jd��hA�OS��)*�       4d���`F�b0L�`��T!ML��L'��=OHb0M =F��Ïӕ^�N�%�T�[R��Ү�u
�O�M&sQE 7��h�� ;�U@	�C�UE���e�%�`��G�A�>��B$
 QEgI���*����$��R�U����p"*+h��m�5�F">]���L�E�@]�q8�0
�H�r�w��Q.�KU9�;bd��E%)�I�{�ۯv����J�!Bz?��F���W���(}	�]�_{/A�}��A�/�U�K�:��!H�4��x����Y�H$�Z��q)�$�W����G>�>�ѽ��}������Y�Vp�C�m��v�5���S�R\k쪓�U�5?�u�%eF0k$@`���ZҀտ��I���u1�j��]�VӶG����椱���
P�dF	w'M�S�v�*Ib:�/�5��L��V2ɢK�DR%$�{w*��sLӥ:#)�R�Eub�Uڌ�tSR^��2�:[�%��n���v���[ut�3�Q�Kj�4,�L���-�4�����7q~|@.o' �}Q��n�/04�6�V	Ԟ�F70���l���EI�:�lA�5��s1�Z��D���)�ի	�d�9MlY����2�IR���&f�[��Um5Z7Fȭ�� FV�u-��h3At�85�Uo��誮5��A/���� ��L8Ջա�sd�h�����!���GK"̥�:�V�a���
QW$w��(%�q��w�bf�kgt�l�QT�mU)Q1�y��ķ\½�����ea��m�ypM���R;�	�ٍ\��O'�۸n�`*����H��vظ�I�0��h��4誻��MC
M<�h�����ȭ^K9�)x°�S��K��#��&�Lx/-a4s+!����kw[������:#o�f �ȄVRՁ�����/NC��㶎��43�����`@S����E1���[�P8�4�^H��i)��^[򘚎���S̸���"Z2�u��7�Uz�ƯJF�ؑ=�C����4^����I�6=�ȳVQ����,~a��v�dH	Q�fҧ��0�ƶ��I{�������$݌Pi��N�����jƬY�jf�A݇��:M6T!c'im����7{�]�VXݕUa�I�GJ�2���[xkvFE^Ѕ�Su�!�FV֦Qof�JX�j)dFe]�Yu0l��2�Vn��j^��o\�f^~/,��$�fk+M�ݗ���hG(UnQ������˷*��B�j-��C6v
�ݺ�Dzd?١�5Q՚QǃU�%$�l�vp-e��p��7���͖A��[�����ȥ�hn�r�k�^�2��<9��h��X&�附���+Un��ȁ���t&�B�jYW�8�2���\�XB�����W�x������:�l�����R�6�q�
N��6N٢gR�-�÷� �EՌ6���V�)���ƴwe�	��3.�邞1)�Pj��B#i+-��.'��X�1�v�����$t�j��rѢ�S�b�5*�
]����l�d��SC�Ƕ��&i�7�lwJ�{Tت4�˿�5�3I�ok4��M��t��P�ƪ�T�,��t��N�U�UYV�0�Ҏ�a��u�mPvCm���xt��\�y�Z�1�oE@�����7.�+0\'�6���3CI!"s7.��f�a'F����S&�j��v���2����U�%іYw��)��ND�<֮�ke���u 
�!VZ�����v,�DU��ŦX�*��ۙJ^(0�����*�v��Kgu%7�5�÷�Sw &靂i��'SFGh�(�ǹa��t��
ф�Fj�-��v)C7t���41OjB#W	�ɸmi��T[fc����H��",�Q�h���L����i-b�ƈ�NM���N5��Gf���'�ǚi���lH�;�.aw�;J�Ŋ���h��ޅy���H��0X����-�p<���茂��vV������E��dÂ��	�X��J���nT2�m���wt�*�U�9w&S��d62�X6^b�Px� ��b�W#Q	�){��RՠɈ��Ӭ���S�Aj��/Yљ`�q��/mKD� X�����FՌ��Q����X���z�]�hWA��,ڗ���A9�E�Zr����3d����ǖ�f"����%&�jiR�Ɣ�fb�\�Ӡ�e����buTs��:8�P�-\�e�F-`b���VhQʗwz�D\�oUң��
fi��.��w�J@p��ǔ)�淲n �ݣ������n�܍��c��I�+�銯Y(�($/ �l5r>�T���+H�wq��3pCV�I{I�U<hDҷ��,XX�[���B#�:ܭ�3~T�U ش#Y��e!�j�7#N7#�	���g(K����KB������p<���YR�S"\[2��۷,K����u��e�r���AńEOq�ܓU�1�;��KEYAB�"�X̫6�lj�R-Q��ޛ؋��4�0Vk:��Cd�j5�,
ĦE�-��)�ˢ�T�+v�	h�X �GP�0�����;`�T�4��sC,�mHn֢�M���`Ul]�*��MQqA3��97 �4�y��Ń�װV5�R-]#���S��M"ә���S&Lpf���1��c���M"���Y�a�_5r�A[��Ug�}Ǆ3U��D���
����mTE�y��ə�@c�.EyX�K�2�uV�$��&�I'!�,�U���h��ĝb/ڈ�ss7\�hA�&��LX��:J�md!S��轣��\ˁ	L���3�����+�'�F��x��lͥ��dCC��&�ي���j%fo�2�%l=�,q4i�gN�e'�F2�Q�9�]EX9*"�*���d��^�CY�tPG+r���;'h˭{B@ke�̫h(�H�`����U��e	U1�p�/E兰ɬ��PPU�8��ܩ�M`ۈ�B`�!`���O��VPʶxU`_�%[�PB�^��vku�����I"b#ٛK]��yl9u�A�R��TM�m�V�ۍ�z�Ie���R�Sk`����2�P���m�1���)�X��lT�#����f�C���.�[p��NƝo3͆�ws�/�JܽMd�9�a����d�S�'5���j��Z��bi�mm+�pƶ�Ц#������J�גm����Y�2H��`DЦáj�Q�&���]�9� -%�Ɇ�{����U��"ͥ�3�dme*�ǮU���i��P��+fѨ�݊�@��FJa�]k̼�Z�[�1C��n����F�[�Z���!�L�D\�mS����	bV�;�Y�AcN��)��wvŜ�X(��,w1�&��5{�1�V�������48���D�ڨ�a&�8���Y]�^j;��K��f�����)ۦ���d5�5�aE�����j2�Ol�]D�d�v�����x�M�/((�4dTJ���Mn��h��P�@���@eb����v,���u�h�[j����[nQѸ�H�{���+�a��a��O�7�he�A ��M:��۱�F��1�[�xJ)��AIe�wp�v��v��V�^����9��Ә\�O���.�0�܆�6I���3j3@F�jAEV�n���MGz�m�WP��
�P�,�r����ʚJ/ecFE���B`����tR�Ǳ�Yu���R�q�zJ�V�J��YW1�ܐ�,�T�6n�P�,��f�M֩�ݼۄ�u\�(.�7��ӡ���q��S��ʵR��3 hީwF	�&)d��9����j���r�1ԶMl��6
��;��[e���[��l��)C[y�SA�ob��
�����(�X,��ʋYٙ1i�(�t%RU�����I�!+XR�5���4�*R�C�0� ډ��5V^��1I�/�E���N��DJYG�}	�	����~��@_g����o�:;ۂ 7`='�7�F7����wc��uq��Hu�#c�m�4z4!hƓB��&�`��^�آ}>����Ov:�{:�I�Кu�I�?}�oc��q�>�F�:ݽt��=�w�{z&JMQ]������
(~�����)���i���H.�:\,.Y}.��q��K�ݖ3jѢ�3�P'2�%�8D�N1����Q:k��Ԯ���ۆY��yAⷩ%��, {��*��N�Ɨ�V�o�Pt��].j�uN����M�Xŋ�������_[�l<�>��z��-X����v�̙c�w�"/g	H�<�s/tTꜸ�e�#�ϵƖoL�=?��5�{xf�Z�ɯ+�,���.�f��3+"Y�&�G�1����_8��k��e�[��7�־<��XHq���kB�q��"<�;X����}���a< �K���[�z-
�vP�^����AN'(L�zL��Y�d�w̚��u�{�E��o��6m)�Ƥ��cj�ʓ��Y{�9m"Q�|�%��p-RF벳����9-s�ɳ���yp���-�G��9���4cW��5e�}����Gs.�#�n�&%fq��Q2�,x{׮��\�Tĸ��`];(�\��y�=�P]M��EWI�`ɯ-���v�󛒕�����)v��B�Ӵ�ܵ4Lq���;��b���.���ε�d�.%֋U����Q��$����[:.�fk}$
�W��x��U�i��G>b���)��k2�F������݁���8ˇ��k0�v��b��d����K����w��0�A�
v��SxxǺV�BVT�Enu^��>T�uˢ;7�į�F����;u�0MY�����
"��1r%�DS�f�n��iQU�FȪ��ow�����?ejy��L� �
�̐]�c��f�!��XD�(Q���g>(Zʲ]�ݎ�㹕�f��ҵnr�w��s��{�L:����9�n��ks�e^�;���b�-�:f/�-�ǉ�o�n�t3. tI��S:]i�,�M�к���Z��sܾU6�wX#��ε�\妸8�e����
���]���I�3R\W�6��?]�N<���r�����gg?K!��LR�\M�T�)�
�j���y����^>�D�z��~��j�z�ˤ��4�M�����,��nup��R���o^er���\�'b:dh���	ٺ�Ӣ΃d��0�q���W����eP�ݶ����.j�ꪁX�2�� ��;bn�- ����.q�'sHQ����a�ёM��u
��a��M,��Φ�{ox���-L�A�ڻ �<�ϻbcF
��u�:+'�{������:�כ��6�u���I;�&�1��@�Lu�Vm\黢�GV�H�nr��]��fse�=��9�N�#u���1K�X*�R�0W]VP�h(+z9>�z�$ZL���)����K��f�r�z�.T³D
o�+c{�>l�%�	�M�"�:#¯�:M-�/,�Ὣ��z��Ya3��=+j7i!���Gt�Uҡ�cul����������Ӧ��2������ۆ�\`�U20�+4w8�OX�!��{���/��&������;"��sK���>�mW3�(�(X&���bV��%Z�x�xJz΢��gA�UE`]3���9=B7�X�U!�d[n�cNb�l�WU�$�|{/��Y��B\:oY��S%ۣϻWs�;Cik������姢��u��sT�Uۭ��u��ǂ!mSK/�s����6V�M[,��O���9F��%w=ԩ�(mu��5ئD�&)����"l�1��r�"��K�G��f��[�c%.H"�A�n�$93y���@�=�"��\Dpyx]Nja�%=[��݅ViV�����؝���;�`�AҤ�-�9(+��nu��ɯ���B�{!���M�௶��nK��CU�'Hz�]t/^p�m�f�7�A6j.�-�B�.Ei�W*
*I�lE��J��;���=ֺ��+�[NH�*�؍�[�F��-�Yu��OxQ9(��ٗ��W*��c�ة���SZn-�Dv�'=�]]V�q�h���xj�mh���i_SC��؃��k�u�.(�U�8�f`J�K����d��A�$���6�P����Zu�d�m�'f����:3��ݐ�I�4>z���CJ��@0k�:Z�)%����FK��v�1���ܒ��l�<����{EI�W=��JmX �/T٣�&v�[�vȭ����fy�*�;\q٭l9��:+zl��W.��Sr�!�V���`��Br.Hw
��Ѻ�Br��޼�D�8¡��֘6����hY����%*�]�����2� iM�7_(�W��S)��[��-+�_����竴�jZ��:䂎8�u
�H.����=�f[l�c̖Ha��t��އx�QPgK�ԟ��EE���[�2RZ�r��x��#x,[>V{�R_��	}g�o�u����3'�+����W�v"Y��ʵ�.���t�ҰA7������wsDq�J��C�3A�K�h�--�'��e��V�%�1�7�ftcx��I��,�ʝ�2uC]�X;r`���>�8ұ��u�ڈ�&yl����IW�N�ൎ���Sh�)�f��+4�S�=O�xOC�j�y6���n{�k9�1��-#���7yl���i����4sM�GA����tmq�;I��ێr;K�L*L�e�@���r�`���u�[����/��l�ɡP#yT�o�Y����m�DH,;$�ڮ�K�:ڭW])aQe���h�J)�e��2��-_A�YU�GQ#l�tjd��%�E�ԎV9C)����X{��vt5_�w+�ԬA��.;�Y�4�GE��]��`hN�˕���W�2���
2�n=\@�w�쇪WQ���F���vk|���qw5kU�N��mWJ�s�x�]���r���'�.��4�mq�l3@���j�ӹ���j�gä㢭d�ԎN��WR�/��%����+	���/	v��]��6�`��t���Z@�ܷ�L��1w�Y��Vܮ�f�����I!�Y��a��;5�F����`pL:�M�U7�oL��>�7:�/���:��kr��}�5D���6r�N�S���5@q)*�s�aL�9�0�wWyo��Τw\y�L<�=#�Fr�����|�-�����v��*x�gk�ʭ���0*�]g�%��9����vU�}���<IY(C²�RI,��I$�I$�I$�I$�I$�I$�I$�I$�I$�I*Y�$�V$�%RĕLN$�I+ĞҼJ��,I$����6�	x�f]|�;�7/�ӕ��4Keˬ��q�)V���bga�\��4;v�=Nk}�5��9|NuwPZ��ĳ����4��t������t��35�7��Ss��r<Y� ��{xM��۾W�]����EA����ᄬ3�9ٹBs�]3�e��ޅ۪d����^�+2�N�`,����wJ;���!Y��Gr�U!�����\2�&���v-��|�G�֍��8�����<�V�1�36ci���*(�`+[�`aV�2�����É,4�2~�������,U��U(~������J�=If�nǚ��o�r�YJ��o.��0	�(=5v��Фf�q�`���U�+.��D�ܧd�Ę�1f�9�Pt�J�o[��oq�#�9�H�6+VU�^Y؝`�/7B�u�LTh��e�-8Yb�U���!`�0S���Ĭ=N��d�2���$����J`�AYkre
�#�$�*���Xu^�}_��PT6]Y���2;��(��A�����3{�<���D}_�ы�jq���W4�W#���b�u�g�퍼� ��<����.v`|:pͽY���(k�5��)%�a����V#}W��O϶g�X2�P���Z��$���q�;e�Va�Z��`2��Vqirؚ�fb����RݙE'��0���\�D3j���!�\���9օt\��<���8&f���7�Ue���*5�n���2*^�v^�rv�)��gC ��ۺ��+)iR?����v}��=�f̔/6S*�)q�7�\����&u�49���.)bY�̲�Јmށ���ǵ������3��=@M;J�Vj�:qw��{�&��h`W׊��]a�jn�S�v�fhV:�+h�c��1 {E�{s(�l�\�{o��9b}1���{�x���n7|��4�2��%���sn��C�V�}b��4��/�U��d5�͝�gh����S&���Vۺ�wcqJ�b�N�؞��qG5��w��R���TN��`�Q w�x!:!lk���e�e�6{s�ʖS��&�g×{D=ެ�]wL���z7#��R�ư��׽�T{ꭦ�� ���Y������CP�&s�X"\�o�Zm�[�'0�Wi]�i�x�`y�����_D2H+M����m�oV���*�P;�{�;����a��NS�ֶh]�D�jlޜ��RL�e�
vu`�����v}�4�ճc9�!_:��)�M�h��}U�la���͗�γ���?&�'.b#5gg�w9e:E��۫v�wWW(B��5�*f��v��z�\���m��Hܚ3���'���R��]+Kt��ox�q�,l���E�h�\���@��������d��pb���`B	?�v�BBG*Q��G,��O�M ����7���PD�8!�]�7zI/9u��۩̞厗�Bu�g������U��&�Xf�\�)�Ő����ǔWRgj��?9�k���pu�F�4D�ӄ�Z;���K8�_c�n�l����IaP~oRN~��ŌU�M����ek��.&���o�f�W�E-�Ev�Z�[��Qv����FT��\�Od��;9��	��h�o>��}����_L�,m��#N�跧,o'Q��{�v]�XWd��Q�Zr`ү��m�#V�Ʌޠ��2��Ec�]��N�ݡt�X�)��1]�=�'V��tv���BRE���)��]I)U��*�$*��v��3y�3��D�j�ٌ՝���q�r٭?�G���%�V�S�&s�[Ůs�2�Σ��#x�e�ֈ�i��Fڬ@��9Ŵ-�8X�n�,|Id��h��J ;��ai��֓��]l$����Ikt#��R�ˡî�q�=��|�@���Eu�n7dκ?�2�O�7�)�:o��m+g��7G�4�eJ'+���p�a�D�>�Oc�a�����GW7(���a�]5���SB��yZ���e��	�F���Ve����=aUA�j���Y �B���� u5�],ŻZ`�t*�\���56*��=h��	l��L��Wջݣygۼ�I+i����tfq��7f����T��hX��@��K����z�,gk�*(�L�n۫��n�h�\N�v�]����B�����C.���_�q@%�����%Soe����ܯ��{�^v��ⱽS��g��T[`1��]��5��_m�}b�q��ꬫ�|M��O�t
�rړպ4۩ֺ)�&Pp��j[$i�Cz�1Z����o�U�h#G�yf��=�-��BHSO�Of���}B���- �N���1�xX	�[�6 UJ��Bl����R|�Y�T������*��L ��$N�T�/�7)B�Z�����)�yyGXδ(�7��tjn����5]��sK��'uS�=������7Q���۶�S_���y��T���p����}�=�iV�#}݂���q|!��@swq�{��$�5>�^aֺ� 2�	G��j��� ��� D�NAS�<��FW�y�1d׼-���@p���uJ�#�	E���{ ;3s�17F�|�v�l�NmR�ݵ�S�����D>["-��-�i��u79�p�<^#��X��[�����^i%��B��-f�4{.�#p��I�<��p��@>Ԃ�P͂�ъ��^󪢬��.$��R�}W>�V+�_!-Z��}&(.i��K�;\�Qf��̮Xh�}������Y����]�*�#�R.ŋ��i��cY�0+�4���+��Щ]|�,y@8�S�����jc�[-��Z�rT%�Յ1��&�ܸ8�&��Z��"ڳ��W�U�0P+�\�Mf*sb�]ޱҵ��{^�J�������F��gM#fg�vՋ��א���Vkf�[d~���k0	�:��e$1����vv��a��ưh�֢2�� �g��כ�T�(�%Ry�¹b��a��O�f�c���B^tH���Z���yAJw�&|+���}z�7�Q��G��-E qoo>��G�'�!��C�޹��Y0?���O�Ӥ�;6WԵ<](ڏ*[�úP���K�(F����$?)\&�P�FzS������[��mb�!�����"��R-�Rv{����t" >d�G�tT"�`>�Xө���>Q�u1��6vW��pA�Y`�J��c�:�WJώY6ie��� �:I�K7�	5̛ߎ;]���}��<Y�:�K	��W8�W�w���U�v>ܘ���>���U��z��W�g�jK��K]n�	n���ask�jUv/��(�ttM�`�%t� �M� ���V*�@�Ll]e�pC5��������h�۠�J˯��`�� �rY�:m�����N�j��hˋV �ek ��_�ц�44�'W���V^�T�\����HX]d;�nv��e�J],/�h;��N�f�왗�*���2��U���$G���J{/���*磺�0�'�;t9�����ܼTFF�b��JJ�0@�d��k�j/�`�['w~��:E�e��j�C��9OR�Tz`��W˵f��λ����OVe��`Z���v��uH�\F̽sp;a���\�[�ٗ�Gm�C�
Z��"'g0���t�^�G���o^l׊#���;
��xX.^u��K3&�2٬�������	Ar�r䣉��뻻C��fu��m>�5�6�GeU�F�;�ݺ �ٻ����{�ڱ�,��n���&�����z���
$S��V9T*��.�Ӫ�l��o�G�d$R�fU|�U���o�TN�1*�-2���]:iq+4�.kÓiy���L�{����yb�*%}e|�y��y
f	sI��f�
���	�˿s4.]C�}k9�q/�f���"8n�#���N�Վq�Dջ}�o]]�p�]fzC|N���P�U����*�D��j��P��i'@FP�x���sƶ\yZ\�)�xn[��@iy��-&szX���;w'`�i�]ֶ�F�ɢv�(Fr����(;�]f�v���Իm�d�xNU��Ju�b��.�ˤ�7k�����D��_Wt�٦Ԩ����<&�u�Q��@������zA���;3pk��y�ǘz٭��Di&%Zy���G�l�:�����%���q�Έ�*�9��n�f!y�"Ƃ
�M�V6��Ȱ^L���8�Ef�}xf�7��n�Y��������U�K<w�e/*�b�N������N]k��i�w��Wq�b�\Afɑ�#��[|��]�gt�� �����E-G�����P`_��4�����08؆�2���	�)�DQM��g肈�#MG"j(�DDp!>F�q(�m��2}�"f$B�A%i�C%��)D�#o�`i(`E�-���_0�0\��0�L��F6�O�ą Ԁ����غ��`��"��8���M�'ѵ��q�b&�M�R�#A�
���P(܈��" �b"�+�⑐JF�)!�H5*$��6Y��~M�D% q��H�-�\%6 ��P��@/装H����
��DU�����>�Ϋ,xr\6C��3C�M4�S����Oܖr�X����Vvܭ�m��b�`�xq�i� �֢XY=�J�X0�-M���3E�h�#U����7i�5f�eb�V�lv���OYt�F,�����h�?Tde%X��5��{/Y�Z�!���Q�bVk[��Wʴ��NDM"zL��M��k2���P1�6�pLr�F������S��ӑ��4l��ZEf��FK��7�^Y�ί.\�zqR4^kfY�j2���Fsx�I$�I%�R�̣�����陌ܚc�N߮�*��W�^�c]�~w��x�K��>����m��.Ƿ]}�ޠ����A~�E��8����]�[�s���h�*�m�QN��N�"m}�U���X1jϻu;]wDΒ��w�>����!ӣ�n����]t��m�J�����wn��tBoYJ�T�%��i�ӡ(��'��7`=!�q��@�����4h�u��[&��:)v='@ztm��d۸4���M.����� �7d(1X���D�l-��@m����1]� Rh:Āi=��;`��g�l�F�A��G�٢���Ob�P����Q?q�~��DR]�N��j���{��tz�{n�c�M�������h�ԟ�ރ�>���������U�E�҉I?L*��>�5�Z��(�,�d�-�1�Q��1������,�A	F `(� ���)��:��Y�}tMM����>���vvk@�+�R��/̾}�j�b����"�$f7��瀐����kҮ��@�5.�l^��Θi�[�n�]jJT\+�p]�	�-�ڹ�[���o&�g���LnM�~����L�c�^�S��y]W'��D�Mn���8�uN;��v!t���=��s�� �*�:z���x,[���S��f���ʹ�!����</��3�v�wI/T��V��zD���I����wO}|V��[����]/aO��CV��t0	���E��z�b�@�B(�o��%�e���y*���୅�f����^����L�i�G=��;ͱ����o=����Oy�p�A㥒w']�2��nva��En��T�����oǎ�}�^~�:��x75����-.{�+��Xƿn�@��}�mV��溧`�ʠw_�UzOi����h���o�����#K�Y�߶�{�{��^��K�W{`g��]����'�����^>��+��\���� ˴"~Yma����:�ܜ
�0�r+"��H��m-Φ1��+u��t��+��k���e���5�Q�uf��Bwr���	�����4o |���tm��U��V�W.^ͽn�#[|[Ń=�;����o�^V�J���FSl���b9{:&rP�v���(4��f�)7k^��M┫T&�U�p� %��v�<P��)	H��(�m�F���	�*qN��Yd�Nw�6%�ZT
m3����ȩ�UJt(�W�c#'�i��(��׺����{؞�Kй0_t��&ߧ�eWz�Т�3���m\�RoV,�`������[22u�k���$N�{E,�����+�y���}��Ta���2}�k�J+��[j�r?M�߄~�KوD�+���ڝ%�g	21JT���^ay2c�V�Q�{ky�y��<D�}�(��h�5�y�X��sMh�SF��s�޻��:]K�:r��0��fQ�z��F>�Ûsp.�ܨ26��xJ���7����\4��G>u�5�'��{ZM�'{�YSg�|��B��Ɩ1e��R�{��^���������g�����&�a�26�,��H¦���^���+��&�M�VoWW�t�x�z���TT���ޘ�wLn�{=+��Kk�Ox�-<N!���X�g�Kǅ���Sx�.�*^��Ǣ!�Rļ�<@���=/�^~����u�C�f��,��r�g��g�y��Vނ���Q�vr����۬ӥ�I��ڞ���k�.�ȟ���D�JW� �V��m%��Y�5|�!�v�WA5]���EC&n�Hd�'[u��V�HC�{K���Q���e֣�4��+0c� �[EM9y�Xs�o�ұ����H�ڝMT��ͯ{��]�Wh~�>ǔ����J��^.�[=�=�w]�����i��	�[���W�S�w��xz��ͥ���%r��R��P�3"�ޭ�ֲ���j�{�����v/9J��EϹUW��eW��.΋ʲ�D���H�,Q�)2�u�N#)�洬t���%��ﯗ��=�J�Ϋ��#GC��F4m���l$�J�n���L+�cj��m��$f��U�=#tJ !��Qb��-������QR"��<6�6�S4�g;%�"���kq�6v���s]����7y.X���Vq���/��m#�)x3(�z�q�O*��3]bz�J����Ϩ���6���8?:Ǖ	U6m�ǖޛ]��9�^_'���x�{�W3��\��٘}�Y���0��y&�*g\DK�;��N2RݙڡcNf{i�E��m�>��/w�Ky�³_en<��|N*?-�!�V7Oz�Լ��~�����.UFz?�{c�u���v����χ�v��
����mFC��'~��˷N����e���+����g�KG�G�p��q���M�����N�1��(���FʼaU{m���U^$G�(�7Q��K$y8������%2���w3[S�F����@����N�Њ�m�(N>%+[$�ܫ�yw�[�%�w���Ug��,����4��3?V�k=�Z�M���oA�s���M�{���^ڛ��E*�u�K>s�[~l~��HԤ*n�7YQBo���١����Z���l��TCc��>F��"^���
s��7��u	5�.��}�.�+}Ǒ���ݪR>�>^��Cg�hxh�k&�wb-��bǘ"����쾙sg�����1��nU+`K��΃}'�wS�oO�sNjoc�y�ė�vA���uj���ZC�r�ٚ��;:�.{���*��I�٩�jv-ԙ'�u�y��n�N_�ۏM�����h�(�w�N��oռ��R<�s�E~=7�q�V���J\�.��o�����ƿ�!嵐%�<}���j���!�x̭s+m���ٚ����\�9�������؃�C��^w�������m,��2��u%���^{Q�V��}��n*[��i��z3���-�L�q��~�p������+F��~tqc�7�0��e<C�:Y�w��P�6n]I�[y�|d�e3S4�?y�+�Ŝ�EEb8J�F_=s6H�MO��Kݙ%E���c8�WɵR�h���Ƃ�f��6��Db���me1w�;�/��D��w�PP���Dyf�nhb�kYkǅ?U��Gs}�8��ם��v��������i���m�eU��D^���06��%4�ؘ���Z�U+�-i�w��q��
9�l�V̞��1_'ݫ«�q�x(��"b�3�0Os�L���c���Y�pI��6;�S����aS;I��ϔ�T�)��,k�dQǚ�xTիa�<=s��U����:V?W<����D�~^�~$�j~��N�ž�o�.bN|��%�&R������5yׯ7�.��̾m�q糠J�`��x��#y�б�Y��Tt!��8�5I��v����;��z�Cu��j�7�ڧ7Ue&�uir˨ūf�r�Ζ��q"��2�7F�yQ~�ʹ]�s��1A�av�y�����Z��+�{�U.�rJފ��	�~�0-~�wyS��g�/j/ngz!W�?_\���WIc��w��[-w��n�^{�tT:$�me�ט�MN�e�.{φ{G~
x^ט��{��_���Uө�q{|bU|+:3�׫��sT׎fOll�K�=����T�-ʏx��j�
;A�ξ�1�O�#��N�ܰ���NY��~�^�ϳ�H�]����_�lW��<&�����0 #�����;�@��%�e����»�Ss��(U�_�,�P43�\����m����ޭ��-7*ɛ�_쉚�d]�qmb߱��N�N�Ot�x`2f"�5�AÞ�%�˨%A����#g.�|»��(����{�X�O>�^fX�u�'Z�����'-����K��\�9�j��L�������2��g����:;ۻ��hV
��eAы[Ai���a�uo�I'oxe@Z C�l�]�$�$3&���*��J�m�r����YقxW���dom\�"�ZMUV�&�Zv-�-7�Y%�kn�!D����7j�u��,8���[Ǳä#n䕬KR�&�7@����+�T4I+�7�:]s��ɶ�S�U��Q˦���h�o2��^+;K�D�@��W˦^��޶Ȝt�y������X�]fpeSz.�2�p�e�k9S�jJ��o;F�;.�5���^���K���&(�F����H����u{�'���v�����T�V����Qj�C��	�E�]	W��au��p'lP(��wT)f��ҰU��(�׹��QԋZ@��.mN�(c��}V�!հ��-� o)yŎ�v�r.�b�ŉ���F�X�J��5�e�j�����ݜ�o�Wr��ܥ���M��q��5&����k���L7�Y�l���"�>f����CV����x�����yܛ�aS;[��s���m&sst/���M�-&'ݣE| 緂K�d櫃��dw�|z�X�a��LEU.Q��ӈ�zĒI$�K�P��+������Q��UP������?�;t���&�T�ma���ö8s~�PB�U����~AA �@�	 ���E1I�G�v� �l∌C���F
��8��ol��:�h���G�1z�%m�稪���W��w�uRUDU���`���C���=8���(bz�݀�f*���t���>�h��}���r�Ӕ��5E;��-�M�����f�EQ\�������s_b'2Vh"&j���2r}���ˬW������& �nZ�5��;:�?Lԅ��j������guP=�jn֢�>�w+�I����\����V�jN�/�X�o��!�e�^��в��/��u���'-]�aw��0���r	�����t<o�a}�<��-'���ћy��tb��k�=�N@�|�M��M����+x�~��4}k�,�j��g	��d�Ga�\uk��|�tjD��x��9-}�}�Y�#���q�.�[@i�khdүD�4x��C��U�Vh�ay����/9ԧc����c������+8���v�
�m�`���0z`lil F�;h�YW{�q]Q�����Yw�/.Me�9wQ;�Utfk�b�㖗$/���TZ]��
��2�+.�s������xN"���`>ᗋ�52�w�1�����m6��|��aN���{Y?c���տ�t���W5�Ҿ�#��=�?���A�՟���h����*Z��+'��մ)\ck��$۾�[U<fθ�����s���7E|��G�~+kt�^��?�/�Sޓ�љQ7�ܓ���"���g������Ny�곽�y��7��~�s��r�A@n�E��z+��g�A��j_�Q�a�N�}hGV2��۬�������J�I�N���+T��(Z�����M������;������wV�GA�n�M�A��A&Wu�%-ߪJyVW�Χ��郺�#23���uB��W�M����#e�ú3:�Uݹ�uL=S�M�cs2�X͂�� �9:.W+����_������ćL���L:q�rm�!�׬�O:�{��k��7;r�׺��ʎ���ޑ���4���SՂ4��gt�����}ޖ�n�2�&��n�v��y���	ǥP�7)�]n�U.�h�Z���ۼ��馪m�4\��gu�c؍��Ճ$��US}�W��R�[�q��������K�~�I��] e�W���r�.؝B{�*�����������E�S���.�!���w5GK�|�RZ�\�Eb���OԆ��n?�}y��o�L�a{�~��$�irK3���I��\��
-�v��{��P��&pͨ[�������sdˆEv�R-9o�9��*��g+���/�T:T1q��0��`�9�l��;�c2Xh魵��i�KT7%_���_h������Ѧ#��'M�F--�S��/��u���.ψ�Z�Yݻ7����V�_�2�!��֝���\C�^�VA9;m����7MD�7X�g��^�CN��W��3�11Ҳ��&�[֙�<��T��Cf���
�|�
$�����6��ո~T��3D�=ɥx�
@�B�~;�Y�OMf%��	d��g4�'�eN��?�5>}b�X�q��:{I��z'��y/�S���H�ӆ�i.�Cc��շj)]�����c	SYM���q���iz:�b��l=�u�\�~z�nIt�w�������ρ}����[3�����e��.��I67\�yՄ'ٴ��kI��}����թ㢣un9����4d������b���G�}&{[�[(Tb�}�w�f�Q?|H���ʷ�s���`狀Jco�-O+��N���N��e�>� V���g~��s�du�+��\���!YX�}B������9i.~_��J6mE8��mu�=����Sy�9=��1�����,�k�P�}̅:�4�q{�q��f�u�a0��Y�h���~a�ݮ�����<6��1�Z�l{�������r�ʍ{�:�I;�6��N������L8�]��9��;����kgr�� H��<�r��kdwj��|����gC8�j0`��n<�
��}��-e}'���:ok�	�����G���6������7޺�ݕ<�[����m�uro$�%2,[�:�x���x��C�<�a�.6������+�틽�8�{R�n;��wJyM��ǲ�S�����[�z%����:pH��S���]�Bg�߽����,�S�m{`S3?|��^�ڒ0�C�SܒҪ̺l{Z����)��i�v�~/9���bG��v_:�1��I]�κ��'$�W��Q���,�����Ǽ������R+��c�9�Q�sr�m��۽�蚜~������/}IU�K�=ޔ��[��s�^&矜WGcT�?���yu]''ΐ3����R�Ϝ��|35u�|��wr_{�w��eV�K�z�8�	i;R��?o7��-{�rK[r�,f	�b(�x[zvk��ѫ���>1̅�g�k�l�MoY�JrON�M��u:b�(�p�EDu_H�"�U��_.|�u5X�4]l��].������9����������z�W���ѫ�b7�ы�Gaک�ޭ:�)c#�d9fR��1l��t��>���@�޶�f�X&�rZ	+�1�p3	�R��]����E��JZ{�~�Vv���fX;�vOF� �{�?��Lc5\��C߯������4��ܤ�[*b����pa�Qq��F�ŉ�ה�8k��,��N�%o8�����nk�\h���W��]p���}~�UO�����}v˱P�f��	}���ҠSh��@��&��?/�g���`V�?��}�ڳpe��Z��_�¸I�D~Z/����o�b�CjR*�ڞ-[^�ڇ�70�[�9����qp�Z�zV��͊��,ܴb�17�8�7�����%�c:B�
�7�U:��Ow
awE�����[��K�3�n�`��1�E'.u���1O3%��5ܱ���tW�U�vO�M��W&�e�\�$������/�z�7�`�Y����F��܆��������t!1�p�����_:,P�*����MQ��D�4��CɨCaL,�C���j��{��v��Ͳ���eBj�id_�b�iЋ� �p��A����y�є��Ţ���&)��8�[5�V�T7���EJ��Q�]{�+^���z���^{:��h�W���#Lh�|��u��y{�(0v��Q�5;�ܻ�oA�d�C��<1遹ʩ��>�z%����Ǻtˢ�+����h�3ͣ{�U�ٚ!�LcJZ�	c2j�dc,Բ"��Z��+��b6�k]a�x�l$�����|.�vŕ���WZ
�%#���T���#��,�¡}��v�35��N�����g�*�RV�S�]N
Oj�q�v�ٸ"��:&{6�a��<�4Ln�m�<���WO;];�%򵖨R�o=)f%d[��o[퇸��� Vm��)�7�ȞF^���v)gF����(��uk4+wd��&���ly�kk�ћ�p\$�b��c�D&��A�ٛ���\*�B�����s�z��E�r�ǜ�<g�P|���04ΰ��ͅ��7n�uQ�Kp��1O�|}fE\�}y����F�|��)�ZL�$I ��|�~!]���[M߄�=2]JŦX�
J�Z(�a��|��F�
�o��s�f"G��Y"���v�OE
\k�D�PN���K���� :M*OfX#y釥��G�Yj�-c�/���Ĭ˗�	eE�gnؗ�Ū�P�[�g&��ޏ���U[2ޝ�z�p��빪�Άw���O���[��J��^�i�9ooK��"��!ڮ�]|�!1A��*�\�adƃ���P���-�j�7ա����V�Rb
2�b��q�J&��
6�s<���9�{�X�� 2�b��˵�И��ے�|M⺬j��%�0I��Ǚ����ի�r�{a.l�[{'֗V����<P��3�ϲ�
4�a�]�O	�zeէ����N�,Ug;�ڕVK[�.�u7a��S;sw�����~^A�W̜���v�{{~�v��v�6��u��(�N8����	�Z��K�rő���-U�65����Å3�ਬ,��&���X"Z�.���bh�H	�۷���o[�ۤ��6��&�N�n\�E�|��V{�R;�:�̥�����Ӿ�֠ZVuȈCy�ݲNn�����@����Ӕ����[�W7QV6���Ьݢ�hg>������-���o,����#bq��&X�������D#C�.e ����[`6.�T�f*���-®�' 5�ԉD(]/��%e䤐x����\�X��' q��mM�Cf_�u0⪙��	�I,I$�I$��+J���Q��]n㓫��/��
���3ʨIb�!�+���Y��x�����}QG�((��b�"��iJ

�����RѶ}h�
i�hJ(
�=����ѯZ���QkF�ti�.�A뢨ZN�j��b�h��C��z"C�_N���	�F��UwpQG�u�dк4�ON��f�ס@]�4��s�Ђ���b|���	�$B\P҉B�ɑ#1�"He2(E)��R@RM~6�~��b�J��Tu|� V;�#�N�Zt�A�u_��| �������(��&�+�fa����nSY�m�0� 	�C�YPE^��6�nLNuv@�-�b��^Ƿ�)'B�*�l������B��l����^��0,Y�oN�m��y��r����7�Kq�J_w���[#�|��_}an"��d�]u�8]�5^�"K��=�W�]��US����WO�|���U�Tl�5��s(E�pm�Ws���6gxET�#y��T�l���{��3��Fi��"D�s����PY8r�]�y|d�[rr�:�{��ϾO�´�&8<�:��Q-�:�3#'�v+������/��TK�k%= ��� ��d�{�¼�I�)F7��{�+�&��N4,� ]Y8��XX>��<!�{Jާ�죓��K��摯�N��;S�ٔ���5�+o;iߙB���ݭ�����i�
��k%\Т�Gl8�哓.hSdD�d�))ډހ���a�h��Z������ɹ߼�}�����%=Lk��yo
_;`Ż��F�l�(>���"�:X�#",�(ng�}޼/
4l0bv��0����"�,.�j�tgZ��=��n�E�ڻ�E���={=��2�����k[N{tb��c)�q�_�;Y��UP��Ѹ(X�)��`qҺ�v#\2ʗ�䳫,b�4�^M�Ӯ�7�-bw��P�&���Q��^�W$J?/�   f�ժ{/�]|ϸ���)�.`��9����Q�c��|\j1��b�Y(�����m��x[��i��z�x�
/��+�����oFf����O�1u�'�wEꎞE��U�}��q%�x9J�������Ȼwe���4�Ѽ����CL�W���g�>D 7e{�����Fv�����Jb�ita�����:7z�nk�|m��~����.��`��w��qo=���՛����Y�yR{�~U����2�QV�72� � ��m6q����v��\CVu���%]Z���2'���:���;��[�h�2��Wz]ډc���aH�V�9�e�T$���� �Eݣ������|W�f�pO�o�ͼC/�>����R�ޞ�q�"����sFjc��t������6�wڽ=��]�#�4�[����V�S"��¶�^X��]�83���\�KR��jN�?U�e	@L����d��K�����]�e8R!�3:2����&�B'�7q(6z���F~��_-'�-n�\m`k�~l{�c��}�A;�U1��sheps5I�F��[�0��'�{�}L��[��67�<�nP�['��0�N�a�c�b-Z�E`Ҟ���xo�������8<0{��nP������WC����d�g���Zh�}&��WZ�n�z��  �1	F .,���Q��iT5g��q�u�d�?�ꚤ1��E��y���M��O[h�w��3�u�7m�lꕛ���b����ٻ����4싢G�#D�����_�^�3�p"�l��ҥ���Ն���Tf�RN�ͱh-��Mj�7��X��i�6��G�f'e���Ħ1��e
��(I��!�!v���h���xL3��s,���y��4 ��������#���wUZ��3t��q}�bf�����XcW*�z6�QЮR�D8qR������W������[���	��tNW=��P�˻���j̸�+zm�T&��
��BtR�����S59{V�Y����f]0C̭��V����E���a�6�J��}�e�T�r7u�3ݸ��8*][n
	��w�R�~��_��l�W���U� *n���u>�"�2�Q���/i3��0`ϴ�k3]��F�6ZHAݛ�T�����1ɼ�
T�c�����e�L�j(s/�n�e��*�~�		�n�ttGZfۖ�O�LF�+Q\A8�>��1�7�~
O3���C������{�ig�+���D6��T;��S{C�_̕�
e�l8�M�%M
�&���e\��$q�TS��hv��tf��&�׸��N�՜T��NN'9���U���i9G&�a����KVf���x{���{∞�ao�]�{yBqA=���P����}�]�sc��+����/����������~�~�b��*�ț����}�O$��mO�����*�q�}L��f��hT�|�T���^)�^�t�ь�^k���j��W��&�9N��Ke�νW�˸�7��Z5Umdn�4�:�^|8�B}\�V+���^�j�d��Y�k��ޓ���j6F7v���\hx��
}�e޴ʘn/�I����4ou�3��J}C{e�a�׷��<��;��4Y���ϻr�G;0n�p��8����r�0](C�����+	gq���У��gYE�^
h��Iy��S����� �D�Փާn�p3a�/��,4��>~��.�7.��0�j����;Wl�w]��El��6CE���p���v�z.*�����*���z����f�	>T6��S�}�����Qž���O��/�;�ï�}b6glQ�1�]Q#�ꗽ\� �_Z��_���z���4����S��H��p2.��a�o{��$n���ö����d���4\��V��j�ћ��z��Y�a�3^?y=�;�z�S}ٵ���":;9�Z�9��k��%��eV7?��Fh:��6դ�3���!���
���B���%=ۮ�����6�n���k!�wUA ��Y�C��P`�z,\���Uaa��xh��|�D.U�)�h�r����k��������ĩ������\;�;���j�����?3�h���ғ������[2�6�#v�fm�I���XJ+"���n�%����\��:���͘1�f�>!��Ӧ���aO�]�{���o��N������)�W|��pi����;䣪��12��vuܶ��UbN�S	yN��J�D[9���E���f�蓟Q�X�6���|_�l�9�T���̟^��߷X߻W�����ɰM+Iݰ���5���l}�t&q�~��Z�����w߻�O ^�e�3�Jp,
WvlOP����n!�f%�Y�����U]Zw�_�<����]3���S�@/�b�u�}s2��8h��wǂ���Iڝo��zg+�ѳ��>ڇ�k�ע��R�د!���Y:����yr�d�δza�u6ɩQt,&ܞ�X��9�����������D��6>��[���r����R{���H���Vc��.X]�L ��;8R���
���g)��:��٫�z��R���3{�f��E�;;ЀDx'�2��ˌF_K�[���z#�i=�U���|�('�&7� ^b�p�0�.D��6V�n)Lyeh���*zic!� R��z�k���@AYz�e�;i�����v���3[/��C�v���!^^��[�����iY��:��O3�ɠ7rr��*^��:�7h�a�s"�*��v�xN�V���W�t�5�݄���dY�w����Cn��ҺZ'd"��Q�f�t����tn^.F+&d�r$�q���j�Zӕ�QvY�9չK���n*a݇�}3���N㭷s;e�L\S�ORdV�i��sUt!�97f��S��������98-N`�Dme�]B�=��5���N�:e�S�Z�в�r�"�8��suG�;��UW�ա��3�����Z��(Q�=`��J]b��f��P��s�ef���]�[Y|d/{��������N*^S.���W����k��I�14;�ћK����QǶ�䃠�"�xM��ua�l���e@ċ���]�=þV)�	ݡ�`�P���g�]�n[�+uB�DS��T����n���'�������,�`�u�D�S��$�U��NM�0������r�4J����j��e�
��UCH����L��p�uC[�Y\�Q�����1( ,qXNR����2�ʩ!����uKM��x���x��6���v9���ĒI$�I;�T�ҨwNv�I�/t*2���{>�A?���Z�t��g�������>��H|	�P�Bi@����z4'�H��m��wR:Ӷ
)i��G{'^��@m�D�4:iӣJ�4'�:B��J�I���B_H�J�8��HtUl�z���>��4�=G�N�S���T*�٥�Q�FÇ�S� {�<��޳����|�
����S�U�3��^|�*9�\�=�d����i�|��k���ÿ_��͢O=Z�R�̤��{��;Y�&EnVB��K�_�7yC�s(�}�2d�go�@�W�;Id��x����|���OO�u�Իd��g�oh%���U���`���U4?���%�ҽ͹7�a�eU��gF��JۡM�q��[�ϱ�^�ǽ8�����i��S��l���)�-�.�)&�{0�0W�5�1oVj����<�� ��4����Ӟ�gW���@����4���N:k�k�!��B�Ց�s����ڻb�
��	W�Yޓ�~��M��Bu-�|�-�k
x�Q7���	�C'���*����{��T�t�K��xɦo����V��m.w[q4h�S�{�sZ繹��P������&�� y��-�{EFGe;;�A��w��G"�:Jšc�YR͗�\���Dl/��Z�eς���Ϗ:�|`;_U���V����7��>1�����H���~є��.���v/Eʈ[�+���s��3o��]�1M��ꂭ��^���Mǘ����gj���qo�����R�ctw���ٲy{��f�O����C��+M�]�)蚎�BuD!;Վ���R�zH�ܒ�*n��A���E���$s��*�=}���*�?�����DԹe�ï,Ը�T�ۺa<��`�͸��=�Gu��kQ$�K�}��*Ćܐ� A��{{0jX�e������-U�{K�̃0���|n���&�Fʥ=���Phg6E�|��=l!����{�E���1����Y���w�����Qc���M}Rc��R��e7o�+m�̠ϯj��/7W�}�s�<�~Ϡm"�S�D�u���}��i����Y�ى�˯��w���e}�J��;�Oޙ���f�u����=)s�+Mkj�U�EԎ����)�Zni�c�^�ǭM����{�ZD�/�c��')妇d�Tc�V����w��;�ō��!�Qy�t�*:͖.ݻ�.�����y`g��.�3\=����^�-��[.��e�f3�;Y��F$�������e�O8�z�P�g��w4�S[�d�uYu#��U�_���ᵡ����ef=4����{1�Ug���]����ͿI��s�Kd�d��w��>W�&s^���}�_ci63�s�A�N�6\�4�Wl��ʁ|j��z98:���>v�W�85�1���=�;�ݧ��w/�׶�v�P��OZP'1�K��r{1��q;{#�zm8ٌ�b n*7�ՙs�8��+����<�����W��V��9��8���R�����y�9o�Q�F ����:��J��Y�Q��:���2�d��f��������;G0��P�Vo4�v��I#�{���&��;龀��B��-������Nf�1���ҵ�%�Өz�(^D��Z��iyD��C�o*v~��9M�L�3��N����,b�,݇ƞ� E��@�h44lM����tU8ԃ���=X�9�z��n�ˊ�<���bq���PS*�͉�	�n���>˲��|�Miu�03j����B��T.Gm�H�|/f����M4�`�|ng��s�t�gR�����j��D�8��}.g�����j��}$��+�o%9��ϦKr�b�B@*�_hV%�]c�x�7��J"o**�����̕�	ND@?  ʪ�jf����M՟J�l�}�;�H�eE�T�`���6Wowrifu��=nNb�3/r���r8k'�Kg�5����%H�z�W�{峎2Ud���o�)�D	�A�>"��^K�i��WOw��5
Ά���A��f^y�<������H�Y��n䖧�W@�fڨp�V����Ӑ��:����5�/SJ^Mۢ�"�9�,gU���[���ehY��.����4��n��q��bj��%��DsPy�yza�����J�EE5�F.�3&��HS�hi��gu��}�Y�6M@����f�S��\7[��K�gou��<�iڙ��h��	|���o���MD�w>���'^��	T�6��gg�˛!����|>����CH_MG������u�k�Տ��VT������sd^Sx��m{B@�MO��nی�!3]���1�+�����z���#�͸.D���Ǵivgb��g�U#��#"{��3DM�}�]��mc�z}���W���?9ƹ˶[z���bn�Ց�79��8ъ�gT*�]�Y�mmk��
^x�+>����1є����2��]ED�DkH��
�l��D,��Og`N#�y�1]	��幘���ºr�D�)]w;[�4�%8��������	�D�/�lՑ��Ĝ�W��*�eZ�e��$�g��d��?*�~xQ�y��O��T1�KV����۝�0!o�<���n�LD��.7�%G�E��knF�c��G9���NL�d������uL�Wb��)����G�Ƥ>��f�T�b�U�PK*����n��{$�a<6�N�i=]����5�6&V6,{h;��y���}��K����H��9t�b^��E�@��.74�O��>h=��#�{��O0��N>s��^�@X��O�&ƥ2�M0���򺦚�tj&�����]��V<��>J�>�{�7�v����=�9���k�3 JfN�wN낐h)�)NeReg�:vv��n��9[go�W�������h�+3{�N��C�)�^���2�6Z/xvE����\eo�b�j�rXu']���C��\�u���S[.�U��y��bz���|�ZƤ_o,:�+;rZd����i}
~V7�:�����c_���r˄g~��o�*$���U�
�]ֺ��8�Q��̃�<��W������&t�oy����e��3��;Or6��.yd���;̺E���=wݭp1�K��� g���n��;e�.��.¶�$$*��cW0�����4o$��B�6�ikV��3�>��a��lpv�m�7��[]��*<G@�zv{o��:sNh�P$�H�UNƆ��e��삪����U[&��+"�����A	$�]���ERV�����Ҳ��|�o'#�J7-������v˧��N��p"�h���s)F��΅N�Ef"��(a�v1�M�q'�Xj}3o;�$]�yS1=�[�����a���܊��O�^~����E[l2�{А/�1W�����P�~����'�t�R̔��p����GlV���7�s�����p߸y}��������$��잗���^�|s_���~Feϲ4����u�ץ����֬܊�n�9�������}�|ڸ���m��C�O������gO�lH`H)��	�\�q��y��Z��l]�L��i<k:�-&�� ��t�n�Y\�pWήi��Gd&�L�箚1��X��NL4�z��0����b<�3��y$�9R�7�����k��'h�g�q�@�o-�z���{ʄ:��u���\��{�k�X��ϮR���j����GN#�M�ۘ�][�fv:-�y�16�"�#L/���mE���ʼ���vS[�CV]��W��P\Nm�ӯ1
�jS+�6�z(�W�̼��b�pG�Y�p$|I�w3o)$y�]AݗkAo��i��{�	�J��6���bv�	);�Je|�V�q�tD��6��7��N�>Y[N�7���A]S/�;W\z�X�9���l`B&[��:��G�8U&
��}���2�n:u��3�B�e�C��������P�>!��!2a$�_��~ο{�G�ؖP����I/i��670�깷�U�l�P̄���fU���I��䨦e̩���U��X�������Ӷ��Z�r50�̗;m�i��Tظ(5_��_X��w��y���7�8o��ż��ެ���]
`�en�}ˡLNœH��{ha����R{0nh��SK�y'4)w�Hc��L��mf����2�����]MKax��}׹�������dI����V⣗B�<Vٍ��/Lz�C{ƺ�GP�ǎcڔIӚt�yQ«hƓzIphћ8�s2����!@��݊�Y�]c�E��q=�Q�f�M�9_��S��`�j�s 9���O��U���a6�ޛ<#���qBQ�WQzﻻ����wwfr��Z1�۵�Ŝ�X4Λ�*��z�u9�2�3��wzX��ւ�?��~�����~p�bbN����Ѯ�Ҕ~#��PkB�t%JP4�#H�MBj�"��Ε)(J()�R��=��bH��ZB (�g�:��)))ZB��4��4@�ҧB>��(_l�T!AJД�J�3=�����ݍѷ{�
A�ZA�$FD_Ȱ�!!!��)���EM8b-��q$�i'�[�LFS>F����i�1G�QO0�]0��[�v���R�tc�Y���:�C>�B~�f\��0A�����M����̸�|��=�$�-���v�
�L�lLT��6!�m�V����h��9z�>�;�i���E��Spl�G���B���E���Tn��=�%;��b��a��%2�OF1�l뽮S}n�t�j]�^�'j�"�ݹ᫦�qF�p�����+Q|�+�ە�ca
���$�QJ��Ud��ſo W��іTƃS��K"��r`o Ӟ�2��A�~��J���i��e�a�b�NgnL7vy?�W����e�I{�*Խ�z���y5�8V��v�c[^^��:��T�w�����Ѕ�������lcN\�n�rW*�2�)0����1����:��a����/F=������[=�P7���a�|�ާ��Ծ�B?e�t��1w����q*���	ؖ{�,�M�1�Ȇ��e�'Q�#��g����컝.#���NCWuJ������7BC;}/�;6��y��5S��oF����ш��nM�֭h���}���=I��V6G=���< �e�U��-��P�f^ΌMB'�K�B��YSZϯ�MUۼ�>y.�T�ݣ��M�^82�%�i�/�)5�S���L(�z�&x4?E[���gߞ����u�����QOu��Wk��Zя�4Z�;].��ۛ�lw]
Q�)K�e ��yK��k+1W���f9�x��SK�O�}��#�<��}�����T)}��p�sV��;���x�G��#û�:���E4�A���Y�7j�۫��[2*���ϧfcw_¶��rf��H;h6�}Mn?j�f1��{V@�"�ju���!Y�^�%�V{>+�m�T�3&��{Em�ܟd�|�lCHl�X��!0#Y̬����b-������-�ʥ1qچ����'�D,���]�u��}p4!��n{�H �y�'�I��Ǖ!�V�n^��7�n�CI��ƟPU��r�C�̾{�!8Ü��j�^��N�H���g 5 j��C�-��`���|���'X�9&��BA�f�Sc��ݦB��E�m��϶e�R�"��ǅ���^�����?,�PÁ��
��cF���]�}�����塎ؓ��X�����Q�2ޑ�ugx�}�K.Q��^/9,)!���v6W.�V�vf��G��f�/��g�}ں�|�f��k�D���UV�Ω�u�R:�m拪�Q���y>hw;���;X�s������#��Op�}��l����j��Wc.���yh�՗��t�l�=%��.�{��&(�vԹFj�׸.!h=�-�5�yu���v�Â)(c��-��-�F�U���j������t4�jP��S�@���Olה<��b��Kތ���x���"�ݭ]jWtzbס�K�
��U	�����NV������KҜ�k<;�=~Y�+��t075]�Ǖ^���~Y5%��N��Qc�d�Kd���s��W�d��N�C1��3f��ؼ��뾷��[4Aك��]��-嘚�a��u�Q���Ӑ�&-�ss�L�s�X�u��!����V
��/(�$�]��wm)��Gձ�w�=pI����f>�8�x��oAu�șQw~j{=���i��o/��A.!�V{r��S0�<8|pz��,�nDM쾈�����\� �<�]�{Mo�V�v�>�ǿ�����'����	|ep��z�,$�Q���M����N���9.Vu5�8�y���\n�6�\Uw�ݟI��y� �f�yE��uz�]nB�O��EEm��em��W/9��L�ͫԙ'G���b�^��O�Y�7r�	���f*��Z!�=�.��Y)g���ԃ1�௏��^�����"ͨD�2��w)�w���t1�>�v�}�h��J��[��u�0�j�ܻ��V��>�L�`V�o!��hG�����/���qY�@FΩ�,��n���}��º���_Y�n�F�u��AdMвn]�ܬ�1K�B�~�{A?�����eV@?��J�=�`�o��)���W\ļ�R^�(Q��v�	J�{)Ju����I�����6O~��{��_>1�����e����ͩ�/4�����W'��,yͺ�����i��G6�=ޝ�Q�(�Z�{:N����E'�M覔��|ICxN�j�DΤq��&��Y]�������92o^����ܼ�7M��؏��SB��۹ȭ2eF��%S�a�����>K^H�h߬d?m(le�^r������Q�L��,�,=Ҩ�A�s7��-�����R#X���[�y��E�04=�.���vc��4f%��{ѵsW�:%�qަ�����N?��s�)�����S{Ȉ�����"+��:>�h8M�w�X��o�����/��Tp�W�y��������	�5��>�|��	���.��wy���o�o��v_rC3<E|���]����Z����k������C~aE���}[U��R��K��vԢ2��u��gg��t��`(�dc+Q���w�㑛������s����}�@���f�}�����Q��a�jyJ7�:����h/��>�$p�ǎY­�v>]���-����f�!.٤��m�Q�AU�/��vD��R��7qWt�5ep�wI��r�[�,J�Hu*r�~���g����hsy�y�jtϿ}�!��o߅:^��`>��DC�B�j1�u(���D^��FP|ueOگ���oZ��b�u�z48k���o�A�U�����S�QC� j��S�Ɂ��0�<U[B��mML��v�$��I�^�v����Z�U.9�K��4<�z�{}�!���s�����+
���eg��\�5��i�8h��x*Ude@���/Ne~���d��M�O"�rB�V-WA���gĺ����J���C�{�ևÊћz>_|�<6�<�k��:�x�|f���u�=�/����~>���Վ��~�Iuɽ�I/' �����:�`y�*����҇���N��ul=?=�Z�3��}�*�'�O�S��3��]�#c�UXڬ���4wֹ�.���xCf�jdXxg��㝺r�M�yw=�b!�o�糣�γ�{�+]�bo��&�\��V���]N��(�Ir��GFs�$�0�|{ˡ����g
r&�~�8u�۟���[�Ɯ��G��e�8�W"M����e��̵3��.k�����d�'C�y�T�-��ػu�7gՊ�4�\��(��V�0y�$i�DUr�{�(QaWq����lo�l����Q�n���l��V��K�	ٖws��JY1���gM��<$��^�oOKd{c7gJa����#�`�ך�c���X����6�噹�ȶGW0u>{�:,��	n��uX��bԡ�sj�`��b]��Ih�m�.	��P�;%��~[��D��j�w6.ev;�3��P��\�*�z��^��r��N�
wuV!
X�)53�HF�U�v�қ�y�5סt��us��q�]]|w����r��z��`��Oz���qe��:�AW�5�ԧu��q}ƱΦ��)��3�bݑ܎��[���4��Э:[<\f���:7��u6��׍z@4X��}�TI��
�w6i�'c�{�=�aW���M䊼fL�Vt��|v�R�G��2�^c
Ղ�P���"t2��a��r�rZù�i�Y��2x,��qL��`�����M�Q3�}/r��A��B��m�]�`��q�s�MV��'�����,R��T��0��d֘����٣j�9��Jv1�&d�`�2�H�b����f핅MF�b����4I�af��웦b�rJB�]r��aj�1�n�.�_aZs?��/K��v�"�E�Ua]۷J��2��S,f'Q*��e����a�F#�ΏM�"��n:7�%���A������ӻ���'-3����JY���C*����Q���a�f]yR5X��T H������M*��]�(ZZ��� ����*E�����=T*R�@�%"Ҵ�f��J&��:��iI��=+M.� ���� ���:�:���/�M+�z��N���z�Z��hӥ^���������o�"��]V;ޤ��(fd^Rq%,�S�/���un��0ޭǼ���u��-���<*�Ԩj���ʉ������t�j
��=Kv7��Y��3���7#U���Zc�׊�;�{ǜ���?*N�����To�=2v�D�p7�3Խ�O�~
�6y�KE�}$����Og�=�LW�F��5�ͭ~��w�-H��Vyxfvw:��v�*R�s.���]&��j��/:���ʑ��]���7#�AP��f��a~BS�Ypv��eu_;Ε.r}g���L^�L�Z}�����qz�v���f®'��6ފ�=���Q:�����K�=�:,L���sb�V�kgV�GL�lO)0��.�e�UJ"���>�\0�+沷�QW]��e=�w[���[��/	����^غīָQ/v�E�������!ԇ�����؇���]�Ҿ���o�{4��]�>`�X�bW6�ܫ|�^��TgWw�sg�4�M���7F�;�">���C�:׮����7��m��nj��Ѵ�x�?k�n`�L��?N�����q/�;�.�=����o+�:Io���>��L�v����X�@�8m��Mְ/�5����:k2Q�M��ed�{�r/�m�5�ww���T�r�n��L>Í٠{:P��~a-SB�1�	��"��63�\Y\��<�:6L��P� i�;����N���.�̆�a(i"�jm�)���!h����Ln�Y���6'i#�q>K��ޅ�٨���زn*�,������[%>���O.O�wfV�}��u%3�ɒ~�������g����A��N:�ݕ0�X��k�
����z�O��{_�����ڎba�� �z��/mW?b���;����ʝ�G����OF�<�r64C�|�j^g#6|�����M�*(�C�}�lW�/")UҪ��@�g���
���n�m�3ǽ�ExuF*^�S"����H�b:w��:�([}Y-�*���^@�g�����JfV)����W<����Z��<=J	Բ�i ;f�R���u�VG�*7W_�.�3Z��[�S�Cf:�����"�6�x+Ɉ��j��=ޕժ9KXz�{���<3q�kD����V��Rʃ_H��>ʥn��W���|��3���B{�SN�E_g/���[��G������w��=��?� +�;����_������vF��E(n )��ឋ��BV	uګ>�F<B[D��ز�0��x�u��&EZ�ثk�X�#�{$���Ч�7Ww�v���ps'�������e����Q?W������1�ws���E@������#˫�w+����8�Qķzf;��]��uj�72I�@9:\�9��>�����P�����{2%L������i�ɵulu+X �e9�A�އ�|h���A�$���I<H���߲���Î?}���Ím�V���<uz���]p�&Q�W���Ԃ)-Y��)�;��`a�[�z�-B���s��׾���ړOۂ��@v�csV��]���;��׎u�����H?h����Ǐ���W���}D{}�a����_�~R��3q�y{oQS�|�J�d;>ݴH<&h��n��V}�`��6F,�7�(�s�]��]��ܜ����yL��R��
]|�E�*3��w����I��h�3�Nˣ���6=�Zp�;_5/:B��[�y��{A��Ϳ��sy�d�����3�W������s�K��//�9��l]m=>tES#�l�ގz��5�u�3j{��Y����������\4�<&� ����t��_j���������[�T�j9_*�s�~���*�5�[U��&^�_f�v���ϲ�{�LK�k>��J�=�V��i��T��V�;/5�}�0r7o��Dx;"���p���N��1�y��W��[�N{v��8\��Qږ�=>���яP����v�+����_)�BXt�>��v�m�ci��k�FsHwI�j��]>�M�������}�9�yu����h�{�|�b���B,��#)��??*�?e}��v���~j٭���so�<����k\tSʯ�u<SŻ�R��nL��7hf~�d^�k��d6�J�����iP�M�4��Ɉح�Yo���\��ۑ�D�Bd�ʲ�2cuf'h��[]�Y)g�?\)�[U|�N��+�B��~}x����n��*���r���.��q�;mq�#�KV�m���a;l��Ȳ͜��#�}t�Y[y)*ӽ�I>���]����rWR�·r�Y�o����\��w}a����Ց�p�O�����~�³;����v��)���\7���,ð�(]3Z�)��:o,3�̢��¹��+gx*��E2���ӻ� ��|�Y�>2<Ǘ�j��dȣ��1���+�i5���D�Y�T��B��7`] ϭ��V���t�F�Er���NO<����9��0&杈�=�O��`�:7�wiV���l���6�ac�YGq!��=qU��D��u�ϻ���q�e�0����G28tٜ�I��yx�Z��,�1�6���c`t�ݽBMg]�����禈w�w7���Z;�O�@ � ;�$Ra\���	y�218������f�^aC��}�j�c�����f(��EX�����m@dou��Rx�:`[�š����y��Sw:�Ӑ(����r�Ĝ=��pU���h�/]��Q��ȵd<�j#��iy�h�I�/{���䔪9�Q��QM�Wx�D%�5m��y�X�g��9�����\�����LUl"�	 �6�i�Y�Wj�崚v�8η�h��c�y1�8˚���s����0��m2�}��F\�j���n���q�	�a��d\��(&���{�y����G�_�H�j������h���,�O	���-N�/HGS��c����@�FM2�.������w
/P����tݐ�h��qM���a�U�ۭ=��j�����'(o�s�cp[g`���ÆG㻷{�:��[ kH�G�L��M�H��-����Nvb:�ܻn�H���9)��5���N6��1�dL���q<J�o|��(��t���r9��ta�O7����Q��4�L0k5ʶ�G�z̘�z���QV5m�9�E��ve'~R{B��|Yz2����M���������ܡ��"��뭵8�kb�+�=ݑ��Z̮�U�.H�{�� [���H���g�l�xX9�D3>�=�4�l�^!��b�;��wz�`�Z���7�F�C�S��[��~B~�d�\�H۳�ڙ3�d��@�@�I�maGJ1�$Ax�=��hŃz��uhN�pa�F���re��� :P��q��|[�Jn�#$9�d��_K{�v� �V�Ŵ���B�c��JۦVt��ˇLM8�	�8�����i<v�zf�E>���+WÇc�DD5ƌ�\"[���%U�����M��º?�+!�P��������L��ʢYWw�ӱ���,�xs
~��v�"��K��M�0�9���5Z8���K�֮���O�=M���&��K�ޑ��W����э�e��A�?��>���'��3� �?]�߰LJ��͊�2ܹg�((�έ��:tԎ��	Õ��̛u.��XU��0�Q���ԱK�;=ϦOE;Hx�]�Bd���rjH�J�1�������O]�C�_.g��C�x��fY���ꫫ�l�#b�o5�]�f=G��I�V�+:�u�N��k�ձ��|�p���ލ�8 �rr�(;{��m8;*�>b���Z0�*$�R��v�z�������}��7�a��7骎lơ�%�n�]Mn	���,%-X�"��]�F\���	�[���M\yt6�I-�km��>�V[�C	�&�x7+��y1���+�j[]l�ɱ��=ܜw���U��tH�6ݣ�@��Ψ����۾70RҲ���:�Ω��\wA}����dV��4�XY��(R5��j�j,�u��l8BmH�f&KP��>�y+o,k�9ʢ;���"K�����̜l�#�:���K�v�fZ�,s*v�l)V�Y�;�3R���jЧb>K�N�8si��j:��p��V*�C�)��踚���9�xӺ �Ŝl�x~��n�؉�w(t|���WR��x���{ʵ�ѥa�2�T�v���\�:��L͐)*��[���P:�`k-��)]�l^��F�����t�S�0eh]V):�u���AB����P7���#���s$�Wؤ���&XlɎ��u]��#�����"��D{0v�j��Ñ�J�Q؅�cL�V9�,�3�6	t�A˽g$
_;�/`���OF�45mGC!̗T�Y�Y4m�k��Dn4Vʺ���6T��ʬS&ê�ĒI%�$���q[4�ف��
�6m���;���o�$���ꨒ�6 ECk��H��4��_���4�룡�V����	�M%>��WI�C�Ǡ(�@C��� t'BP�	�5Д�����G� S�M	��zP�:@h�"
P�OC�����PD%RP&��!��B�{�F�O��%1'@}+Ht��=������~��k�H~{�W煰܍22'��H�	FL��a�)�A�m"�a��&�,�1�Vvo<�������DQ(���l��M��4���G�yCRʼu�����M��ӭ�F6ֳ9Q�@�z���dxr�S��$k�g֊2�#��ŏ����j;��+�p��s<��T�O�o4�y�&�'�o���d��P�����p�r2i��ĉ���,3���G(_�y5�<5�Iͧ�bl(�`������e��N�t��]SJ8h3q}m/���;�>P�0�c���2��X�.{y�Ho/n�(�����axu~fCl���zN�@j"Ξ�z*5�.1�:nf{m;ͤ!�":(��_[e�씩»��0�\�hoQ.6bHD]k��0'zc����(WNbXq4ڛ��d�F�R9�5~=Hx�����Z�+b%=�����Ѵ�jjo���6m8�!]rm&�mJ�{��O�,F�<~p]-=J��/z��z*02��"�x<��8w$Z��E1���5��������d��{���r.�sۈ��<�0C��:Vt�Ӡm��ӆ�*���UN*К���tp��,=����G�,n����So0�V�_%��8���"sI3��y�
k��4Cn�#hL�29�t=�I��Q��
b,�\S��uY�1��]��p싈G S���-��c�~oY�费��/�S߇{���i�l�:D�,���Ϫ���4���ie�)K�/��]4<2�(���$c�i���@`M�=0��.3DT�oeu^�Ϊ�p�0G�(y��8�Ȣ.{I�d�x�5���9��6��<�������;�a�ƛ:t�zg)=��ə�o7��k1�2E�qo�Dq�j�W�A�'%��e�J<U����[x�P�-u87��e��W7�<7�����f�l�TƩƹ�XU�e��`��x
���֞��,F��0��ĉ�uA0:�	�)ƘY�-�F�m�h�f�� ��sN����]K��F��.۟�߳��cTG�x洞�- �����C��m6vm[dh���Ǔ#ō�O�9�>R�H�Ɓ
X��KiŎ|�!����/M����9q����`զ�Yz����Ң���P��t��Ól�M@��D?4[@|P#1F	�sA�V���+���qI���Y圿�����o�c"�~���6:�S;��
��n"��FS��2an0ްs6�x��U!�Pe�qY����"9��sW�r
d`��o���L���i��{y�̙�8�N0�\��2/�d����d��1vL�4�b�G9�.\�|�J	I�+��%z�0U㕃.��y�KԚ��s�G�V�#�l�q�3��I�EmJH쓹��sVn��败R�a���R�W����9��%������ K���fHq�B��9�w�����\��P��M^5��T�x)���Ȇxے���煳��Ca�j$���m�,́��a4;�*�Ǐ,XԷ��,5�8m��Ȗ�ne�{��f~��G
1�+����
c��3���A�DO8����,l�i�sY�oqF��?����s�s��-뷣�'�ن���B�v<Qz�t9��s
���4C'E�5���o�66�?�WG{�p�7�O���R���D��iÇ����u�'�D2���dM��r�K3f�����a.:�b�<��� s�./\?6Krm"pE`F�f�۾�Z�?��*��[3�!�*d�{��������;s����A4L6�f�k��3Q���D���7���#��Ui��`��R�������;���8g	&c�׽�
!�}��0Ѓ�C�*��Z�}f�w-xS3=aJ��N�l�1mVѴ�9"�ҭ�$��3��'���w��f6���n#��p�k����tu0G��}ə*�f�|�~�|�i(;y��ac�լO>�6B� �Ӊ�M=�[E8�}j���#C��~/���$V3��a���3���kus������D�(�P��1�8�ka��ɶף���d�'�Tuq����@�d8g"����x�Xr�?���m߯j��u�]5�6l���ܰ�n#\���۫�mP��$�\�I�`y�l�G`l-��2@
��{�(4����a���iPG�ፇBo�{�ۤ��q}��Ɇ��YE�5p��D���[_���>���UW���MA�i��}N��ļ<��'[3!\s����>.�Y���B.l�a%3�A��"�0�����1�g�͵V�o����K"yC������O��li�Vr�ob�z�v����:����
�P�\��os�v��a�i}W;\���yk���XADf����A�CѳDR������g�=Mg`x!�[��tg�A�c� 쳁-@��{�3t<���.:�Kk��3ܞN=�Π��
�SX|ɭ��1&��x����+h��Ѯ�ŵ[��r�'T�Q�f�d�$��Ю�#�*����'ZCO>���qO�g�i����K�&6R�i��3�$�/�T||dZ^8E�A��ek�E�r-����ވ��Ss�#�U4�����dC�n,���&<¹�Я�CuE4����L�� ��4n<�������]�WQ�까RyFZs�;�ŻY�`Mr�N��>�:;���������\�X�*��_{��=�0s�|�~�,�)g�|p�m��GYs��N��F��3��H�d��0lͻٍ��"q��xӓx��-�C�����_3v��L1s���1��N�T0W�=Ԏ�Gn0u*����%��: ���؞��\�=\9�
�.�¦��!�{*1�l#S�d%>,�8e�k������~�}���u�
ڂĸG�;vD)�F��e�Q�{w���E �m.5��L2[�l����
���7i��\��a�;�ყN�6<I��I�{.&a��O����Yn/����ζ6��nd���3��ʩ�����;X�"��p��4cd�xyÌw�ӌ+�{�^�P��r0D� ϽO]�v������֓�D��5ܸ��M+���x�jq��sL�[6#CK�W�_nT=:bt�['9�U{c�=�SsWz~��K�#�3Q��o��g[�M'��\�������7�<���V<�5�/!Z���c��8p`��P�vu��fnm���q1���`H!Q�GL�
g��K�C����W��V�F�~���I�B�ݭ�ힻ�8f(F���+���>��]˹���0����t��捍l.Fح���Q�lM8�#[Cm����&�8Q�ƌ8v��ٲ �?�L��o��2Jz�xg{T�ݿ{�ތk5�]7��������
��Ȼ�,8�#��5ɖ��c@�aZ�T[Z�g����XH��[7�V&z2�Y��q0ҍ[�=M$(`�٪�s`J��@l��J�)���
b����DeW�l:RU:	1��y�����"��)�Ss�N)�{ϖ�&tW�Ō}�O*�t�C�D�������i��-�ۈ!���	�á���㱴�F|�{|X'�F7\Y�4;�s�MGnbEƀ�\�"���_3��e����Í��f�]F�D˾G��~:�ZQ�Qa6�����P=o�|Ǣ�2�5AD�f뉆G�G�ǘ��'�з�7֓�VQQ�3�4�Ge�9m����e��4_�ȿ���5�:c��=[�[E�O� �j4-�����+�FP(3�M.��ߛ�c�i�0��^�݌8�TL���ֲ��~���$'�/�V&]*����ucl��n"���l!���P�6��[��;�fY73��s1������Fty��fǍ+��=5Ր�88�x�Q\s>[��q�o��j.!�� (���X�n~ �I�.�Q�uM��ooN�/�Ff�Y-�U]Q9e�Ʋ���¨{C7�u�d���aW6q�m!~�7.�jQ	���7W7�0�0�G�JϿ!4ȺP�������t�����λLw��Z�q����mŹ���g�+ih��O�����R��?t�C���o��F��>,rjSO�.�*�{�t0Ѷ�z���K��hh���\3a�
NM�W0E����\i`Egr�hi��@��@r�F�ҏi�����<0��c͏V
�b��;dW*�o�������5�׬4���N%f���#�A�pî��͟i�j'YȉN.Ov[cVs_�/�����D�փj`�c����`�C�:i��?Z=���Ф�y0>�ǩ2n�Η~b�Th�����T�q�W�� GR��0�͉�9��3ZL�aE��&�y��/z�� ?P��:'�߅�d�<�������]nH�^�"kǠ qپ/n�Ĉ:+��
�1HHWbL)OB�`q2f�&���*7�q&mM��JK�J�fփY�����[�=�$ޛtԔS�f��+q��/!/u�f��L����h��{�{
��Å��ĸ����p`�F��;��e*�xw���W	�E4h��6��u �l�A0��#2HPޙ�H��X���X��ܪ�c����
�f��׻
���2oUj�!B�k�(3����6����n�o\��S!���B�kY5��VB:st��!s�\:���,H��y$\}\W�ތ=�b�9�q�J���(h��;S�ڶ���T�^����	�w]���; ��6l�]M���M�u��ܽ�=��wa��V�A��tY�]�à�S"e<���C���6�[�r�p[�xl�����S�Z��mA���&�
tt��z(E	�t,�P�0�TjJ���U��Kɰ��.����Y�Gc�c:N*�Zq��\q�����@�׷G Ghw\Qu�:�D�ڤ^(R@�-����5a0p�#)K�ǆ��Yw�X{��}VEp�%��EɉmZЋ��e��b����i�o/��Ƨ��<��7M1G�5�������2Iu�	�g,�srƆ�k
KMi�Մ��C(���A�����|��04~�.�v$&��<vlS��J�v�[y|���	��b��bI$�X�I�qӊ�c�œ����Xa����{�T���^�D�&�I#/�|V7u\�
�@���O�P���>�{-���G�4���^�)}hF��4�������h�����Pz^���q(iq}轗B��=%	�ҷ�����@����:��Mh}h_�:��tE/@ih~�(
�ﰇ�K���B�u�>�҇Gҗg��?A�?K��t":ẬR�Ko���mܧ��;���u�t�M�f�w� >�)U~�#OkA����l/�P*S�������wM�s�����-$�QD�Rk��"K��"�Îlֲ�#��y]��ʴ�y�P���gɑxj=�G[	�~3��筪XF��R���N�qX�wZ��L��=���j���}���L�J���9[ǅ�0p�;��y�K1�k7��̑F�«b:�gj�z�D�<� >@�'������q�^�f��k$��������M� �ٌ��l$氲�k�(�>7(���/�f��hg-�7$���B�������܉�5��a֭������p{�_���|U-?��HW��%��~��{[iG4����hx����hF�G<��q���?�Y'(~�TY���}+9��)�k4'�Yl8q�v)���^�
�T��e����vr��>�Y����볯�GWgCk�o|�9|žO����_�6^��-�`y�3"3栔�����'�Q�2�k�-��Xȳ6)3�A��M���a�Ƭe�b�_["����V�L���v@t�`�A��j��s�b�"3��<h�&��H�×�wC����sz}��F�&�ٞ����>���a����Fe��s�鴄��7l�9���Wm�뗒8s������������SiR���<�%�3E��6��n8d��È|L��26��}7r�x���K�����8Si�j<tٌ��G�%ۙ6M5[	|q���e1=3vˏ�sNۍ2]�l.a����2=����Q�dr�j��s����ۆ4x�cт2���%%�3
�o-:s��߆������mG6-a]h���z�J��d��J�L7��]���9i8GY�p�ǒ�z���Oz~K+y�Sl51$���`	�ѹ�2�H0� �y&_?��uᶼs�lɃx��L�:�G��l;rr�!m�����9��j7l�6[���&d��j���Z;M/1��~�w��!�9g�HwP�G6s<������t6�U��*��֨%��;o��17,��_4]�k;!��vs����Y�yk�/[N�����Mnؚ�N��O�"hQ٩���P��,1��"���Z���r��Sm"�Ci���F鑢4Ō�~5��O}�]���G>��.Q=9�]a�`�V�c��a�i����`ɉ��L,�Í�4z�=)��8�b��y��y����*�x����(�U��Z�ޞ#`{�)3՘��y:�A���cQuO&�lz��n�&�i����w~kL>:��u��m�/��N)am�Pl�S4��SDPS6❫��a�\,\�}�f;�[{�%���iD8������H����,}f�ٷ.�j$��ʰ��sY2=�mb���Tٗ��M3'��n[�g8F̨��d�l#*]�|"�.���)��j��o��(�׹�!ð[�ھ����I�v�MH�m�g�.�NKg��t3��.�YC��ÒQ��z��r�K�1�=u�c}j8����;�5�و 3�7L�Üs�°�q��w6�	�aƧ弨��0hɄ~/�%���Ć��Ϭk���5v!���զ��$�c�p��[H�8an'{
����A
q�:l��ڒc��^�쓆·Iq�p�{8<��?�%�0�
,901�_�:K��EAdz���v'�Ң�[w@pP�Gmqj�i��i�P��*�l��v��Q}����t�ݼ�����9�V!����Ͳ��ؕU��/�HNs�xF��s6�BN�[�n�t�}r���R@�MuO9�u��{�s��<�_޶8�/��ƯŊ��`u(��w�m�~��A�:-��W6�M������	(��p�������B�ĝȾ��E\�\���<��^��Jj�{�M�e����d��f�&�%��ԜQ�%��.��F�-��T�Zٹ3��K�"����[#'N�8kjX�p�j���EǸ�l��Z]���x����.P�~1�$�dq��[�\���t���3i�����zz4��h�[�$1t�_��z�͚�-��ݾq9�n3������#�u��p�7��,�.v.�ƍ�i�S�Q�&=���A��l9�`�;�=�3�>����v��w�[u>3L�@F�Өl(�E3Y�dC��i�{�v4�h&�u]*١�r�l��%�.��-;�U�33�u�S=Ѝ��6���g]'Bo+[���U�?M�n�G�Rh}��_j��B4L�-4�<C�ƭ���c���56�(��̎��]=�[��J:h��mDa����t��~@0%��	k�;���"�i_���)���og��7/��^[�9`µ�v#>n���(�pf�lx�x���Ȉ��o1�k<�>�����W8�6�;(����ĉA���_P�R�@E�2�e�^��-<|^�t�j�����c�����MeK	��Sʺ�!�1��`k�M��c�r�ru��
5@�1E���ze͔��XF��LL;QC��4�t�q�1Ѿn2�y��v�t�ƛa�u�ك	�7��`[Q����ݿC.��gz����d��Y,�����y
k��U��ZY	dK�~�|uxy��NPݧݘzf�Ig���"�������w��ۋ��Yه	�\�kN������&��X��̼�����b�N=�im/��r%���|�?�Q
XB��ь3 t	�0���n���!�?_R��f�d�}�����	}o�Yp6	⹐��SFK���!�����"��X+i0o��4�φ�����C�\_WV�z=$�R�#�t�z/.��͚(�6&�`�
�9YSM�י�܎f�޶�&<�\ٓ�sI�i#�v��24Jv����M����:����p�V��pZ��8E�(S?t��޹L�E�=��t�>tQ
[�h.s4�Sn�����0h*�m�'�Җ����:��"畏�ύ�ʒ����dq�ځxȉ��$H���O���d�Ğ!����L���A�f���聑lΙM����0�c�gf[�I�7%�"���82�Ƃ�m�u;R��\�^��ܬ����y��G�t�}��w��k�����.y�2�.P�ʪ�G�0�M���4�0p�F3>P�n�хx��V�o�#���C�~GW�qx�|��nF9�olLBD'��Ӻ$�CO�K��o'O������+�l�=�շŲ��Q��N�YX̵��
4Ri!���]�Ǿ�h+���D�6vy��Z�q6&���A�c)護|�v N!�;W64n��D�?��)��E0ɵ��%zy�	�1����4����8�u����0�i6�p�
t{?�2g�x�G�����#%���K���f��)��M�N�nb�R�Lv[�ƥ>��C�I\�h���.�H����oR�V�d^�\�;l;8���;bi8pܰ�j8;��}�~K'����v��VO��,�6!{w6mv[O�*�ux�`�m,��S�΄��݌t�NV�x-��/��_-w��b�WZ
被�Wt�/�rO+=����X��烅oXgF����XiM�1L���$�oX�c�aUn$&ӆ9:t�m=���Z�nju����!��U1K�F������pB�ĊB3���o5��Z��X��8 -�ܰ����.0+덹z��/�5��=�L�pܛ��y��[�5��SzC�l<d�,�D��.n��i�dy[�Mb�lQ���jގCg���^F��O�~k7�wx;��58��Fy����E{E��p�A������q8ȌM!�߃�֮m�w�H�n�8�a'1�Sbj��V��g�9�⚩���N�:-�����	��a�Ec��)�qO�Nc @���X�k��Q��U<��V1<������]?5�7V�R�t��2�=��gY���eA�+$�Ԥ�v�åX��(
�Ii|H�^0���"����&V�j�!����EtIj���V�:���0�aF%l:�ζd9��š�l��ߕ�Gc@�M᷏�ٯ���������KA��0�h�jEŬ�\�o�Xa�D���GO���������#[ڝ$6�]�jm���!�[!���_	9�+�F��\�g3�\Fu�?����v���Μ"}z�h�����xߚ��3
ws�J�뵁���E,�ɡ��5Lt/��o�C�ڱ�uut^���4y�7���D�;C����ͬ"ZH�N7��&~}��X]���v<Q��'�a���>�����cI[�E�.��<z��!��m����er��y�8,<I�E44�������¸U�	xW�?��F��$���X�����9ږt��d���4��cv�p;�F`�N��6�~��ʫ�̽#P�yܥ��IY5<ݽ�&���)[g[����5��E��+�5hd�9>ӱ3��[`�i0�w�3�T�5D���/'_.���Z�qd;�j_nVw����Ў�Ι3v ��O���L�NK]z+yt6�_GF�$@޾��3��G[F7�ˬF(�JW]G�Kl(�f��N��d�u��+��xm[����\6��^�����_c59����vwe�3Nbw}HIXI�t|wn�ǯJ!<
ti^�syO����>�y��Sc�2H��|XЛZq9׹�/n]�ͱS��2Iڨ,����}w�֔ģ�k�3�n�f���[Q�LWj0���=�t7V�)b�u��&��X�l�M��e@�m$I��
	[k5Uyy�fdV�Ԣ��#mH��S�����CKR���Y�n9[y%ɸ�WF�S�V�X�z�� ��۹[u�ۣ�6*�^j��_M�#��Yy����+Q�fDB�����D����
B�է�Y���b���Z���-B%Q��e��2����{C����u�b��g^V�3;p_K��E���C�X�-s-��k�F_oK�*�$����8�"��4#.�x3hs��$�*�=f�]a
9L3a٪��$�j�\��$�KI<�B��.�V�'m_g���7��P�#�eE�E�Q��(��ʒn
ꑤN]����z�ץN�Z�o�����)([��u]�l/�E zt��O����a���@�Ѡ���A��Bt�j�ۤ6�`(OA�z�쥬���;�z:�F=�C�z:�{�Ğ�OF�����:�:�Z�Jk�讝ũ�tj��>��o�ղn�����G����G�~����]�A�=~�l(kDP$B�L#�D� ����B@�!-B��"��$�F�"�E�sZ�!�U�Q���E���n�	�NQ��s�$�����U��L���Iu{{�4�C���MM��l��pk�Et#�]��P������Kh�S���.p�"-����/uF�p�����l�p�c]
��z���Âh=	�2��e�6r�� u��Oj��h�5���v���1S�ooX�9�;YD�0)<��~�2�jl�vѢGtN��ӥsY�2XB_a���E�fL:�cb2{s\�S��oN:��K^�ȇ��ka�����d� �!��ڮ[�:XO���<�V��&��s���������u�^r��p��l��p�Q�谆�(��FJ���WDWhB�蛯NͱY��?�:j��	g�ɬ�f�(^��F�3N�3��Έm	��	��[�l���W=B�p�4X:~�vɂ�������!�ЃcwX�X��J�r��{A�}e%:�����ͫ8lL}�`'�H����J��jЍ�i�ͥ�6�\���HwQ/�X�N����E�\7b_�����>s���t�[ ���m2].ڻT�}�&�a���_����p	�b��;�"��4u�L�Ql�^�Gƫ�~�H�+-K����[�]�~g�A�XX�7�}�u�<Y��m��\������f��c����N�#�с�q��tj[N��-��a��j�uG\DҼp´Q�J�I���V�q��L�4��82�kV6��r��k���(�0tΰ�O����S�M��5��}擙]��Й��~�q��,8�~2%=��ؒ/!�0`հ��E}�g��m�tKA.�`y3�i��ɷ�V�d�l!���~�>�y��Ku"�=��:���9�,W�ԥ<������8�
���V|C5m(�j�g�̙�"�|E%K�&�u���mn�OR��%g��Z7���NK���m�U�6�o�?�6�DrrV7��f����[�׏�9�F���4�N�Ws�zǥ8���F����Ȇ����j�O��g^��b՝=l��q��M�����%�ؖ�ѯ���1��=���>��2�j�S�G8��x&L0�Y��U5"�J�2�c��z��"˂n¥��n.1�!m�íq|���iRS����l�7�<��b�
ʎ�z�4�$����ra�{f�<����i������Eg���7�@j��ko���id_uG.{݄9-�5��q�5��Έ�E�?g&�nm�3�N�H�d[e�M�}9�G}$�=Jp��r���'LȂw[M�7�*\I��� ``��*L��qB��AJ�&=����[�6��{�ԋ9���e��L�ϻعꢹ�Nz�}yx�r
ܬ4?,>��4;v�<��r̖��K���m��Z�$U7�oj��%�KG8�d`�'�wr�{~<�N(�@(�z_�f�fR���
$,��
��,ղ8Qh�ү�v(MG�5�d�:�0���$�FSi�G�쓱��_�eX6��nցt�U��]N�zvk�Z���>�/���g+�u�ƫ�<�{�O˹W���2�Q_|�U����c���ȷq��i3��e-4g���1�m�/��O!�����թ�C�)�����k��
\_7�Eo�����/�_�פϼ(� ����~U��G]`¶��t9��=ڼ�<�n3���5�,c���� �w�ޟ���NAd��O�Mjb]��n�q�e]���d���ϋ�ԼAp���ٮ�.�]s";��Oc�k��:�qS�\�'�U��8�3zff��7$5ܚI���.��̒�����s`�G��!��>h�ܐ �x��3)��J;Vĭ-�ñ�E�����x�G1 J��ϵqy.���cl�~=
X�c|�%�C��e��w��3jf���ƃ�G7fb���ӺĄ'����`��j�L#k�A
k/-|�F�H��;�g�0>�fpV[�Y�7��4n�A�w7��}-`�I��͖:a�5�h��7��^�-�M��:�$��0�sMXek��r�" r�݉�[R���{[��aeΦ&�L�(��sp;=�n�Q+��q�� 9#�t���|����ma���G�>���"��Qx����J5��.s���
�?��j���$u�ҍB���MG���w6+ <������[#�O ���_�uյ��;�2�y,/��:��47ZB���fb�D���6k]BN��N;����&��B��#�de)��n��ju�$>3��Y�ηO6�oӚ+���a���<vq��5�F=��-��]��Bv��o_T6��G���������0>�z;��P�N���!M:Ly���=ȿ�{9!���qj�#�e��9��� ��ki6�0�a�/e&
�~W���룻#�0�Hs�͵k���!�}0�vNM�ck5j���mV�s�s���aX� ����#5��,.Cd<%l]�*-Mǋ1�%�t����\��[p*�3�m�ڝ��8���&w\�8E�#t���!���&j D�kh�n�:�j���XD��m��X�Q6ȇ�ȣǌ�&�32�;d׍@�ֲ�OXh���:���F'6���34ճ/t��x��^�qt�E�?����VwC�]��]��q�0�����r��2��Ol8�i<�Op�s�������qT�}"��*6�:�D]���&��3I�O��A�a&�=������l﮽�!�[��`�c���Y�H�c)уy�@�_��y���C����'�>�v��ˌl�4��Ə��49>��Ubӓ���,�h��f2F�b�܃��Zj�2�����"�Kn%�0{S������
ܖ�k����(�S^�����	&{�:�?V���h��v�h���J�g!���h�bרL%��k#�f	��t�sQ�N5�8��+��: �0����pz)g������^Aai��P��M�Ɗ$��*]©j�����Uzu�h�j�.g2��0��QÁ��^�p�o��V����*|9-��38VuJˮn�v������[r���(lޕ�d�涜��1�����,�J]��Dx~� ;�Y�t���8�$9sfl0�mfgqK�����P]O�͝���N�k�����ƃ�a�N�鎙�9wiSY�ֈ:���L�m����[����8U>9¨�<ۥ�ͬG&�\tđ	���y��j��Q�-1��a{Kiֆ�ή:2�iҡ�&���y(�˃�r�'dc����Vj�H�cFI1j�h=��Ax�l=x�X��Վ�e�s�̬ug��e��/��JУڬZ��lVj�p� �s�7�~/(�2�p7�z��͵���V:��C���QZ�\��!�4*�T懅ryP�qv3�Y�=�?E:���_[��{�4�k�+�������^��9�	->��FK����!��,vA��؇tֳ��x�([����١Ʀ���S4!גA[Fg7*΋�aT�y�����{�'���^�:���5D��$&�e��m4�M�x��}���Z�]S�f��	�S�����<�t�0'=8E��s��\4���#
��&^ �x����=M�G5�X>�>s|�,04��Õ�hӋ��z]��aL�l�c����ч���KU�9���-��b	g�<���O�hm/�Q��1*�H��$0I��smf		5&���DS"�
�*Kj7��8q�C�m8pkq|���:�mgN�0hdw�����5;s��ńxu=0z���摑n�&��8�����9D��OL�Ӱ���~��ǚW��_xȬh!Z�ްD�!0�Y��o7R��sq�n���CN9��a���w���n����r�.fq!�m%��$][E�KGf�����j��bW��k{٢�과=�b<��$C7�M6j�K����դ9T��#�hMɅ{y��iL4�m�k��"�3Aym<=�s��x<U��Q�(�'x�lQt��M8�D8Rpbł��):�NeeKPe���Lv0����0�q���u1{���|�Mutq�731�E�����2*���f�;�L���"@����C��4��sѓ������nU��v�Vï��c�͛1)�<T{��zޛ=a���;m�v�].sǛ7_���l��p�ʖ�G��{4r[�b�Dm���T�V�d�$n��#�ץ¿zH���fӣ�9��]Z&#gw+��/gz�4t�4��Η���8FJ��������$/K"NsH�t5�/S��_[N-q>3>��� p�fG� ��} ��r�T׷�u\�JC���:�L3X�Z]��%�����д�́�K�U���B����J���Dm@Yζ,1�w���\t���l�籚ʺ��75�HG٬��P k�8d*��\�V����D�S�7�Xq��� {�^f�p�hS��������w7���h�U��$Σ�˔2�x��ޅ ���AX��]��a����e�Y�>�����K#���K���IѤ�q��2T�;y��Mc��Z79��S�Ta��;�ѕ�RVOyTk��LCs�(�͘���;�vLT�:��J�\���]Z8�f�v��4�I���SJ;��O���w�N}�����7�2:����G�]U�f�P鯶�9}li�g6��'Z��g0�V^=�%�ͺ�p���:Z�HU�=;��	�qLk�+�2��2�Gc�[C�}����G4^	5��O��i��M:wWZ"c{����;f"ˋ,�=ݼ�/��/)�Ȼ��9ìc[z�',*V'j��t�y1�+�~�ޜ �9���/�5]��-��Xb���ŋ2��l�j�[J�[y]ڴR���s4���a�Н��7G"k�s�W�Y9:�Z溢�/��P��^fN�y�u�ڰ�&H$u>�٣�kJ:���5E3z��/�}��,���1jY����R[��=͈����+>�c��36�`2����%��]D.�W.�r9��PW8�R�ٶgN\�]�a�EAt"�Hjf���1G�NҐ�.e�{�Ś�s�9v9�*RI$�I$��h�KULJ��N��L���l�W��5����}�}b����C��.���멼�V�Q?
?h����=��MkG�_뮺�m��z.�}v�}�탶
=4�qi:�_����c頮��{m��i����w�x�[��ݏu��[����WTn��>�t|O�QE��=�������*s�����>�)�z�]�`ﶚ�gLDA�x��Au���(���j���ګ��Ѣ�����S}��<A�7���4�%v�:^5����$-9{CVΓQ���9��Uф����G��4�?�C7H_��8=���"Gw�^u����̾�xW���㥵㦍Q��PR�%�f'�~�o}ޱK�^�>�8`�8��s���5��\�4��mVc�l~�{k�W9�љh*������"@Ƃ�;cA�e��aa-Ф��tU_X�cI�a��%��ĉ֣�>��8P�O;�	�Uʋ�����M�os��
5:���w�ME&�F��}ى��q��=n8�Yg���r�(�l	��/%���;��S\�p��q�&�^_ܚ)��L2m�ж�$���O(�~m"�^̛#vr	� �+�S�4_v��;��i='D�'��e(���|��צv2_���Y��|ƌ?�5����Ϥfo7KSN���g���o�A�f��ا���'S
��@Uȯ��nvح��OW/�܀�a=,>��P/%fy��/"4�Y�a=�}4t�ۗð;�q�`���@2S��VD�<�S�i�m�	��1���{6[�M����]�)���6&Ε]��T���1�h�z!^5�
��q��2$�0���rev�Kh�j�Z�u�Κ������Q��8C�@��ם�{��m&N�D�4w��:��""����"�����S��[���RdX��}L�ApU��>�����b���3��F�
� �U�����5�u�������kmm�'	�r#Xfb�v�	�ݱǱ�|Ǔ�dNA����fCA�M�qo�5b	&���� �����N#�6W����`��w�ì����!���W��:r����-�x�30���w=T����q����z^F��R!�9s4,�"��V�ܨ���x�ӣWWF5�[��	|3qB�5)9�� ��Zm�L���h���o���$��`��\g���jv�_�}�D��嫲�Z��*�lo���8����	{2�_�������I��������,}�����{���[��l��g�ɿ	��}]陖�Xd����>��,�K�5�x�c�݊Z�R�����楰FF��l���?��3H�|�Bm�_�c��i��ޞ��z��ʣ��Z�u�� ��N]Z�l��>�k�9������wo���۹�1�U%KΊ�|~4��S��2k���yT0����=S3���2�ɕx��P^�����Ü]C��K��`�o:�BK.�7��
����b��T��[Y��R���E��Ǉ!�טн�ں3��3���!���k�a�\��\�g�׊��S�ͣ�33��!��i�^�^Y�U�&���k��,W %!�� �X���s�+݈�P;,nO����fN�|rR]~]�ZOz87���W�`s���{N眛/�b!�{=c�eZ�7u~�ɱ��k!ѕڵ�~c��)�b��4s8���ʽ<E?n?+�R͢/�0_n���k�l�~ܾ~M��}�L�<�d~��ee`��Ff��WH%뾼h�Q�ʀ��]�.�y��e��,n\���Bx��gc֯כl�]�����u�©�Z�	�ޛޫ��Oն�U+�ә�"����<W2�Wug���C��MYg�R�I���ͷ��u�Ya5�<~���D��E�_��{C�C���
vun��r�O�<�X1u��F w��vV���51T��1ڌ��x�bwj��A���EN\�d�<a>W� ��
��=FR��HG[Sk�ٮG�Ξ�����b>�c!��޻�G<rH�]r쪒�H̒�Kg=n���Ӆp�.������j��n+�,�G����;�aM�^��;���{hA,ĮUI�̬��f.ڥ�Ч��8�Cy�+���8}336k�ϋ�|��/s�k���h꾬��ܓR��u���]9r)hҊ�|O=��p�x�Z���q�'�cݪD��~^���V�B���������L���VL�1�zY�n��M�R
���L�x{�>�[�h��K���6����8�z��C3b�ԧ �C_.3�66�e�m1����z��Ø�{�u��~�s� 闞Ԃ�}�߼�c�_O*�0y��g�Z[σn��s�MD����@eh\�^��6�b��@�v2_RlαB9Ï����ϫ����~Ҩ彂���z���T���+��b87�"$m�|�[�ˁ������\�2��C|���6_7|®� ���K �z29��>��weDw&.�wj�S;d3�*1�|i��5>n���q�-���DIC^��'<ks��Һn{�={U�������[_�/��L���y��:�M��:t~�}NīJnWN��w��݌��g��˜���u���
_d~][Y�8Y���I������S�d�����=�rE��=6t1�~��O1;��+<�׷q*Wk[��B�y^��ˋ~���,�''�?c��\�I=`P�\>�K������ꉓ��3^�&H�g)�y��uU�+���jOgu����,H���Q��1A
�e̧���Os9m_a��d�����6E��x$͛Osz&���ծ��˦���JT�OWK�x�{Z�% �9�>cJ��Q�X�YCAͷyh����)y��7�~#���ػ;..=�Hg3�������NU�g����Y�
#�ٌlp�W��{s�8�ɲl|�拠\���Dk���=����ut�8y�:��XH��ؔb��=+F�Dde�F{q����J6��ݟ&���T���K�'ϸ\#��ں���������U���|�{�G��Cq���,��X�������L������F=�e�E���J@�q��:��"7ȴd*T�;���^������Rk��]m�WI�IU�ٞ;�Av<��FCy^U�u��F����538��c�k�E��ֻ�E�)�,Sq��s��{Q}v5M+����~��M|B�YU_~�>!A��S�B�^�I��A�4�������W��Z�b�8ts��p����~���ձ]=�i8f�~�Q�@Xj���18�X��Ǿf�Y�B�����9��W{�~���R^1g�;�I�"	�ݒ�x%S^f;�ش�;iL��v�^S�����c;/o��v7S�</�g��^�U���k����k´V�*s�W�dN1���g��{��o��מ�K�/_gy�X��z7���t�[xv7K�������V�/)�䈌��� {I��h6�M��)&`"��z���M�3�s�z|�߱ʋ��^U
�/g�0�^��mxO[���O�*@�vM��|��e�l�>��c�j��t�	�;*/��j���,�Tlx�u��NLPO[����Jؑ�����j	��I�u�Sy�X���w?!5o�����W��죝��6�ݫh�}cۜ�[��EI��2f������܉�I֘Ø�ܟS��[㈏^�4���z��ȑ϶���s��+�v��zA�{e�i�����??���Q�'����"���UUUT��⒐�(�NR9�EE|�VA�W�c�H�����;��� ��`��������{��pJ� ��vQ1"D�,@1t���(*�_d ��?�A �x�TH""b�i�	���@o����'�?�(~W��o����J���"(��@�l������l���|��i�<s��/�H&�(��""""*"&"f**��"��� ���h�"J��"���*���f�*�j*j��*���(�����h(*
�(�*"�H��"���� �"j������"�"�"$��""��j*b������(��*������i��"�����"b�&""����j��ff�����"J ���" ������������&b����"b"����h���*"���������(�������*��"����&�*�����">Ԉ��u��L�H	�A���bג�L���(ՔD������pjȨ��
h�����(� ���Y&	"f�(�I"i�$���J��&a"fH�d����I��"`!��`��$�&��H��"d��$���
*"�f*)�) !�f��a�""H�h ���*&�"`�$�ad��("�b�	i&
h�(����Z�)�
	�������&j���*d�����������B������"���������1�>�dDQ_�����}�l�_ �1H[��"�+��eDQ�N
BIfv�����;���	�lb�����"�3��CW�M8����� Ď���DE�}A�K�L8�BD��΅�LV�BdgA�o�j̨�EWR����_�(��l�z��>Y�$A|eC�0����B��ŉ�"�ƪ߼���w��_�yt(�@��2'�"���U !��R��Cc��ŏ��>U����ia��м�E��D�6/U�9�$EW[��\>'��[H ��f�g�&�`��̢�1)�;�hwOO���2��QV��	M��Ce��.i��2�	�g)�H���wq�[ju�Ш>��/O#"z��-�r�=aq�h��+�8��~�.A�=F��}�P��{FA�������TV��DQ_`zzH�E|�t���0)���F�/@�^U$+�P:�t�EEl��D086dg%��^Q ��DUfLEV	��f��M��T
z�'���n֜0Q~@~_�`EW��~JA�;�~C�~�O��O�EdUY�n�C� M�oDE��>au:lSy�?-c���fk��S��5������I{�@L�α8brt�!;���:���n�䧷�DE�ss�Q�f(Dx���SO��>��/z�D*$B*4�� �P��BP*Р� R��P "�"�#C@%
�H� �P�� ��%ЩHR�#JЊ4 %�"�
�*�
�T --!J Ң�R�H�R�H!P��*44� R��(�C@@ Ё@- �H�P�%�/�����|/�����G�*���3�4�b;S��2���F�EVȐM <�ИA4'r4� ����R�������y}߁|��ՀQEW8U��"��bl��(w.#�k`��Uy$(���"��̉uв^A�pH�a�2����d@k�wKm�@�$��5��z�XE�::0�o�]ѼEW�������B(��`n9RBX(k,�x�jłH^B�}�Ns�K�A(u�ؐ&��@�6����"�(Hf6��